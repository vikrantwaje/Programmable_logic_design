��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z�����4��������8xT�(�h���/�<�F^[��V<v�Lz�=q{���ˁS�=Y��y�
��+J7�‿��(��ߑ��gƄ���'�j����/��b	 ���5��G��r>��T�CFT�8g>ڑh�?��H�&RXA��z�b�}'���mR��z�^��"㭄i�Y���	�׍Q�H�q��"SR�D1et�2��7���������)��M���%�dd���q�1��7q�x�(��SZu¹Qd=�u���j-�>�-��R��rG}�4|Yڮ�B&E�%��q�C�>EÅ4peш�)� ��I�|0�z�9�yw�������s䤧yM?lo�|
a����
q׷הUƸ������mn��Y�yθ��B��~��MrG/�OH[����rs����SՅO��
ޙb�	f*�谻8��>ZH ��O��V��v��ln�A���� �x ��
Cj��5���)�{g����|aM��5���={��i��J��d��c�f�aɠz��X�U	م|�T�a�f�iw�mc�Y~�V�$J3'IK��rQ4(��0�m����]�ZbO��R�+�*��56�����s��(4��}�:��!#P�Si����H��y�X.�����*���v���v4&���$���2��H���.z/wճbϻK���̮�6�?�^�ά
<�҄����Hg�$�����N���I�Twj����i�%�;4	�T�j���M3��H�f�����;sSf�q��%�f���7�=W�t�z��r�o���nn���̔��#$���Hί(u���������^��aѷ`�g����2���o��|Y��ۃ�ë�9��UƏ���-���˴$f�zS��:��A���YTS~.W_Ï^��/4�T�û����~��x��F���2��ݪ�g���U���#�zEuH�������	�/�@!�ة�h qřy[�FS�iN1�1�o] ��_G�� ���w��FÄ�����A?�
��� �+����m|��w�2�Ƒ��QP�OB�;{�/�!���0����̐߷"�N�,"�a�]��h��L�(�ROx�NG�ݾ
KmЈ/�z
�}JxtmGq��e� ����м��Z^p�$޶H	m�oQ�7�O?�S���߸�X�Tf}��Y��N��w�-��r�yؾ;͜�[M��A$S���AM���F��.�_�=��Z^<����4�YD�,F����x`7`bM�P�h�̜8�k�^�<�W�����'���.�	��0�':��;��TP����\�T3�cX#/jD�jt��1�5���/�%
P[��������%ៃ�d��Fj�pWO����K�'��iI�6���:����C��h���ޑ*A���=T�����?��7� �D0b��?�O
9�@W8���9��@�WH��M�u�����@��uJ��K�y �z'5���g�v�lTc�4i��X��`��j#��5�˶��ZT�I�^��A���z2�{/�G$�D�"��0M�L��z֫5�E��u�OeT������O�D�3By�?'|�B�Ǡ"�� ����
d��sF/���tk���)�N�� �uq����M�gC�k{vDYO;N�'�F!tG��s�$�jȅ�CU
�&�FL�;��3$�--���m���{)u&U�>-7Bm��3�?�7?W�ؠ�1^Z:���^��_]�zl�Lf��/&�� -KӃ9
D���_��V�)�sl�k�W��	Us�n:�3�����[䩽�'t�s��.NT��bA���m=<�i�f�z�C󉱛B ����e� ��ad�B������l~F^��"t\����Y���T+���V�%�0��Z��j'��d�.v�L�ٙ1��`�ɛ�_�]9g��䷂"&71 ̪��f�;���D��qN��(��<�W�9��$�@��3�x�W ��{�px����Fa�'	���P�|4�N<%�v��M�BY��r�p6F�k	�D�Ss�p��%�>����� �I�8�+=��� >���]M�a%��L�|3�jF���+���(�Y�ƺ;�bj������4��e_��Q�9$\�d�=o�4���Y��ԍ��h��ew��N�R~�&K�ˀ��xv�9WX��?�kݱ� 5Zz��v�4��)����
���5XT�V/�BV��[�Ҷ�������B��9����VY�d����6q��cW�!��pӫ��e�K	�7ha���R����|�U�y��5� �[��,kG�����v���~nՅ�=����\K`U��u̴�+�G�sE������S:�Η�I��t�4)�3|�9�gs3��eᵈ��e����C��l��:� ^�]0�W���?A+j'˃~�_�r���?OyOP��֨��F��7���TU�?����������IP�:<V{�>���ԕ3�0c��i��+
gPb�?�(�'rTWN����d�}��yṞ�l���:@��1��0ΔR�;�d)#Ri]M<�ƹLL6����=Gm�'1<.H�1h3�i�L�FSe��߾9��D2��˄��9��sL�^|� � �qVE�)�D=׬T��_`a��
EZe��(�E>��0(:΄�D��$�2���d覤�OKT3:Q�v�t�"I�a�b"�o��ps}Ò�L1��/P��B\�]�m��*]�*Ln�轴2����A�Mx|W<�!g4~ӯ�4ܶ��^_'����M�I��#qf���4����������	���e&��t'b!�k@F���L�˘��Fɫ���@��'y��־�B��IadOn}U�8�g��%Ʉ�?b�rY�
P@�����^��U��8���·�8j���.�p?��gUb�ոq�o��& �*���V@#+^���������~�ϻ�U^��7p���'�v�u��%���x��@*?��	_���b�G
���0G�c,�6m�e�I�C���y����2�D�s[ա��m�i����eT2�Q��kMf)k���;�ņ�=���/��8 ����19�?�"�˯�א�j���H燈2�.�\��Sn�)���:�<��P���c�Fg����@p	0eZZ��m 4%x�l�������!fD6��4�v��ۅU��"+��w~S��̻����B��|�	ګqr[�~^�ff9e=�h�5�(�o��� ��^��x��HS"� ��ʷP��VWq�0����ۓ�jtg,�!��J�DN�w���G�qb�Ǫ�CyW��0�6�4�|��*gP�WW��,�S�u�<E�[ܝt�p�	��C>]D���c9X��)�I�쥄�C.qr2p��G�P �%?��_o'7A�"F-]3��;g@~�]�ԄL���|>��lF.�~�����XE+	�{�������*��������8��p8?E��0��~h�^�_�:p�#�篬�����2�:���A�_�k�l�B���>Z���m��nD�X��x��hS|[G	�N�}�x9_`�2(Q����1'��ZȻb�:�W㐙�6=��,c���;bɲE ���>��I�������� �q��
o�B��`�g&o\b�7�^��3R�$O����R��*W�����NJ�;�����=�ohi���}�Dl� �����e���DQ��SI�5��D�5J=!�4'���ʬ��s�)���P�e8���C(9�=��E�
Ҥks����i����y�u�Em����J��:U�u·�<b����R���k.���6�L�O��p8��`�QsRC�(��iN�R���@�sp����Jڶe<+����T�#��;>_c(��>�{���{z�"$�� ��`թ�m]��S�5<'�e\Y[�����b�<+����t磒��Gf\3 w>�\���Zo=hcO��P媙T�`�sv�(�V��%zy�_�y�t���]Ά��z�z��C�橀�"��D�:q�y%>�!�s���E���5�M�Z��%
�����Ǻ�,���JFÐg(!�=A9��)�r1X�&Ya���N��0XL	h��<���3�k�nׂ�.5Ta��'A�+u�Y�災z���(��L�X�\8H��N!(��d��?m���'8q6Ǿ2�K�{u��� ������� �MH��_�0�n�;X	^Q�DT�4��r�g�-�fy��<GB��3��J��|��"(�0�s�N2=�;ʁ&H��wg��9� +ޏ�_��#6ާ���8]5��WK�J1����YP|�d�jG��y3,d¥=����
z�D:���Q�^�/�@$�����[�鄁�3�M�d�?jL��+��
����:�XA�l�joC��R淎<�
	�e����mį+V����n���E��n��_��|�����5�: �陪��0�=��8�k2�]�ԆT��7��d%�g�sdjw�%�d�N�	=�YQ?��7k��~�
d��3��#a�P:~�e��ǜ�� ��by��k	���@���O����')����XtN�\Z�#��v�G���g��ns-�t{8��[��bDu�>\�]H��&?S(O��5��-�p�5�2Dܭ"��"����d.�����S��t2�^���!/9�����1�dj��!��\���#����˥)vr�~�-�$uo��=�i;����E7bg��v�6�9`n��V�ʥx�.f9pGc�yo�)�{�d��*�To�J��'�'���NK��B
v���������l��o]��ѣ�uO*���oP�#��?4�?���|��ӷ���hl��-NZ�Q����vkB��i�Do��������2�;u6�|4J�Q��q ru���~������)|hrtU��:��]��z0q�+��G�]I0Cᄡ�Y{�UH`yqh>'��]}���5P���9ɇ97�f�n3?2q���}>��������)���V[�P�ſ�Cg<.�Q*�󈠄�������-�cL`C��˝���>��3^��-�c�D��	��.!������ ��"�r����jJ-%�VrXi��P���$�������p~�>�^�����5�6]�atV��[�?_��oWJ�f��N_���d=6ԧ/�Z�sP!J�����r�zX���m���o�뉳���\i�����_�d��G@M3�ಱ���|��lwy����w<p�+�գnˉ��j��b�63���G��̑�7Y$�)o7i���j�F*<�x^�yd2ܘA�q7'|�8�T�\�K
o%_��}cօ�Yd�����6,��,�\Ĺ9�,���J˙����%i�zDi
�"�[���@�^c�q�S��b�v�}��?�pSi���Uԑ��o�4P��������q)��̃���cTB��{��ME��~+
�jM*|��=3�
ql�0�_y*k��O*���g��<�Bd�I�[AɎ��Ca������1]\+��y�[ڇ����|i�i˚:���a��7���|a�����끩��������@�"3	�G���U�H���
��q�'�����0��I#�F4�@w�4�ʞ*�ņ��+`������K6�G��o�N m���v��MSt������j�i�:0��"D�� ��R��6헊���Պ�%qu��У�u+�r����`��O�%�K��
������lt�F7��C�a�+�b�0�wQف�Uԩ'`��3����ո 0Q˽\J����ژ9m@�b�.�3rJ�A�{����F�� ���N��)@��4�i�Zc8�#t��w^��`]�,�W_R%=\MQ��y�����czLГ��������wen�u����Rm~N��4� o��	�Z�U� q�+�C��:�!=��(�WM�T�X�ԸB'`D"f/����P�C�0�2m&f'��8N�Q�ƈY��?9���(;}d�{��m�8��5�_��uZe��4�Bĩ�t�������-��
���"u�����o�>eA[�;'K��]��`E�9��?W���W�^��#�G�����ί��z
Z���	�(o�ƚO�ȼ齆���m�"F0�qS:;����(�f�F�y�[�Y��wn<م�>��A�1�lq��Ṇ�+k��0a�$��j9P�,A�D�Fg<X��� ᳽A�/�@浩R�wS�Y��L�?1�5�4��R�U0`֒T�ی%����O.�7&��](d�w]ez����P~9�4����/@���FK�#%��u��i�4����ÿ��?�KwɊ�#k��U�a(j�Ь�Uq^�}��[�ˬ8G�=��n�D<��n��"HJL�;��J4��g�����2FNn�O���aU�d����FZ���\S!��w%{h	΂PC\GY�a,kXR�"01�~�:�f.i�v��6�-UN����٠��KUSr�+�T
e���%�����VՎ|�૬��= ���gE����X꺦�ؓ���n�-7��RD�	��4:#��l؆6�KH��8$죭+4�%��$�C-@3w��I�8��P��(��=��ĴV���oȰ����\m'����6B�l<� z���L2��J��6 ��w>�_�I��N�kT�-���wWg�jg��5v�{";���������j5¡^��6�U��/��Ʉ� �ҘK��=�
m��]��FNS��\��?��]�cL�ws����!fj��ïk���n�#\���FȃkVP�j�SuN�7�gG^�X!�%%�?x��$��s��iL�U���j�� �߲�\x�ar�K���bFǢc)�nR��6@�x�m�|W��q���+����X${d�Ŀ��6��?�Ք� ���cV����Eq����	�D�&DV�3��((|���#+)�?4��9�h�����t��������F�jK�akg\e��0����h��=��L��˩leA���ȟ���f�5�YX:�E�s�3JfH���8A�r�ʫ�:{t�4
p��|^�6B�1������+�zI��0���Xs��MO��,<�˅ל4�~s���qmk�
-#�Q|�ZBʍK9ܿ�U���Ͼ�m�R+�-l�J����G%����V�D�=<"R��?�48q��>
�Y���%�N����+dstRp�\L���8����l����W��z�u��k�2���R���M\�Zz��75���;W�<�3Q��/cy���k�j��i���ʵ�� �#�������w��v���N�z6N�ƿ�S���٧��y�^[�M�I�2�r�/���D�� ��2��vbyI$�s�I���z��ʠ�v�É�b��
���4>G@�ȇ�ʉRl��T�����7�H��.X2G��i��.B�Ȥ�u�]��\���R��*Be��a�ޠB����(Cl���\/�C��1?5�ǚń�*��ǠeＪ���jhː�LqY���&3�#���v&cE(����o���pgw��ʾa]����&�V����)A;9�~x��֣�H]��`jo��=�Pd5��(�c���x���K��E���u��G�c(�̛�vY�gB�:ހ��������Gӑp@₄ˎ`�T�y(ɽ�aݛx��"S��|i�&<��sB�r�PS����V7�cm`��;�s�#EW�pT ���[����K�N/T(x�]�-��p��%��K�vQ��2�l��h�[��oq;�Ks�I#q�%��W�I���%Q�r�:$�X�\���: /��^�יHӲ�m���84�w�,��JQ��f����lPcR�I*��������+ ����ZvR-DN���z�1�^��D�C�^X���G�r������oX�P�'R�����X/�w�	�A�_�	"*��K�+0��0�g�7<xgg0S(���k8uܔ�U���c�R:�J�Uo��ӝǓU��Wv(K"����L@n����p���Ȓ�+�k�<0�vC�`�uS<�'�O�G�~�L�<���M#�0�9�8��s��K������xR���p��mcm�R+��s|i����%>c�+�e�� ��j"��P�<�@���yR�o�k�2��.Sl�RՃ�3��+�U�Z�y�F�}�ɧ�ִs`�(�L#����T�<�1�D2$Sbך���E��{("�����3уHʺ�'�8sh��pB8����D&�) ��~�V�mz�M[p��+�����G�Q���0�J�e���p(�: ��P�-3���������.�Pٶ�סfE5�����o}�gTe�U�����tnu	�������8~ �ݩPg��P����^��U�mY��,�v�>*x�R�q�s���:�yF��������R)I[�0�r��L����4�|	�կ��P�z���!��D7w��q0�P��r�<�h�)ܺ_���f~���A��*b�������(����Z�1n��D�֑�_U�/$"�j�b�M&�97T@�%�\��a�%/B����Y�w��o;(����޳։O�蛹��ؽ.�j~v�6���I�9��ɁU��H��<��ų�l��ra�$����R=`C�YVMZ�H�eS�8�OA<� Z�یeЄ���i�5���<V�筒��l�U7ђ�88�%aW<��I��\ФM��5X%��z�7�˧�Ů�r2Oȸ1c�d�^(yH�U�ݗY��d�غg�0�<p���][�i�33�+�u�	.��E�{�j��jߒǱ���S�vه�١�0��	N���ϛ\H�ڥGx�j�Yh��v���%y��D�w�_�>�z �>�/�Q�me{@�s|V��;�B�۔^���{���wH��e� ��E�7��_lB'e����.��� E%03���vf�i�V�ȱL�/-�h��h�yEژ������Q�����BҾ��~3�'��Ȼ����j�
��S��X���'O�a����=+e�y�g�E�f��M�VN�ie�ߗ�H	��_�����{�<�OPIVx0r ���8v�-W5��� 5;7r|�]Z��{�����H���hF\������[;��S�8�[T��V^�cj�P�B��S��UH=�(��;Cs�F���	��>B�aԓG+i�������LX����bӯB�����bQޒ��~b�W�N�&w�����q_J�\7gj�{Ʀtf���7�m�xR���+�,6e����Mܠ~>�Mq�SC8��d�.*�hQ\)�C�@Z���>�L:<�� �!��9�����N
�]z��`.!7\涟�q5�����"�^��sq��^h3�Ӵ�[��b��ҭ�U22����ha>D(K��Z�,�@�x��UJm"��K}���5=@�u.�TX�T0:��/q_�h���b����_>;����Ⱥ�R�$=ܰ�2�%bG���i
����Y˼����s��q@jG�s+Ҽ�v/�t�F��*��ՙ��j�S����$�h���+�.E�q�|��DWfI�c�������E}'&yJ�ҿ!�vY��A��B����M����L@��]^BT�(�N��?$f��Gw�oަ��d����]�O\��?�[���m"b��� xYx�@]J��nm��7��H�|�)u�9��R�Є���H߰p�2�HJ�Jز�l<[�T�Gt�b�Sf���f����
e��A����%�ݝy
z1���Zh���FP�֚q�\(�V<��s�!`�7V�-'�`M���b�j�L]pE����[�E���ȍ������U�P[Z���{�����KwWUt�uץ���D�j���-H���c�V+��^��Ǿ��[ʝd���^tW�{7�Z&�a��Ų�!<<):�����}?��LaP����L�������~�坬¾ZP{��B\c�`{����w҆9��M��e3� /�3=�����u��.����7f�8K�� ��hL�!!���B:�⭊�*T��l�+~��BK��4LD7GFf_@�s%��Q.����!�K�g=�6)Μ�E�]��)u�N�[��Mw�*�gA*F��	���O����&�f
��q^U8	�RT��?T��+l��U�b�|\��U�dG�(�V��	�y�A�Xh�\vߠi��D�y8g�|�#����w�t��-�xW��u���� ���4K�[:�n�+��ņ*�����b��ֈݾ{�ҟ �GRkFx!��� �����u7�M���F�:-��4OF,J��Չe򿹢ζ��)~�්;߽�F��a�u����_��/�cx�-M��Y\&�߭���N`A��^D���O	��ߎF4��v�!��7�u;�:��0	oO"w��0bx\��٫X]�8�qm�,�@^N�5����c8 �>��	6y��"����`�x����+��^&1��(� *�D!2��%٥���ś�_q�"�D����GZ M�qmY��s�Q�{��WPJ�o'��Ϡ֓`�6�g�p�"�9f�~0����а��{[)Jp9�D��|�DmN!;@)��?ae��K�S��N��V�d�i$�/g]H�<�?	&����y�cA���4Cz:����L�E`\�/lD�C��U����+5f&[�S�y�1}��O��tS� ���8P|r�S�ɇ^P�걊�F�I7r��������r9ab%򣱀����1ג�m���������hE�I��(��S2-�z��a�+tNkÀ��l#���M����~e؜÷�^t��*�]
�00��]�s��B�B|	�߯uq��2��&2C��QUl6w��.��!"�m��r��K3��@��n��Y�����Bu�N�Y��_AL05W� �듥`
նc����\����&�j^�r&��J�4�1�f��GB�L�w9����KP:�`:Yn���AR������։+t-�D�x���W`@G�)Y�$q��Z5*����\�k���CK�M"���K^���h��*K4:6�B�ghsD�4	^����;�ϝ��@�eR�H!�r���Q��@6�|6�uni�
8 �_������~�F��c58���.�����E�����;`KE�t��lj�_Xs�mH�v��'H$�tB~���"��d´T��B�g3w�����J�8G�2Q�Ea��ʖ4���hF�k�6"x�Btƕ��h�qRI�hW��_�9f�x��$�)Mi�����T{�Xg.�
��E�)�&�}�VԧN�H?ñD��Ƀǅ_�d�U�6�ͱi��� .�P���to��G�׸��VF�ٓ۬ �!��;ڝ��l_ъ�cE\}�4��u���Y�^�d�b�a�P��Q���j�%T
�i�E���nI�HȬ�#��7��}����x>|�6ZO����z�-��v?U�7��c�V��UeNې��DCJ��ڝ'L)/ǆ��z���U�
Vܼ��vT��ٸd�d�z���M��j�S�[����Θ����&Tf}�0�]�G��v�J"���YV	�P�Z<���
g�R� �����܍�],�%��zE�qUDK��4�X�l��u���m��T�[v��j��q�B���pX�L����)���>�;�LR0Z��3#����7�m��)Α.'�M#vq"�п��s���\9��ۃlu��'����7P��А����ف�Y���"A����U��?�@���Q��$Y��OX����R>�9�A�����
�ExӔ}(P �Z0Ђ���6 _��_�Tk�Ҁ���(��Z(W�s'�9[�c�;>�5�F�-���k�$/��)*���N��~�$�G&x���YNy�T�ֹ8�)j�ra'������~h�<�T��<\��������R�X�w���(YNҞAr����Ms�M�j.���d�+���V4���M۸C9��AM�n��xz�����Z�)��q����B���u?7M��@����V@�.�?��O̭�N�����	3���K�Q\�+��
]���Eط�p��0�"�z۹(+��1�g���D׿{��G��m,Iw��H����#�8q����%;�. W�l��!F�|?��2<t�Ԣ_�ҾɁLg��Z0�pͦ��� 9!�����Q�|�#�Jq���AP����t$S�I�@|�駠��oԣ�ҟ��@�9�z�D�z�����7NAx	iI��l=Gw����p�Zw2FjP�Ö֫V��nQTVS۶����c�Hrv�L?͟xw��vljL���]�{F���,I�-Og{�`�?6+iq��P7�=i,\1�m���i�������#���a͞<jb�_$Iߡ�#ݥ̦UCe�ϰx����`��̵��/�_���*5��խ�d�4�'D!,�(Mv�E	�����%SkD#���4q���y��jX�r����`.j���Ü'Rj��K�����m����>U���a~�������W��ā=�s�p_Vz`�L���a�S^&��F3�f��ՙS	f��;��e�z~3����3�%s�sR\5*z߁���8�&�ԍ�[��4�P�a�_�v7���t�xv���l �Y=��]��,ץ�C�ܼH i�h!շ�2m�"{]ȁ�Q�7n�d9-O,��ਸ�F��>�j�Y>j�V�7�P4.y��i:m ��8�I�&Y����>5�p�� ������Xa(2��_w�fL>��R+�G�w���\����;��m�[B�/=E�X�!�FM+���h�;(+'���}laIv�{��&�ೄF&�-BAsv�9�*�����nq ��:e �9�d1��qܢ�F���ω\8��UW|U��x'u�m�� R����I6�0��B��j�n F��1�`0}׹��Ɏ�1����]��� B�ﴔ1�����j/��s%��z/t
3Ʌ�_$\(���������M��G�'8��0	��:\�%�ڵ6㣯MO��Et��B�����	�.u-�3�̮��3ߠZӁVBv���Ӡ�TʄO���Z�P��or�3�)��;�G)�)�]u�`M! �_��)���h0���5��ԣL{5��j�U*k�������1�)����e�L_�c�Cs+M�n܉-4��3��2��
���H�����	��uYJ:z�a�U�W��9�t���а&��㚹������K�-�a��7�4D@���	��昑xJ��oȦ�B�`=@-Mh����A�,�� �{�-j���odggV'>&�Q������ǀTQ������ ^"�ҏX^Zr_�R:Z��4��a.*̿Y���M���c�ڏl�A���[G�l�M�OIg������,V�U6t�\&��rĳ�N���O����U�D���T���$�z�_U�g�3k����t,�E5]�wܶ�~w�/�a��]wc�x�����io]�[]�7!��e�p��w[�hP$��v�p%��B�ˎV=Y5������HL%R$ �-��X%y-���e>��Ny����/��l��S#��!��?3�*3`����q�'j�tJ� �~́�q��9�2��
Jtg���'�z�I�[�<�H�i�	+��<u���i����$-t�i0��z̴����$=U�s�J�ܢ8
j�O�Rt���;ʛ�_.���R%hk�]�%��mK3Z���x.M� ��h@�%Jݮ�i��M;�9����A��~�7.�l���WE�lؠu�*���	�Q��ȡ������X����2Mhh�3L��y��QE�\�СQ��j�eVA�8���|�X2ۚ6���-�;5�N�	{��L��驏2uk�y�����䠼��H1q���C�+�:z/y���'߫��ߐ'@jS���D?kI=/\T�΃�N|ީ���Wx���]�&���]E�r� �ӄ�gsdD����	h����"�/��h�J5�+'�G�����ד�xiqS�ٛTE~MZ�sL���޿SeV��!��R���Ӣ�,��l����_�
�B`x�Q.�|��d��{���w(�~VH4������0F"U8	�ll��{n�v��[+W��a���WO����5uM27� �6��.������T�[���}��gÁ>��?� G���՟C�o���[��Ʊ�p���*��jƜ}�����l��	bF�Y�g����ַ�(���XTbд��`&5H�5�%�F��-��c3a�������1��I� EA))���Q���m&�F���v~O\;�%PS�r%.�����K�_�K�G*!��AÙ�6�@×�, Q�^t����+���Ϻ{r�]�����$���|U�C�� I�OI�N]HC���=��=#g���n#\zjd6_vV[��	�GzX�A��K�lSP&����>t:4J��r�;]��ٿJ�V���<�/)?f,e�6D4:7:�r�4ï��*�!���P*hk-ռV��](G��ĩ�1?���5��F�Ԏ���?��l=�����RS�5B��՛�%P�
�R��S֓������F��i����N=�;N;�-)�,��"�V>P���S|��5�S�tvdH�����T��d,��8!)Z��9C{���t���-+��W�g����N.��$8�pt�M�z��H��/�� pͿh���9�	��lh��0��mC�`��CZEB-��tc�]:S�ikwE�:�Z
;�h��k2��Y�*�{t��h��)X/,�N�l��-,�A�Ʌ��.�z���Cy��F u�r��/�� N�,���ܛ����iN��=���P��a�(�}�����ݙ(�b��u"n��K�Sb�7⟼,#lc�OTc��j5?5��Sɪx���9.h�;��\:O��]��ʱ���ne���~t%Z����W�B|�
h��ۚʌQ��縈'{��!��g8�jKS硘�C�o������4�'1��|X��]�9(v��C��������0�#{�́}�A @6�
�:��ZԊ�����1��Y�J;o<�v�w$C����V�\'^p�� 0Kx&��N~Y�|���m�>C��*ӼmjU�#%��.�a����w*~i���ånvgs��5?H�u&t�H��G��K��D�/X`��=1���A�x�y�<��mWE� ��:nx%��t.Bp�2 �&��3�*(����N��5����W #?g{ ۅmW,,Wt��`��?I�c���L;Y?
v�n1�A��u�Y0�����z�q5�U>����oy��XV%iW�ҷ�Ǎ��=�,<ޮ�I��Ihvw�=��t�sƮ�1+��t�b����؞��j��P  ��<D�ӧ��BD�,n��2 �I�s��t0���� �k����|�-ec51;�BI��|t�p�î���IbhI��(�-��!+Q����h�mu���9�]@G@�j���K�vro6�C�s�H�NC\N�ʿؕt]��8��8�j�4��0�8�z��s�����@�~��($*<�QN׻uT��C�6	2������8P畣^�B��x.�)��l�"�a��銖N�|�b.����w[�]�Nm�;���՗]��E3	���hc�>R���tiJ"n�Ǽ����.z���=���xT,�����=��B���7b"�*^��T;A=�\W�Vu����V�fM��M��ED~yg�^1�55����&��m]�-%�-dh�����+���5����݀θύ2U��z4A�Td8����I!O�2�-EUm"N�ycRRN�n�ZBB�bՊ�8��ܪbg�3E�*�Ej2�F�aN�C�œ�f�Ŧ�g�ΐ�C	**{���P_3`���>"��.���o��y9�N�Ȟ-��%ι�-��_r�6m�C�	�)Qu#7�I�����{�r���)���߂�n��HJ��y&P[I,2B�?[��9�!L��Ǝ�yz
ŀ��B��]yW�K�� ���q��
����w��m ��b$��QQt�.`A��\s��b����4����.�wXħ�^�鲾U%����~�\�(���ݧz뽺�$��z#dSp<��I.��2��|�^?��ح�?�p�
�hϔ�T��8���m��j��@mUː@��⎢?�|;����3}��p�[�۾o�t��c��"��$��y���i��^�h��E�#=��u�ğ- ����������R�3�5dQT &�ŉ��0�v3��쳍�5��O�}���uk���@�p��238���B(J�!�G���xg�ƿ=ĊYИ�M��>B�h��������jQӠl7�b~��M��U�V��������i�¥�q܅�����ᒈ�[�ir[���{���D>���9�W ��h�ȫ�?�_@��Y��y�;�˹�]*�o����n�_ɬ��M�)��o��o��n$�ף9�jDx�-�e�o�Е� 0h�?T��cWW���K+�0�8^��֋J������Ϳo��p��.����P�I�}��t8/|4�GU�����6{�ѳٹ/4 z����TQ8��`��a��t����� ��ɲ		�� &��Ė��-��N9�p����$��A�	6;z��qH���� �b��S�.:q�����T&sS���T&��J�k�<�Iw~jթ˅BH���������a��+=�Uy�Ymt�#�����EN*_�ƌ1�[��w�6�?;8oGV�h�M�:����r������}-͠q���3���K���1Hx Y�l�c����P��l:���M����Aa��:���J��Ҹ���B���7W�	��ڂB�����f�ʷEڙ�K��6�7 Gn�g��1i�Z,�^f�N�������,ɗ2��6X'�H�JNL��.dw�[�`������ow~��R��d8���Ɍ]���7�f̸��&���qN��`G�k���Z*�`�-��(ORg��b�s��3���ՋEk&��D�,f��CAM^(��Ys�J���t�&�a��?V[�ZZ�'��Y�z���t��<_�o �BX�c�T�XYYS���+��ﱿ���s���pcd�`t�u^�?�Y^�ź�%�B��8~���q�)�)X������H�_u=��i����/qPs�����J�&�v*�o�ĺC����`O����6�0�l�F�HcP��X6ǖ�_�h���x��E˱��1����!�e-�.�ĸ�O�C��X����U;��v��;X�T�Qޮ�ކ�xg��W�g�C		.��2�H����KO�##:=�7 #�"3�쾷�a�(n���U��չ*���XԒ>�e�ۡ���|L�S����m�����*��Pt{t�]�>�m
amOв_47[^:�M���<���ޱ4k*T��t����n�/C	0��~%`��q��J��O�c��ƌ��9�l7U��o��/���|��V�h/a�u��q1p���2�
�7j�tnU |���Ui�r�P��A1�#���;����ݫ�r_g���� х��w�ec�p�����)��l�`��g��#Y�����e2�[岁$��4�B?��~�_â�౒����i�Mܯ7��B�7f��Q����_*�����Q�U�j��n�m��()��n�����ַ@����2wDvf�ێ۪���yj����1J�yp)��7�̈́�
Њ�S�<A2�� ��Y��\�̦L����jѧ`Ѩ�`���q;�%lZ�P����L.�n�.�A �?����Ν�&����.��WY�(�������uo�{�줹�m�U���׬t�f�G��6������9
�.ـכ�븼��[\�u�B����'�U�0o��V娸"���/?B^#wjĖF���v�\,����4NWyFN23�(x��v)z8��� ���_P��$�-ڭu��:���n����%l���Ӫ's�L=���� >����ޞ-�@0yZ�R�MJ�D&�S!�HѨrC�M�v=R�a��╒m��ȡI�S�%
?�}����PP��QIfU]'����K�Sæ���C#���-u����pI6�eD��P�n���y�y�6Φ�<�?E�N*�R���(�̎���c*B�.�aZ8��"�@���g|J����Q��ϓ�
�IX�렊rf͝;��rWS�u)��9"�O��`�������k�I2x;�ŷ`q�b!���%H�C,~�#�?��8B~t�w�3�Ɓ�nw�A����=��4�c�>�z�#Ȕ��E�>GC�����0�M�,��m^	k�/�")���%�N!%&:8J�G׀�r&��2B�e����-��o4wr�KH�8�hr�#@c�i������[y�[b��,\���".I��*�3IH"|����Wߕ� Ƚ>��J���3:
~X�E�!�q�9��e�؟튩U;I-]^Iv�w�E�V���A�������r��qH�t�����j �����J�D)���il��_<�@H ���"M��b1�2S��tN)�V���O�0d�y��H���{�{���n�Y��r��4V��ր���X�|ºt��S1�9^������>�85�[��p5��?a��YlU$�[�Y�(O��z�ui��Dv��}mԈ΋���"�[D?�3�Vg:���U�xq�i"��o����
#��%�D^�S����ٱ��8��y�"�d>����F��}�E��z{�2<�զnRf��޸;}�b�hy V�J�7�g0�O#6y��N�ʚ�?�\0O�A�tM�J���o��lT�k�>��6`�pZ����O�[���Wb��g��v'�ـ(���z�}���nx�������Qs�b��S����H�B� ΃<�Jg�PB�ő{��
2kok|�'��!0�����Y�z�ȋ[�1���D�X"���%��
E� �Õ����r#r��K� -��曻,�ח��wA��(# �ɍy%��X��Q�)Q��h�ڐ�f�)(�6Oe3��G��	�LV�l[�h'q0	
���K����L�wxly��"i��kQ�@-fاj�(�Lsn����5���M��q䃃�K[0�a�`nzԍ�
�O�d_�f"�d�K��O
-ې?�!��s��M)���OM-7Ύ�����DQ���[k �a�kU�үf�Ns-]��j�k�D�mY��u3��:�B4�=�ÖS�3rm�����*��nD{$L�rse�x�ư.��[�(�%E�{'�#b��0vp�;�[���)/��W5F�Q>�q��6К��(�D�5�}���e	�X�\ꬋ�!&v�67C���O�ʻS�7�5�N[�Fל���@ɞ��'е{��|��T��N	;:������[��Տ/T��{Z��%���7O	�&���K�D�_m��ib�=�9������x�!K	�tv��Cg!Y�ݸ�n��1���	�,��u����d>
�5֍���k���>���0��7mM�f5G��f��&�[���dR���CI��ڡ��ݞ]��T[R9L~
����CD$�8RdPsٙR��d�M�$���i�eri�X��oD.{���'t�d�4���~���||E�(w%1̎'HP�>��(⤿�IV���K	�E%�J-�lgKv"��&����^��;ߖs�O���R�:�����>��"�9�IC��LwC"����@��ٙ���*f��ԋ�6��b}�F��B�ߥ�Ǆ��sg]�M��0庖:����:=�\���lhT�P��9���}�|�hQ�A�3B�%��O.�L.�7���@�f�=�(�(�/t�J�&�u_��Ǌ�Ӱ8��W:�ԭ�ΩUK�#"��.6����Y�f���;����}�����P��͡�J-bL�!�# �����+�� 0M��`���y	�w��!�6�0�3�]��擜��V���+�\�uPWG�G��}G��5�/�OeTI�>�.RT��3ERJtdu�F�U���*�35a(Y`̵r�7�����������>M��ݚ�w�����c�B*$p{Z�^�8%��-���CG�!�u괅/X�u�����*4/Q,}��?�*�_��.�$��t��((P��~5.�EOܿ�-x�Q�/5*�i���vl���~,�%ݿOůVɃ��v���c�Ҳ�e�V�7�����0��I2����{�=gF쉧WX[�َ����"D�#�R�m�@��71��X.����6Mn��N
o�'��6d�"Ļ�S2�m�;�lv6s@Q:d�&q���������|R�Ui��[� ����k����w�|ee)N7���hN"%f^�ׁ#N�<�dE�D��y����Z0c����r��@�I���֍*��LSSԧ��g��u��i�A��p@v�5:]�Ys��V:xO�RA���
��6W�I��/	��< ��pĽ�&v_@'�|g�[�~:\b���Km�Ľ�u�S�@���o0�XD][�����'�}8��VA��<���D�
�nd>��P@e5ׇ�N'�Q�w���\��Cy>��|$�B���羑<����f�z���'F/��v���7��*1 +_���x�7!\�W�}���g:���>�H�t8	�ꏉ@��}+�p�һIꨬE."��E��O.���ұ���>�n�﫰Y�:��°��*��z�A��J��Q�E���}�I��>x.�腠�T��b���g�D�f��3�����Ƭ�v˿t(�hz���hr)2G�8V��FN�V!���Āי�d��5�a�Æ��5��FJ��Ӧ�R��\�T<	_��'�-�$o1�9!����~��s�`�{њ�,ډ��9n�d%��&ē�\����a!�1K��;X����@)�G�D�U?o�)��b��!�6�>��o?>��tN��L��~��^�\����9\T��RC����aПՠR��U�S�ܲx����M��ޥY&i7� �=1;�m���UKӗ�����P�
��e>�|�j5	���R=f6^�R��%�R�M- �aH� $�*�C�*��;	}��ɭ��2�n�.-�b���F�u7�?�G���i�<A�?����gu1�����
���������G�3~����ױ��Dg��1������t�ݾ͢���]��:���3iӫ~������Տp1�A\Nw�^"��k{3�6������I��qM.Ma��R��J�@�ȔhV�T'g�\شSg�O�\�?�w��m�u]��P�0��0��͎]�SJT�(
* R1��� ��ZR�P�ZVW��~4�v�~^���B�%.���t��w�4Lq�t��ݐ���$p/��|�e�I����9���4c�-�dv[�݊]��ݡ�c�!"�;�s_I��aʛ�l�G����м��1�8�^>��.��S��I�Rax�."�a-��=MvM:��%j6&����2��<�
��T1�ˉT��B�	 laϣ���T��Y ͓�;�c��Ȋƣ���C���{�쯄Z��*�w�gLoa�
(���U�$?�)0�/
%*��܌*n�&	x�%��0Śд0�/ .C��i�\ODX~���K�4���|�C�[K_�E�w�\�J�!�1ѤΆ��hy��뙍�f�t�?�c�dt���#K��$~����֓�I	���2�Z*9�l�"�;�4��}����.��裔v��D?/��Q�9�*<;@�\>�Z�KA�p�8�plm%�����@������6��傺�}4�q3��jshO��e.�/��Q��^�4i���~>�^�G�Fbt��i�;��2O.,?9&G���r����ԉ Ys����?�3`����c?�GF`$��ͽ�V��5V���l}شY��4I�u�s\CݥK9�i�拴�.��"[=Z�w���t���$���r�W�t1�{ EJ���mr�"L-μR$�����h�h���˗c��
6��۵���Ċ��b�D-YX��H����Z�w�9��l����ж>��;��W(�'�����ɂ߹�lv`��>�lndFB��u�*2/P��*�2�D>�+OQ߸A�z�����P�� �d�;���fE�g�b�=Ӑ���h�����FVHW�#���H��\bBϷ߄,��Jڨ1�g:��M9x�"Fd}i�`�=���|�n�_����m��RׇL�N������+�^�NtBc,D��:�#$ɪȒ�{�|�:檫��3���Z9@ϼ��7q�%^������᭟�2��d���
��;;d�Or06�²o԰)��������ʽ����c��5��,�&���1*�]u���~�A��8�q"8�ZlG|qU}�l���&�[B �e���j�����:5�'��V �2 و+��R;���u;�)�m���sN��gj{Q����yro�'�Ԍe�E۹�"-'��p��Q�AF,�k�>db��e�:S'��8ɸ�l~':PX����6C�Żh���k�kaum�(3ƌ��.d��䜣���P�)��䵳!oj���*��xu�!U͎T�Jc�
��s�\��&��4�>�:��g���w9���M��$��-��6.kZ־K��9R�ì��^�~����g)��t���p�<�)�HwB���nC"a��L�>�l�!-ko�v=t�l#��l�ϋ/֓ uί�w]R�0��4��U !�a/L_��䪤�*�\�dj�Ia�#��r��ߨ�D]�����P�5p���<����x]�Yn�,!#�b2�}���h���q��a�����/�4l����̖��c��$��(Jh�9@E	�!p��B��	BΉ�J0[4E��b;�0?�	b��Ip[��aD1Z�8ڌ ��qO���L�����ѻPf��K�2V-W�������R&-���{�k��-�~#q'����B�w�$�yj�D�	��|jvи�ݓ�}���r��Ǳ���EÆ]�,#�Q
'�]��D���U�{Tk{d#�w�X+Է��4+S?�*�
m��p��Rq����s����,}��8���ۙI���d����� �6ixXBZ�����FJ=�y-X=��=�N�l�b���!�o�\��$��\�'QGg�}߳�b�����[;M|r�n^��0n��f�Z��Z�	�>Gʒ�FGb���8S	�h��|{K6h�`�����UzDھ*� ��x�\� �M��� �[ǳ˺�rJv�T�RPY8�qo��]���F�e)��<�d����ް�Þ���&rF���,�M��j��(���a�GN��U�;ݕ]�~���;�%(G8��'>���{�����Z��˩'��H�4��u9��8@�'%w4��3z���������:a�^x�v�8��ЌZ�;�RX�S�����ܹ�0H����Ƃ�cvtXtL`m�Q3�`���+��2JA���}��fom����|��y�U�R�����	�
��ԲD���?��B��ul;uV�zQ��}y��L���IdZU������a7|���=n,?P��e�h���R�iK���x�;�:�@�3ϱd������*�>$#�]�b��6��A�^�*k��5]�@��r	9Bm훻��@��JM��N�<����vMr;�D�͐�;B���Ev82G�W�J����T�jوu[�ˤ��n��E����'X�W5p�I]�';��:�6Lչ�`B.�X4��M�>����Q��I�U)�;�#�^V{�T�&�z��l�6�o��St�ݜ,WY�B����2~sK��A���`����3^,۹�d���i������(�B��]��(U����fb���ǅM�2%( Y�����o���(+��y���n���>�@G��A�E��+�c�~�%힚�/�I�WGf�]�M�n�S)ނh��9�
F��!8V���	����%+z��g�0�UИt���.��d9uZV�w�r�X��<B��K�c�d	���@�t���9u�<2b��6��/���;*�W�;?]xq]c�*X�����I��z���p�n��3��޷1Ɇv���|U��S�J�܎���L�c((uݦ8������x�)���W����G�X[,��v�E|t��	��4\���_�� ��O��y�n�&^����Q�*3C���r�<<r�|�e�������������/L�7��_0�Fрo&������ݖ��T��Ra��M����x�2�,cO7oC����,����b�W��"|*D�r~%��PR͚J���`�`��=w7w���P��M�7�G�QH���x߇ �V#�T�̨�6Qo�%܊����������Z'������N����_FR��<��t̉-�)���q��6���z�DН==y���'�?��l�/�_ǀ|
�>�K䑲*\�r�wз��P�|��4�ήy�6f�V���dg̸e�����֩v��ò���u^�L	�q�㾹#��Y�[��G�x��*{i�������^��֍�S�t:� �P��B�e��.|dp��d�%����oZ���:8���z�!����'�I��/��c���纃N���}�U_R� 78�~5�q%��P�sh}_�ЋB��h/�Fw�����o~��yZ��,�����O���R��İ'e�7���c:��������׆�9��ÐG��
_^�̯҇2���fJ���1��aq�&�]@+�=��⠥�����C3�k�.5�3�  �w7�qµ�3+��,�spP��/ud}�3�y7j?�K�ö�����M��0�]>ڐ���\S���κ�L]��A̓�Y>�1� �Չ��¸Z���zL�oQ�,��#��2?`_v��mi耐Ȁ��o�y�5ٮl��_����J��6:�C�7Isz�k�SJ�;��;����j%��5��:z�Oj��|����w�4�C�	��W���K���q�����6 ���b��/1�2���o����&�����dX����)Gp��_�T܆��i=�Í4�	N�!/�?�c�733�@\%.�VjA~�G���M�.v�0�(�t\:ȯT�d���E�*���]3�I yPbj���*g�#���8{�j�� �1*�ے~2��~�����+͌�j�=F���ebj���ۓ�
LH���!n��گ(o���)�"�Z�	�m`��������x{� �0�ep�E���z&>Z0��5}��O@�ߐPN ,�-*�&�q�L ?wJ�PD��Fv��b���nO�Q�@����Ƨچ�"gJ��O7��Q�`M7�"N�B�H�^�|��ʫ�v�!i���G��g,����Qޟ��-��ﮋy��x,Z��\��������1�U�}���$���=A^�;���ʊ�Jz��X9
f>�S�v�'H�XŖX-��z��Tw-�\����Y��$�##�̊k^�hWz�|�ۋ�F-t̡���"Z,�����9�N@2���ج�)WG�� �>ᒭ�?֮�u����8b]����1���Ty��2i����A�t9R�^��k��\���EFxþ�z*�	�^�}��&�	S���2�o�G8,T[(�c�˻�H
d�o�H��) �+�x�%٦���4W�!$�oa"�\�s2ۺ7J;|�N}.�Ӎ�Ʒ����C%G���^w���;�ڊK��pq�񱓭�?r�WHmK��FX�c\�e5+�^
h9h�2�X�[�.Y��h��F�*H/��GY/�%���,�mߧ������G��k/
�$$��Vq:�ze����,��Au����P��΢�H�6 �pԺ��cDCU��q|I�����Æ�%1����&�3�|h2�����=)S&�5 ��q�O(081g�j��ʆY1"*�a���4�	�9WvRbE�BDxI3o�A��P\�U\[�حy���l�O#��,�$i�Յh/�ԋ�����q�d�f!EQT�gq�����L�a��S�͟+(�?� ��K�2�����S]�Y|M!?:A�ND�m�#D���UαX�2"��GA�mz�*�`���J��5�0M
��:b�qT�][P�E���}����4����l����5UW0RҲ$�J��%��";%Z]�d�(+R����l��!Y�� !ϴ���NlnX�iM�5Ҡ�Y����o�1w�8�&����}��,��&�#�1/���O+o��5"�Z�R+�J����/%H��E�Ø$��W:N>�<t���l��Z$i������y1]R������_�%�E� �� S]ٚ�Ѱ8���@�Ӻ����f�v�F0�:�����Lz9+��+���d���_��NÃZ�*z�"��/8�G٭�W��tZVl���6����NQ����;'���)�����i߈&]v�ܽ��K�����R�"�py�i����M>���D�����"��r�)��-�E�r��{s@W��X�0V\�x�y��^~�6�1i?���PH�����c�o���rQ*�`���.�|_]r��_G�M�h����6��q�\�gT��IY��ךkq�mс*<K�@k� ۪��i���yD��f�-�6�_Q��C^�5�x�`@��c�i�R���?�sd���������m�y[�K2����))��r����p�,P��N�8)Wzux�܇�S�l0Đd=3)��E]"��潃$�I�bF����r���-�f(t��������y�mϱ���/��+,�W��I���c�YY��h��_ڧ3j��2���ôޢ�R�����I,�8z.��u�Y쳌xg�|ph�Q�9���d�WԘ�N.� ���	���θ���#�CJl<Z�[*���wu��^�xNB�x�9�MC�'��z�G�� l�����~g�5� |�"I$�'N�ֱU����|bV`�;'�����+גּ!�N��:��\��V�9��ĀQ⒦����.q|���S:��� �M.����vں�X\�H)ݫ:�MÇ�<��*jV�^�[���D�]RE���)Si�<˾w-�v�V�<�ÖF�!���q���#S3�O��p�&$*o��^���$b�]�����3�Z%}�_���7���E R�HF������5\�#���$Y͖���o�[[@�������rPm�����DN��޸;���z�S%�-)<�8�.�@m���,U�K�}�<#:[c������&\>+�EJyXi�k����x��2�,k]9:W��ݕtlp���%K�Su�r�@m�xg�1M,/e-�1H�����5��j<(/v��/�	k�� �	f�:��a��r<�:�+�/�T m�I�:V̇�Œ�����yF��H�@�{�����y���m��ab�T���P��wL�PR�ʘ�ٱ@�Q��h��������.4C=��3��I5%���Q���>���;�o��>��Q�ۖ�N�����I�>��9�n^he�x�Wㅆ5��e{�Qˇ:�U[ɂ��м�z0��)��M'L�HF�p4T�b�q����˜:� ���@�����ṢP� ���40�3{)Y;�|��x�1U&�Ѣ�����O��uU�D�N�w�ݴ�*��.3���4A��������\�
Zz��h�+����?���O���s��3v^���1�<���X���y	�ğ�I�+���A}��B��=z�(rA�Z(�/���$��oiqڑ����9�.�&!?����l4B[����^�qf��j_ ���F��5�I��[X��
���j
N0�����Y̍!u93C���2`n�o5Lg��>�v~͚��S\�C�Ǳ%�	�C�΀ �ͼe�,�2��j�u�@�KG{		 ���P�R�}�3�&���DU�?���?.
&P�f�YS��w9PI�5隶ff#�Q0��� T��k+IF�<���q�5�$2�}<�UE�ӿ�] C�κ��[�m�p�t���i�*<t�������y��~�Z��1��4����"|oGB������v� �ۻ�W"��i�Pj ƹ�F0�'�+S�v��ڟZ����2�q����o��P�� 	je>ց��he��&w�<�i[#Z攖��y>G�����l�ή�~k�L��Q*�H^_V��$xőM�@>%�9nBo���?iQ��1���J�/�ebGg�!����M���F�(\\���	������[�f���ܰF+��KYˊ��?,sW��ǎ���jx"�	v��<�X��"�ɏ���i��᷸�"g�� �P�cTlӯ��޷� ��U�1�qa~�m���P9w���e�X�6�B���\�ᣗv�7��Fl�6��ܒ�[��H�)���X�qر'a=���+y'M��(��������Ӗ��ٶ��j���M��U�9C���4���&�g�N`:9�YL�a=��iF7�xu�����ߒyc��'���T�y��1����@n��A-��������4/Ɓ6�^�Gd�1yH�&^���&td7�bҾ��Ğ��!1ؽr �u��B�� 9�!ܟ�1�Z(Xk��oϓ����}�a
�~�У_��숙��J�o��XOj�I���;I�R���J-A�0��R��~�ucmP�1sxdē]����pȯ�� �*�
:j��'�D4 V�P����{�h�)(��KU����)�x.`����4�j�.E��~��}3��?,�e9	��с���!�����C�a����+�&Hy��Ft�-C�t��P}�`�j���4��)��6 =�]���@Fk_Dot����~Qщe�$����Y
����C�V�j" @g��6�g�� �ϟڔm����,i��u�uU�|6s$�!��4E�e������\BQ,UF�kZh��Iȋ�e��V��[���z�?�p�K!fTB�QM}I#�͑ {�\��V�o��/���`�×����N��l@�*�$��I�N1�?�j;���:�mՑx��0������r�a5�^rG�nN:���vaf$D���𠯳 $�b�����軱J��Mz���k��1_t�K�,L5;	%�����J%��-nB�#Be�&�mH&��|ſr�"�~��`�P:��%���P�1�uK%IF����Ѳo�Q����|ﳋ@rEh�+i@:���ڐ�����$c�\X¯�mK�`�3{@��������|��3��(+HLh�	2Z�uѕ����˵�1��������c�_��᳘ �oB��:sO�V��|A��f{�p��)�0��b"����h���@$�*]$�K>����1x��o���&�������FV_ʗ\Y�s�WM�:����������PAV^����A�h�Qd�җ4�(��X��e!�H	G9�"ܔ�k��cV�ٟ�ټ�{�F��5E}S�`�6X��O�W�>!s�s��ϋ�/F~B��,ˣHו( F�V��&"iɞ4�qV��@�{�른��G�Q��H&����;mq_�q.��4{���_>�cI�G��ȱ�M����S��_��I��8M;�w�%*J�(��R5�'4�l�j� ��u�	H�o�B�G��"_S��ЅQ�,ih��_Ǆ	i���[t�����:��M���v�U%=%��F�$�DɘF	/�V�bB��m���$���[h
�e�=� ���w	 @A�y&��PWH����ˆ���A���I5����z��u�Q���{��sߩ���ئa~�:���V¸��0���w�"N��
֋��q]�4�Җ�%�����'�f�ڟ5��.7�g���|f�"�˛���U��=�]�iVA�A�w��B9��]�]��@����#�'��$�)-�h���..w�rc܉^�c�2�u�DV���&3ud9|.XD��)uUWq7�\��,v�]Hxk�����
�6LOІ�LZ&���*\�`bW���csF"�^]�<oTb�t?��qƊF�M��#q��?!B��
�YU=q�`��WǶ�p���82X��Ƒ��}
@
�ݿ%sգV�;�EpiT`�*B�o�V7��Sc�3����}��:�fsd����TJ3�&�6��S+�UL����"0Cl[��ͮ:�{�Q%��:���h�sڳq��}��t�gB#����X��4�7��.�J�]u`��(!ݶ #j��	�G9��� �!`�w-c&�N�{D9K��%Ac��Y�`���p>� �+���6D�[��.`.�Bű�g�=7����p�a�4a�xr�B+�DN6S!��F�a��Z�JH�X�L�sKací���R5��ǎ�4���	b�W��#6.Ȏ�@T��R$�KmDt��|�wj�'��MHȘU��H�֐�B��T?hZfw/�K�n����sU���16��{�i/��ui�3I��^���/��
���+c�6���,�B� �͞��i<r�W��`!v�t�:X �7�<2R��Tȗ�DcU����+Q,g�4z�����exA*���P�*#D�y1{��
4u�6֤ѽ^�)����~;!͙�������턒m��An�^�M���V!�J3fg�MtY�L�%W���&��[�j>�AN^_3��im�W���I,�[l�o
�NvS��s:�X(�&\���]\!{Ȁ�����!i����-��X�����SGu�����(�n�G�߄[Q��w��M� ��	��x܇����VDj�ߍڨ��4Z��{"	MzfC��v�j�3W�_@�����R\K_�~b��!��NLk=�Ϛ����[|R��˽��%��X��X�6���}q=���r�,J%(b�<��{C?��=�ج�L��DƋZ���C�����������g��7c����etW�����ڊ�B��8z-��nR�_QPc��n�lJ2�y�xz0NbH�*
�
�a'RNZs+�m��3��&V���D �'�����G��pD{�(��u�\G#��~���]R%q	�S0@ւ��r�'t�ڜm�i������#o���-E�zu�c��[�V��a�[.ؕH%�*]�8w�s�&a�������]5�\�(Ï�16�=�o%�A��e�H���C��&��{x-sN��b8Y���H�r��7J��� �5X�8��9E���^���r7��Z���\h g�/V��+��U�kJ��L&��Ho���ZG�1�@�3=E��T�;8k���˲M��(���ꌖ��+�H{�>ܰ+}�}��q˥j�}��2�T+��;e��녩p�~�7�1R���-��+t�1�%4<�2^&�/	��O�`9�?�������l#����㭻& H�`�_��z�%d���O���]n��`�Ó8	$�����������z[�8{��#��~�@n_���D�h#��V�y�ȣ}}�up�h6S�b���g� %M��
a�3�`\���:�>;�9O��KP,k��{Z�)	�~j»�Q�C����Ҟ�?Üfz�J�
/Q�BD~^E�u;��K�֬s ��B�����"�M~x��/��re�ޣ���S|?�Mܐ���Q��M���ZO�TI�	5� �i,��W��(Q[�/�
qb9��K��s�_����E�@��C[į�0ĕ�g�E�gQ*�,P]��'.>z����9���H>u9mm(���?�E�!�����U����Y<������ %�)ظ��_�a�� �݁!4+�{�r����-���X�Q�Cg�D���P�땒�������I`���!i�.�����0�n��ٞ���s�أ�_`b��GM�U�HX�������tLJ�eĤ���O�l-v	|O�E<�@���g���D�ʞ/Z�x��F����T��{�>�ĚM˶'�  X2����T?��[ Z��-\�)�1Xc��j5��g�.麭�a� d���xփi�g{\/�P̳N�MoV�N���9����Xa4�*j�6a{}��,7&�,��x������1-&��	n*~�HR/����?;��/HF�];����pL=b-<z
(�,ࣕ,�Vŭ�㌭~��i�'��Ռ��L���	2�x;R�vY�a�{��v��Nm��'���Y#!+�)���ow�i0�/���� �r�I7V#���2�n�7M�F�8'愼��Μ�R�Fa<X�	7`;�z������l�N��;{�� ��ߒ�X�o�xn�۹�I������;:�bZ��VCV�����x�'@D\?�$�u?
'��waNT%w��&����X{e��h�D2�֙�L�d���=��*-�Ѣ���\��>�Dj(8�2���Y6R����#2Q��z"�e�����ȰHq�|N� �s�j��}���v���� ���RG {Kf�(�$G��`�Α��7�4��C��c��R[�dլA,�h�ZO*�p�����TP����Tԙ�i��k�X��g��J�z!���C�����p���]h}E� Q��s�}�񡦖73�P��챋v�~�����n�����bր!ʕ���ů��>�!��v�v<�ZKM��2������΄�`�S�,�����d�ca1�C}���(��C�W%M���������3��>����?�?0eٓ��F��b�ZL�Q���v$���&<Q�>o��Cgșh�\��6� F�Ð#���8�é#N������Q���&C�8ҽ�fD�@�e����`��1��M��k >86���1��ͥ�XJL߈�/�&1;K(3����4��]G�R��7X�2�Ad�-s��otHC�K/�*;��v�c�d
BI�o����Q�$.V��'�$?#��͎g�����Z�p�].K.^����g�6^��3x�|:���$xk�1�Z4ɺ�#�R;{���Zr�Jň�r��˧Q�������n(b��Rns��H���48�b�,W���k:��Z�/L<]���Q������}M�Q]��ǘ�8�����d��8J��1x��U��*J�=d~���&�NV�;���U�^�]M�gQ��LF�:�]�=%}`��wK����(�Q�+BS�6�ۆ�))�3�8<׎Cm���r��{�9�b���ʅ���H�Pѻh���m�c�Wf�1i�_�Ppl�C�G�3��H��h�������".�R}��W ��4Xb`6�u��S49쉦�s�ӯ]P��m�HY��]��K,},0�`�dx1�e������OI���$炙 �ծ�Eyb�c�<0X�t�x]_�H�r�l{ُUq�D�j�N�>F�I1�w��2�oxYe��̑=x ���0����B[�#;U�yXrRCU�I�ýP1�o�d��1[����3wbW�QF��ns��y�3N�:�-�}�@>���~�|"n=@�ք����pZq�_~�*`��
��D޷����'�k9��Ҟ߻[����h$ch��,R'�`�`�{�QhA{:���g�{�S�a�*p��60�!oh���	Z����=��*B;.]�����8)3�����QU�:bn�dc���Su�>Y�S�39�]{� NTi�5�'�{Z:�.��Y�+q���Қ@���N����-K��,'�&#*D��͟�P��� G�T��etZ��	��7�m�� � ��rP�c�GL�{�(Ja@�¡���<����pQ��>8ɫ��(#ߚ|�������h��_�
�7"[/i[��.GwёFoP��J��_c|\�q��m���GR��5C*	6��g�d�����'��}�+b*��L�2��k} �8��:əbov��z�>�S&�<��[nCͻz��\Sff-{$�縰X*���t�������Q9������a����v�k��$>@6^&t�V�,nV1=��Lˀe�x;3�rr�����Gۃ-����!�E9}UJ����E�i5^3.�,ݞ�����003!	 /=)���t	Zw��i��K�QQ:���;���9�Y�Z��;=,��y��A_Jg�������#�Hy�xK��s0����Bၟ<�ʥ�[`�:�v35��PA�byeLv�~��ī$m���|����v}I��%��~�p���j�t凧��ޠ�A���ai�i�+�����ı��6]t��:̦g�+�S�Sr�c��Q���� D�:8v75��vѧ�\@۔ǳ4�&FѶ��@?��+�̲/������ˌj8�j��'����7��g���c|��;6����Z���*ʨ�&Uc��N�|���4P��X��`] ��4A%_�tH^����Y�m
k�ҋ�z��ۗP�f�=c�F�}jD|*�+1�U�m"��3H��:��_{G��Au�9O�u܄���r�"���`��e��OjA��Npi�UV��N�h�8�V�0�Q�,p���~�+����ɩ)X�'��' ����Y'����Ap���9]�����i��4����{��~����Q��g�E��}Bv[-�A�D�L�vQt�P~qZ1�<��%�غ�k,z��8+�2̟U��?�*��GE�����q�n��/X���O0�F�xG�ѷ�d~	�(�\�k�=�������|$/J��>�\��s�å��l5ۭ�%�Թ�{�3�L.�i������`�CQ�3�t�VKy�p��V)M79،֙�z't4����W�Jj{3�7�e?<b��P����F�BR�̆	��˖�!��?G�Þn�<�a�9o�A҃�u��X N��1 >]�|Y���}����
r�ݾ�8��?1%��w�61���
p��u��o���#u��Gf��K��ޚ0�͡�P���fy�Y��������V:e;9�r�,�9��J`��-L����M{|B�̏Y9t5N�>)��}�+m���)�m���jNM��n��'�7a�f�o���-��/��f��Α;�B�04�+��{�9��n`-�n�{����1$G�T��Ѽ�Y�'���**α�Χ0ehێ]O'�����9E-�D�Q�y�qG4h�j��	e{b~��m��Q�L��W�'ardǞ����btщd����h;c�/_V�b�kD�;�I+r��U0���c[����?D�&F�n-�"�l�s8�.4ԃ(N�klP���	����"z��y�w�3Ο�L�6
a���!/4AuM���s+��gZ�ֆ���K~����)�G�!�1�ёW�;���t���?��yaq�w�;�6����k�jb"i�!�q���8���uٞ��5��ժoc�	%0]�3Fe?z��=lF������x�����w��U�f-'�e7�9*4��
��ӫe tӒ�e�����Z�:� ��s�ʽ�l��=��M�d�v�q�3Z'�����I�H���dF����q��&vJ�tu?�w����sf2�9j�69 ���B�m*<	B"��РH��VӁ4S�;��A��3���c���KNd��X�\����<Of:�<~2dJg/US��O�3�^�w�����^���)�
�9���a1kC�50��ph������/:@��	�	�0��ZoJ�vY�B�#�F��K �v����?� ,���wQX�N'��fj��9��uh�W�(�{���P��>�g@\$R7��E��Q�G<UjUlӉ.e����0�t}��+J7�>n�V9F��l'�q�m���ݑx`��/6Ľ�R �eಠ�1����$��{�w�-!0L��tø�V��M�d%ݫp�U�`.����hL U��&ډ?!K;�Z��3��p�x�����{����.�x�y��a9����b���<�`����;�$z�٫�<R�C����h%����)D,}���$�+*��ή����Y���$��j�Ó�J0|�H=Y�P���>
t�Bp\�;L$`�x�-���Y��$☎�>�Df���^��[�uw0dGhP��q�z�$ݎ�{�Mxw=`�rTى��M���
u9;�Z�oK[�BZM&�6����O�S�ڞ|6�.��"$‱sz���u?!��y�1�uɾ�s"=vB�ɚ�5²�{��j�'A���h�L)�kH��!��i!�2��źO����޶@��ؗ������l�)7�=�ѷ�r�]!�D!����.��o��se���{!�M5��'�gi#�י�{��j���L�j)�3G��e�DcZS1j��i�>]	>N��9�il�b@d?�@w��o�i`�Kte�yD�U�,}4@������r�gb�>�3GUm��{�M
]*���\p��\�d��u����L}��?�&�����Nr��1������X�(h8Hĵ����o�n��¦]טԁ��-E�{�g:�-�מ"S���Nυ㢇�	�.�L!����%P[��cy=����x=��ШI#��UQ�ߑ\��,,P2M����2 3�t�@|�I�?,��nB|W�U�1X:c�U����n�aV��dj�2KA�#Xs/A��0��&Ϻ,��\^�ǁ�5I�g��������63s�����h �}��c%�B,<�G����u��b�h I���"��V�khI������7Vqհ�����o�&�NZ3����E�����t�9��bx׽*b��~F��������e5��K@R���[�B]�~��.���h��}�K;����N�W�g��9�E"�̘HVx��
���� ��Z��w����=5C��1%*��ش�/�_ϗ������j�X xጢ�s�4�a6ϣ¦ra���v�̉{|h*��iL�~�J��F�g"o�8����Q���s"��=�N���O�����8�����?8"�⇐@�_���S�n:v���&�SU�k�r{���L��W��������Q���H2��(���W��
xߠ�������1�l� O�rӮzN��0g6�IRC��(��
�g�[ 	��ǰ�X�[�n�ZђP!���E�Ó���;^�rKh�E�~�\��]��� �X��f��v3Yި߁�r�N4��r�	b3�����EzDV�� n:Px�^�J���̫w��DH���&�����%4�=lo��0`VMV-.�E�b��.AMzZ���3��j��hnk��+sƣl���O@.��Y����aIKC�s�NHU�x�'@�^P��L�ϤK��Q�Y�33�޳MѶ��R�l$�/�Q�+ ��ծ�'���V4�0�fl�/��C�#k���{�^�� �yx7��>���_J��eN���w���&+_�݋�?��_�Ov��1�|�`���R�G�� nrŞ�A�8��͕^@;
�w�+&v{��mdKP�X�u @p"ۦ��$jo��50�{�v��A��fB�J`MҴ|�'�nG�8��#�!g�2P��8�M��Wy�:	U�jYZ�v�5rmV�݀s��	>̺������6���7���n��=�h��h����a�l9�����ɕ��<&�52	���0M�SP���C��4p+��[�G/ӂ�����>Q�������n�A|FF�`~k(o���8`|��]�9�����4r*�]��|f��TZ�I~���EG|�A.������C�7h(R�آ�F6�l��`�B��h��(O���s���\�H��T�}�r-l�����R4��Ђ\L>$}H7kC���`�����c}Y��N�D��`>�:I�BG-�PcP%��쳴�^�Q�z'J*1����=PZ!9g��_��#�O�8��:�)���
�o�=�?�'N���H���DW��䨅��1�I����&&��躹��ȯC��J�q�f��YVAhqcugrI�=W��r�y�4�|��:�}'�}��9��{���u�DwBf_ٸRy���2���O?�hD��c�l8�p���䉭0�hs5��������e�r�(����aNt-)M����<ɇ
G�;rx�.R,���;J\��aMLԓ�x��D���Xђ$WdPGmEdR3J����{��U?�� O�����jM�f�U�Ÿ���&��񅙭���U���QA���5��m�JB�2I����!G�O�Ny�Ɣ�"AVQ�M��m�(�R�W������K+ye��.�S��Ͼ�M݄��ɴ+ތ'q�9X�>`�#�K���'�K�A��%/�WS'�p̪F���H���z�|���H>���vۙ�FjƵC����R5)M$����fRgc�W߁�8WN>3uU-�ڋ�3�:���H|�*Cv�h�"���q����C	.�������♙�].f,{��~�j����x�\%)�r�u��?7�Tj�f|�?���˥j!�}�˂�M<ĖE��@ퟎc�����aV��<��U�g'��xX�[��5s&����YDȺLʺ:i�����M�����.d���\�����э�����W<��(4;���k{[^,��,B]D��V��"�f�Te̯����ħ�O��]6Pڒ�}����ѹ�� c+R$G��,��E�]�A���h �d�)�[.A����ph��<q!�{ f$zK2�����v+�ʒ�y[$G��I��S��W����l�wk�x���]p݆~/�, S�w�J�]P��W��8��s}�N�3!.oZ��~~�U%���\�"�N9�9��0_�J�ȳ��r!OVI�n^|��?��;� \Ñ���p��.��q����0!M���eцb���(B2/i��^s��_����U�	#y�/�Ga^J1��A�C�6h�+-�8M4�x%��܇���Pmj�j����
��u��d]B��bD%lۍ||�$%<��iF>���Z�\*���F��ƶ��t^�3�@��� J,�Wj�I�z�L��?��L��m#��;!����r�i�G^��ڔ�;d���H��8Ҿٱe���f-
ӞKtk)SpG\�G�����i]j1�����(���r�'��Ū����n��IPppظ9n��F�R;�7��	s���m��2<7��W�nӷ�`ח��t
�eZYj �'+Y]
1�ĸh��l�)�}��۬揠(+�0�QФ�R�,w`�l�پ�D�������N����l����n�&=m_5�=�qR,B:��� VI\Ki��c��ףF��(]�K��)<[�<��,��M���C\�v�m�;��P��y��Z��3��~=��k��Jɽ�<��R-��^F3��Fa���Q\��X{��e
�sD�}��n��#�)�wNv��<xևB���f������	BƐ�?�_ܽ����,H1{��8�5ovz��a��Uq�H^��
��/DK��1ƅ�$´� ��a%<�_ :�ET���&;%�+!���iV�a��׏����6j��>���Q�h��0�9f3�L��O��SЈ�^rMR*lc�jラ
<:^��C֣'a;��?��x���OO�/����+���[��-:l|���;�^��5Ջ��گ�!P��-����q�Y�t��BYzVԃ7���J����M���F��@!臧AŽ���υ��7���`�m��-���m�e���A5��Ί?|���������t��Hn�_���E�y�[��Sk�i�着�>*{V���z�Z�&�� ��7\��ۻ�,]p�FA��,�t����hm�2>@?I���HQ�j�N�b����uk�Sw�Ɣ�k��'���f ��T�e��ߌ?
�lVH�0o뭰���Gw#�Щ4�0��a�����:�����׏3�!n�t�����b�icL�5��=No�<��`U�����RذX-N��!�̲\�^�3[ �z�����<��ʺ��G�p�A�7�ޕt���@�NY蒢Lv���Vܖ�7ه�ρ�ӕC�*��j�pm)���~��8�����:��;օ�|���Z�L˕��A��\P�Ԩ�8�ɛ��p!����eѪ���iͤ��#I��M)D�ż���G���a*�H�):5+oME]}�Z[�^!M���J��(��>� 
$�������n�׉e��p獐�q;\2�9�oM;"�/�q��}E�RA_h���'e������
g�R��L.�������|u8~��(��Y�X��3p��k�J_�P���^g�
H�����:ZY>畇�.��cz�68�Y�&	i(�/H�c�ʙ�or�⇍'��j)at��۶QnDDxAss�Jd�!1�{CMc��ɟ$/�ՀP�����#��T��I����aQ�U�l�����������;�ZM9�����6�{�p"�m<�X��0rﬄ�Ħɐ=z6�Z�t,���t37~��[��q�i�{O�`bQ
�Y�zswy��|��mԻZ�:��|���CJ��׹�sE�뎆�����Æ��*�H�8Z��R��Y����)�XL]�� j)�ːrP�rr{J��Mea�v`�/$�~��#��X]��Vz��-���n��/(�+_�87�V�`5
����pra��4_���xn@����٘��s�ʢa@�IqU��7JŉgI�q��Rm��A�tx����g���8�Y#'�lV�����p���b�L�Y�;Ć��v�+�E�Ҩm��͍��h�=k�����kQ �j�_c��w�3౩F2T�J���ٍ��A],�O���0���T<�b⵲4R�_4B��\xH��#�"-�����`��a�Wi����0���BϮ+3	�_S!�.{r��ZH��z�%D���Ӽ$j��M����S$�l�r��A#zŚ��?=��56kB9h�]˂T�>�Z��%F'f����+�{%h-��V��^EVDmZU�@.��2IHR��g�y>�$����3�3S��{�'":\M���`�:���N3��t]�4yӝ��
�sl�=��iw]T���s�h+�Q�5M��QI�}`ۨ�5�c���Y����(W3�ފ�b��|fڠ�G���#9Q�T�u=����Wٺ�}H�04"�յ ſ�U���1�D��퐟RG_[8M����g�9ڕTM1*�b��k�~�8-�!:g\��vƦ;����9?��!������k�(E���g�B���2�zc�_<�#��uF���;�\���~[S fuu	M	�Mw|`8�����P��a��
3�l��V������]��V	|��v�/3�P���'��V,"s���c�����yK9ّ�<t{D�̽K�z�\
!���^c|&��V��i ��fv*I�����}�l�4����U�FΪ�-�\��1���ч^�2�D�_��,J�bÎ�������C��c�C��Rr6��{sɪ�����F�L�"<�R0h&��d�Nb�|��oz$�M��%��NT�Jy�n�
����������X2H����wt�Y��j�U�1Rh���lI�T2�<ݘ/�zY�A����ŗ����q����vn�"4�O�B��ld���s�\�aS��`�P- ��_j�۩k!d�8�(�d�!K�\����M��h���<�x�௞.��X�.�\o�a���.��.��hK`w f�c�.}B���Ur��MYu�y���;8iҫ��2^�#Ӗf~��'�����l��������RDr��F�=��)o���<е�H�*Z؎tV����(����n�*٤l�^Q;�IR��v�����Ȭi1�5��g'ҌQ0Lz�y^��<�oޯ3āCad��~(x��O��f}K�]�����j]�f�P1�&�@9�$����k	�
MiA����eҙ�o)ţ|nxنW��#�Ց"vW��H�$�{>W	Y��������n'u�*Mб�F�����2vM3{<����]֛�z-�1��y	���-`o���|�ߎ��q�r�����DT��^�C情��z#?+)�^ !)E��.zQ��S�e��(�g����XM�y@.���k)�$X�ŷ�^E�(�*�fc���l$v|Au�5�f1�[1�f.�/��F�'��J�\
򱔁����Eדrn��d#����G�b�j��'!Y��Kb���Ch�Kx�T3������?�r����$��oR\ �H���i�,�����
5��+j'ߎ(��F�ު�ء|cr^q���P�8�u!�|�w��YM��ŧ_�\扉/+�d�^b�|���&0�����Ark��gm�reE��o��R�q�UhWĔ�@�`�fk�E��u����I�Jf*c�EM����ai�]�l4/[��p:�w�.&M�K~���F#r�Ō�2+�������\�2�qj���`a����x�DN�4'<�{7ڟ��
�SZ�\)&ӂ/E��x<ar�|/W( ��
��v�&��O-��>�c��n� cl�ڔ��
Y���9V���@,V���R5<��j��H��a�Jv�YqTd|�ڊ{�`13=�#@��笳M!x�['�����GC���΄Q�7�ؤ�!�"ffA�?� �A�ya��P*��e�'N���3,*Pbf�EOݗ��3T��B�]Z[	�����Bi�+�|%�r\�i|�3u�������Π���B�l��؊�?s�>�R	�
ո"�����&׈St�[ �G۴�%y���B�pW�@r2/N"�F̚3���kM�h��ItO��-���'r��\.D�t�����Oe(N�� C��)s�Xqu<�8���X_������M]�R��,�T�]A�P����W=ւ��Z��C��4Z"�(��E���e�(�u¥!����D��
H}Rԍ��<�ҖYգ*�N�\*��aZ����`eeh�P\�=�q1|�ib�NB�9���� ���i5mV��25,��^@1�2��
S+\�=C�h�h�]i�2뼾DD���.�O%�r�m��~Vc�J[���D-=!!����'vl�	[z��K�Mޠ�t�v����v���'T@k�q��k�bK�$�$"��DLw��g$fw��oy�B���V�n�[�1.���M(K��s@�ܼ�E� ��1������0-b��,�L���8��}-�R�DJ�RU-�������C����.3ո�w{z������E;)mml��(R=kZY��3q������߭�8�k���z:�#V�d�]4����-��~���������k��W����� �M ҇{�sDv���#%�4��.������c�{�N��R�ҭ{qRL��+=1�+��;3@3|���v���g�C��t�Hx �+��� ��l�V�Y��*8��v�'�x��p6��c�W��Jt�1`S�����b�_��RlǛ,L�-W᧬���髛::���Z���j@r���|[η����J�	����"�-l�. ��!���V��@��{�`w��v?)7e�-'��3$�ʔ���C�& ���w-�bQ��r]ѿcaB�������*�z�cI�d�]<%�sϼoE�vBD��z��}��mB�h�����^�se�l�n
�J�J2r+���i�
V���!�W ںq�>H<�I�M�l�w�hCI�	��N���5{���ORz���Kt�`�*�C�N7-!�JT�I<]�����"f�E�4h��Of���%���(􊲫���	���lC۟��y�*��wZ#��� ��KG���o;.Y��N���O�
#ں�5DI�5cF0��c}(N�,*R�hKf��Q�!�9��lj��%.����<�F�tq��&}CMk�2�+ɜ���8�}Q���O(��O>�]�l�x�8}t��NՑ��a���#hi��篟�4��-���3m΃���ppʡ��]y�!�³��W���
��Ӥ�������,����8�y���z��wN�;:E"��
��*g3N(۠��Rh��]�����zu�&����p��fB0�  ��	��C{�ޢ���.o�'�.�?�@��-뚉�u�H3d>hlfA��92�h4[2TO>�wq>��)Q��#jA8����9��QT�8Jq"5 c�LJ�Tn��w�rsc�U�H��Vg�|�-kI�Xp	�\�7y��nb�t�c�Z#"��ϮJW�#ژ�\��+�����"N�����&} d	���w�7u|��{����8��.Q����A������Z<T>��ɏ3����FW��&#����\������FZ���s�l�5T���6�k4�R��e�ů���H�m�ܞ�2{�4�,��][��s.v����#i�K	=��oZvԛ����D"�\Jy�h\����1� 5h�j�g�<�*Os�?SdTG���=͍�ϰ��cK�;"Ys'�Du�66�!�L��C���[B��=R�o�����nZw��m�H"�`H���9�w����^4�8���u�L����,}�y�ᇥ�B�<������8��𖳱���Ϗ�*�AB���M�80V��W������6n��%i:�����y��#c��C��Ǽ��cE��z�4 �g�P;��,���0�E�[��{�[Ifp�%�8�-��
�`�3��"��AK��/mC���^�d�o�ʧ�c\K���L�x��W���4B��$�ޑ���$�Z}o�ȶ�ħ;Q�k8����_	;KJT� �X��鵭�\Ԍ����M�TX�����t=�V�9�0e:ie�8�&EKod��R�N����.Y���f���m��Y`AL�+���<kbs�H���v=�]�����6l*`2�R7�������b� y�`��|�5��DrOr*�o^�����2V�\����7v��Hw�e�����9��\�h����7τk��ǵ3�f�[ ��T�
�+�ļ����O�<�Ap�Ħo?���pP��y��D��Xn4*Rfg:t�!��cC�g�@�R�xG�ӳaR���Y�`����u���ƀ�Zi��NSIA�h�ִtn�	h�x���@�=�N��:)^,�2��V���#LL��yT$�B���L )������'��>5VwF��qz���a���|���S1d�Q1�F��*��@�MΏ��Q�1j�Z���k]�B-7��Y�j�c��}�8F;��:����F��H�d���*�Ǹ<�b�@��i��W�y�T��Ã����x)����/M�u!�#��O����f�Utp�3�ق[�J~)
�e<���TɿYޡ�-c;��>��8�@���y^�i)}Pm�D�e`siT	4�ة��߫�aQ!�.��=��{p�×�#ĶLMǎ��~r�)��Y��#�|��Z��߅��4��_��fs�1-:�L��Po+��V�NM!��չ#oІ�R���,*2�VO\�{Mt�E�"3oF���u󞞒k�*r���+t����l31�mÆ ����?��2 %�0'%У��o��^Y���0]Q�v����alr��ln��� W�c?k�X�����aŌ���<����c��В�BQ��	��v��KŲ���Ѵ�Wl�L%t�<���c�zc��5p����|�y{�;v��#::�A"ͱx"�?�)i��،��J�B=d{�P����Z������h�T���6��3 �f��+��k���
psKM-PS:�n�t���*G[�;�IN�k]�'Xv㨕�HK�7lNˌ��D��tG��>іx�vΞ����{B*c����]m �^[����y�]�1�����Є��㪀lk̪�v�E��P��ߥ�R~�Ӯ��݉6������xJ�01���*jp�G]���aԺ�$9b��W����r-Oۺe�����ҐEaĬ�_���Zf�0�c/�/rY�mp>D����b" 4�$�e�A}i�0Z�y�����}�5�0�Kof��F={�^�֟i�xI�RC��ENGE�W�MG0��;�0xU�������Xn[��DZ�尲�s@F�-ݙ�4� g�&�~���y�X�1�@�����\ o���٠z;��[!նc�[��s�OŇ�� ߋ��e��&��+ppN��&¶�Cī}�M5榻��{��M�n�W�yr<�%�Ҟ��__�ߤ��p�{B[��Ö����8�:s}�&��f�xF�}�3R��S�P��rY����3��r:����u~�9(�a��.^W"�qN3	g%-e��y��Z("��z�?�7�����	�]�5�鉱��Jjr��uM,�j�l���o�����oe�/^�}�#�X��LWط����Kn�t%_��Ei�	����?�æ�		K�yV��9:����c:�B��\�ȩ���5)��[Y�i\I��t����L�9U���m3��1�2_R���|��h��Q�e�/�+����Pn�_�L#&qu������-��5.�n��W�d�����\�Pz�}��l~]c9N"�f'��dê���ٵ�X��9;�oH���3a"H��m�kn�QBg����]�_}Ɖ*�KX��	�-���B�A�H�������b����?;����xM����&�B�g�X��8��DN��w�)���w�ݍ�Lފ\=�p��B����kL�3���g��r���p&�^����'�t[po�U��J�DoJ?���d�_���c���ژ��fO��W���D��P���E~Ğ8h�����CD��x�ث���Yoa�U=����+�P�_QZ�нlA)�RMmFG�������5�ҿY|��rt
��bY�ze��7� �z�$�NjX�e;��zGॺ����C��ߠpƓ���Gi�'�
��i�$���0
xxŤ��M�!D"\ôQ,�zO�4Sl_�7�4�?����?��i?�Wb'�ر���Tz(������J��f��
�^]{���A�n�w��}�E��[���Z�i���Z��E}_��B�\��$T��K@��T}��Zfp������'�4���KKޜ|qog���6(�kɁɝ����y����L�ʲ����kg&�m�;���I&�+͚���%���)o�
�aYi�ێ۔R�ĀU����/9�|�M���n9�E�A.T����4�/֪��4:ES��w��$%����."�^�nM;�}�A��IW1
�7b���Ac&��f�\:�����2BT��LwoM�+=�y�K��W=%xXI�9���b�/:�U�ͥ�-/�zw51ap�}�N�p~��_[?c}9$�oRAd��8%�ٴ�h˵N�����x*���pe�� �\a}�Տ���|� ~>�����C��qj�u9�(BI�J��s���%��u?�6�܂�l��G�Z1���I?�s�����2�H�[�S4�J���8ݚ��@�s3 (�O���!ؐ.�b�hc����7��
@0<���I�?h�M������$/������Dޞ���6r��9�bW�|yɱ��(��%�&��;��e!�a]4�D�q%�)p*���Y�A�1������:��Y7K���8Vz�+ԠC�vz�>�L�+v2�]~�g���<-	�q�G'�&�hY�BL4����g�+#�e��rƊ́���vu�Q�>iP=��/����8�T�z�$��c!!Saï��0ڏOa��D�c%t�"�4t+��~4*��}�,q_�9��臃�Wl����pj�T5ȃ�����i�4R���9q3���]��F�zد�/,c�ri�Sq�ǁ�H�!9��?�V�W�ױj�Sʕ�>�*VU �g)h�5��
:����py�/pK�F�0q�}R ���7V�c��b�/�"Љ��x���uT��,�c��P63�>Zs�&~/އbA0�L��)?�(��@��|�Hɖ@���nR�c����#�h������F�7V�JW�6�8�A f�ṣz�A�R��-|����j��	�V����ƘW��:�Y���+��%u�0}S�홇�%	����0���B���Ŭ�Z�}�Y��q��Bͪb��4`\�J��:�:T�op`�����%�I�Mګ�[��C��Z�pV!-c�	)Z ���$�y���^�W�~�`�w�#8�A
�zď&k��O�d%����Ǻ�I���S�����C��a�odI����\��5�ܽ��m�������78�)��֮�\R�p�o�pI�	�ED e��6�MV����c�8��%)q�zS�JVۇ��@��	�,`%���l���B�q��kI���e�	L|��hi	��;~0$��̏�f.���7|$ �6��o�dTpb�+�g`G� ���F���?z
��>0��ě��Xu��5�_�_r;}_'���'A�G#�H�
����yN�?�ڻ�ȣ�����V9N��������$ae!�$��?0��`*�V����8�J|�`�} �A���^�E�H)93��Hf��(8����4"yP5����[��N���b���WK\N�Y�W�NY��K����A�@S���E���%���.5~N��
R[22�F�d�%���=h������
��$j*�����Z*�T�w��,�3�e%"F���ܕ��?�Kw�P�9t)"��0��w��BT�~]_�-�%�/X�8C��"�>����y4vK��-�#����қ�$�9CN�BST��3�`��F�[�|��.����&���{����a�^J�I�2��u�0�JeI2&�ʗ!	`\�"���B�V@r�:�kx���$�'���	���T3�5�P%J�V�������@��${܎�j�1Csr~����<�(�'��/�28&�t���=aGj�{��}A��S;"�SX�~y03�K�G����C5ݔ���'I�lG�p���q4��%���W��e �g��@���W�شze�㘑2�ӷ�!ʳ��1IUc�Q�y-��ω;B����D��0Q$�c�E��&]��Ͳ%�w�� 6��j�=�yVO�j7�e�L���0��� ��x����w��C����Dl+5�#_l�i!��Q`5�$N1�g:���ʹ��0��z�v.rY��@1n���Y����eͼ�rl���Gܚl�N�3��.����@��"��W��dg��03�b��h��z�zub��p�1o6�G]�h�(�#��oRJ�v�B?0�!T9���͕-jV
��Q����P��������	�t���y4��Z|B�Ϡ�KЋ+K���m�dE��h�n��k�/�ڴo�X�?G0[�z�n�cC�Ĵ��2�˨�È��=�$9�A2�}�k���f�<e�ۉ�`;A�!�q��E�d3����C�w~_��b�xU�D�)�9�/�cVJ1%�Mqo@�Yy�x"�tr��&w�ex��2�O���N��F4F�{s���q�;:r(���d��p�җ��|�닣mx>ɾ�k�ܮ
��g�ۆ�k�d��΅Ԡl������`�NP��aI�S�PJ�"�Ȧ�^U�O�١�����5��Sյ���,�-�₿x�wG�����
D����^2o~�}�C���ҕ�$#������~`��b-��_�R����������#�E+�M���O�4�?Q��Ԝ�a�L�/~�V�������LK�B�5����zb$����׋Ml�u�`�X���ƵO�W�YX)��])�! oB}`�  OH��u�n�j]`,�Ruޫ{�(�V�~a�Vد#;��,����z�����_eg��p@.P��$-�����n�x�p��(:�żw��R���E�]�x=����xc�h��QPϘ���t
؊vvB(gӭ���bF�Xe	�����b�A\iV#uӆ�f^'�G�2�{���V�{j��/��b[7��9��u���4ON
�}����!C�X����y�%���&�u�|�l���$�ן�2�Ng�fw����s?���K��^�{_F�Q$�̈́Ӟΰ�@P� k�ϵ�9���?:e��t�F %M֑`�Q�>� /����kȝ�Ȇ6�#9���2�D����34��
��Z�&������z�^P.]����Swd����i�y��rl��sP%�1�?��x#IOd���m[�`�-��ō��$F�'�YZ�bC{�a/�`��md����]\e5��)��>�=D����'��aƢ ����I�#x��,�+�i�+���jG���5Q�H賘,|�w-�N �]����	�mV��L.�w��;!U�����z����r��@9�>#����N��c��W�#1"�oԹ��������H�_T��p@�'�e��{�{7�=냢�e\���mEtN�-O_2[��*�˄u0� Ż{���pB$���b�������F���ٔiup b��k�.��$|�b��������=��)��:�DsO}ԳU������+��F���gW�P	^�؟Yt��,c�(��&i�]`�]����e��|�"Ɯ�q�;b���p}���4��3\kp�5m�#��^**F�o�=��𽂫r���hY�u�<��_l�:��?�鐾�����83��\��W��E��m0IVu��r}��οĠ� �[�����l/K0�	� �#�*���D���.���=^��=� ����w���7�W�l:r�[{).�b`	�-*�¶
3�� VVHeV�Sӧ�%lVF�81�=�v�ˌzK��s}�^RF�~u��1�&_�h�+�p^��z�+Z���c)c�[g4=b��VÉ+F|[�,<!�t��(kk�bᬦ�
W}�"nq���G�$�}�>;�����ì�>>�s�w�r��s��OoY�����|>:m�<s���O|���.>��?T�#}��;�w�¬�Mo��cz?�Y���&fs��D�T�� ?�>ړ��-Ȱ����~�w���NQ�����5+`�		�@�=M~7�y�+	͔�=7��P6F�='�)y֋�B��-qG�8:��O�~@��#�T�(���:h:���))"����ܴ.���s�����/�ȅIV�Ռ�bJ4n���1�K�bG�X�;.���ۥWv� ���L8M�ǙڤǺ��_�'�k^��v�|�uq	��~a����J�K���y7һG��!Ժ��O�YK&��q9�o��-�f�;N��i��9�_�������9������'v�#����.,G߮��Օ������ms�B���sI�"���3b<��O�-Y�s���:Zh�<S����2Zzil���Bz�f��Y���sy����M��o����C��9I������r?#̈If�W'1	�4X8�u�x4j���1ޟ�Q��1�E�NΚ�xM����B�f�����3������Z��@!K�5��t1APp?�I�}�ಇ�E���X��cM�}�*���JCus��-�US��T�(�:W�kJ�=��aoM�O,����i\X�B���Ĵ!��cP�Ž�+�����c|��S��vG:/ۨlU��BF�˝k7`��ހ�XghpLH!Ya^N({2��\����ېw�ъC�n�a��gZ|OSU�[��6/���Z�]ԗ:�?�c�ʹ��u�BW
R���*��J�����g2O�3���Bg���O��А���
 |����p��Sz)�T|�[2'���v/)r� H�s��o����-�q�ȥ������!>8G�:����Iw��iU��#�j��!x����C��'-�1��"+��8�k��](���'��CmDҩ�-n x����\�b"�}�>����ͧ�:���e��L��ݤuP ���A�fc~��6w#΁u�a�+Xǜ�$��Hyw��G�_8�)e$�g(�����~o�b�;�� u�0�Q�� x�TAՔ!w�m!�r$9�:�:���~��<�~��%�	U�#D+����Ez4�r�Mt���di[���8��)�l�?M(V�����7��D�Gl���Wrs���\��� �P)��wU�b���Q�'_�#���)S6���*�c���x6�{N�1���S�M�b�abs���ZE�ot��<�,@�?r���jF6�}t��y����%JĄ��Q�QV)ܝ���9���=���R�����2�:�r� ��<:,:zG�	h �&� wV�(���|c��`5�O��M6�2)�F�|<��}�W/��:#3���m�'�zZґY�B7�n�%������OTkX�:��tT+�}"��T9������04d��_�D�Re�K�ICHk�h\;B�Q���As�g/˔�%�E��N�$� �9~p'R�P,���#�=��#+j`��L�x �O��罓�)�쑢�^�(�P]��4�������x	��4��56�HV޳�_�?!I���^V�4��_���2���B����K{{�HN,�Oo�EW�P�Vkd�q����ɞĐ텵߈�?e�b+c>,:�	SD�*�@�33�=�C�fq5S���ɜ�h�KC�&�=Cf�Բڛy�z���hǚ8���F�B��+^��f��������sw��q�i)Ir���m>d:W)�̙��%��1b��v!�*ńx&�)j����3A� d	1~���0��	�����v�m,ǿł�1掃ٶ��C�Y�L��f��r-t>�^9�Ց=�2[I�[E�2��2�쩪��W���*'RzX��4X�� XJLtN:��)L�x���j����翁��j�6�Na�k��/E ������+Fz�0Tܱpp��%(|��ιU�$<{��"݆��BO�N$��g%=�6RW���O�9�?+�`-/����]hd�G~c�g����p"���h��*[e�Hsf'*xP,�Ό���Ż�A�KeN���<s�DOV.ɺ :��Z��5(���_%~0A6<���o{�e`��uj�R�����p���y�4�2b;�-���Z���EOf��z��e���V�*�,>�-����.���������l���G���b/;�d8^�),�Xnz�;M��������C��8���E�2X �� �F�0��U�&�Ыc���_!>W��HHR����x�ꝱY���{�k9_7�j���*E*Tu��[�Cv��Z�wǗ��]ۇ�I��4�Q�P��k��x���i�O���I&�oo�^���;�1c+������H���7G�!����pn��,昹����S���~����۞M�qǷ�h*�)z�խ�Ո��X(�s��
�\���m#F��K�"���G{�p�Q�Y���8�7y@�ڜ�[G�\pP�3?�잧���3���j��"�$�
2�x4n�8u@ˉ�)Κ0��J�I��}�q���{{� �o��^]��j��ukкK���0�ȶ�KZ�3%	s�q�c@�x����@�}U��L=r����s�����LT+;KwH&�	�P���C�;/���B:�����,��&#���k���+��J��w:7�f�����)�;�c@C�}���%���{_��X�|���qk�;�q��q8�в�u�km��,�>��r�+�@74!}G�I ���LK�/9bF|H�s���1���0�Ɗ�Z�y6�S�2d͈�	���z�#�/�@jy��EP���>�D;HՏ�7�Ű�锗X%*d��%���~zw�-�BG��D���'w��c�Z�۠6�=^2l7��r������.c����3%������Ĩ$M�j��l��+���&��]���t��9+7$/,`�����uˠ�_X	�,i�6>�'�\L��ǒ!Y���oسW`@z���U�����k�W�P@��zz���r��8�M�{���ɪ�x�R�<�zcP5gf�e~V��:Z[-�U��G'�&��؄�ݱ���-��m�53�0�������(��)z�m�.�z����U�R6�ú
�ٹ����r�[M4�`��~�3��A����������)l��
�G�Q�g�D0�z�6]k�+��D�Y 4	e�}�ZfK"冴M�seQ��CQ���LV���K�e�Z�ބ���D ����6�!���T}�1!e3�)��ՁJ������#�I5��s���B�qd>U �$3�{]?(�\�7�2��ˋ�,��A���t�=�q�%ozu�=�Ī�es~���F�-:}՟g�L�k�~�G�2�裰N��ύ��"�Q���2�����^b.؂v��Όˬ~�x��񁯬q��D�{
QClJ�8$�5zNs���6S���摁9Fе�u�׷�y��9HGueJ'�iW�b���,4]��Rfa`W����X6�C�A!�芼&{7,f���m �'�"�R1s>�S;�!U�`���E�aK)D�편=�j?��^Nt��5�����,?�������^��k{6_cD�������-uJ�z��4��@hU��z��,ǋ�D�����m��S�~M�:��v���x����P�R�N����*Ri�6G�s��py��>l_7���nL����F����!Q�����^���F:U�8�S܀��ݛ_����)��z\3��a0��V�ҙ����i�f(-�'�g����1�Λ�O�!9Ɵ�͕A4�[�/qhY2�ҋ�{�
d
3s�pi�@�m:�i?T�y,�$�f�=L��� (ajPs��`��#M*8n����������AG1���!ն��v�(G[(P�<:b�Ӈ8�]n��k��X���'S*=�l;\��-I�� 	VY�$k����� ��~�?��F�"��?�#c�ƕ�3G	P�z,��tR�I�F���ň�#���-k��2 �%/����,fZl �[a�	�x��A�����<��2,��^����x�?�
�[X�ޅP��s�pK(�-�IIdM┯pWo�5
�B6�*J���v��=��n��qèW�H�/��aߜ��Dm���ά.�F�ݞt����w��zJ R�M���~�ͱ�f��B��}��ޛ�ڈJ@4��[�+(�J	��y<���S��QІȓ���^�3�ϴ�&�dg�3V�-7ԩBPF���
��;�����%�&<J<~P�~��#~�δ^���S�Ѽ:�	�t�8�^Ï�����c�:���!�X���e�L���t����Q�#���[������9�38�f ��QzI���
���x��#V8�`~���KGrmN[�P���>���-el��?������0f��t�>�ko�f*�v�se�5c�]E���,Y=�eKb)3���
���V���T�r����4��H�-��c�BD0�p���O��R��:@��Tl�u�=���ٱÚh`WC�	u�vM���.@�Tq8�9O"-�$��F�/�}�Y��,ϓ���\��~����̷d��coQ�N|;r��&{��b��h����r�1a[��,j����j�����f�+����jxC�!P��M]Њ������>��I��Z�:��k��&	"�]���F��R��3��M�w�M(�u��{ϹB��Ad*�b��Y�w���槜l��@K;r�p+�*>"�o"�k�Hz/P�toryW�d��6�*���p��]�.�l�I��H�	����� ~�ڮ�6����|�(���6n���<f4?"�E��-�������5-؊ମZ�Ya�;8C4X���D�"��ǒ�af�t	���+��8�w;m�f�sf*�@����U:�ʛ�L]ӯ��p�hOu�E �?���2ז�mY*1c�.�5�!�/�@�ph�B_�=���g�u��!��ʈ��$�c���3RI����KU�hmI^-�Q8V����|���0k����n�;�7�2��FpJ���Μ23����"X��m;;g��4�$S�r��nkY�f����k���`oj��_��0�>�J� ��h'�(lW��3�o|f�"��` �
[E�I5U��{S����&f����Ņׁ��z(�$�3�e�\�t�'w{��}8r<�h�ʾv��z��$�;(�(����;��.�r���F4�GzȝY���k툉S>��q�c˜;g$��Z��(<Jq����Jf,J(�Q�%|�ͨ/��%�	��c�gFm��VWY����KUW逡���&�R��s��<ʓSq��9��V�I��A����߷z|�ڰI�|�)k/XxJ]�R�͖���T�I��	.�;�U�q	���W�,���QK�RE2�_��>�Yu���m���?@Uh��Q�T�jŕ;�p���<.��jo���q!^0�@P��LZ���95N!��hV�P��f���e�+�1[��w��c�����~�F����-��9���2���q���<�(.��M(��By�[�J:/iJ���� ��FI��������%h�N��$:��[&����ع%� �i!`��m|� ��.Utµ@%�O�ѽK ����L+}�# �0S��Jx���*u#��������}yIU�-kẐ��Q��A�����BƠJ|��D�|�;�60~F:��g�,_)�^l{݉�*z��(L)��@�&��?zjb�b�s�V�+���Ř�HY�z,>6�R�B�C�Ff�˜�g�ӸʭA���AY��,�w�o���}����I^�a
,��W���x]��#䥠U���x���t�|.Z���q!I��
�b^����-:8��I�(G�"X������#� �;S%��ʝ*)+����g���;���gͽe�I���f�d��*4����Z��h�N���?���$?�yq�5>�b ���5H��b 1� /�c��gģ(O��9�p�.��B�%�E�p�/t@z�&��CѲ,2������M9��!]� �3?=?d�{8Kc8�ʕÙ��X�ZF��(��52�MF���b�܉��Fh?P�rzǦ��"$��!�n��0U��t���܇��&�N�A+�^o|��m�RR�|�\Q	�j��ᩌ��@���P؋S�m}���b���k4�����fl�hg�Q-x>-bg"�{1�e�[�����i�b�B�'��^�W�M��I��8͹e�����q��Œ#��[!��95gf>�A�MJ)�Ʌ�� �ӧ�Z&�<�G0����by9	���co����oi��f�hɉ��}�Q��#�`�KRqƶC�z�� +�MG�"�t�0�ݥ�O��h��[��"C-4h# Ao8�JPS�E�`�PD��LxP9ڬ~ 6��Tu�����df���۬G��d��;������ [!p ��2��[GOz����l4/p!DP�2�}AB8�FFkp�u`Z��j��m��$�`�#3��O���l:�9�e�-� kP8-� QJ��߉�zێ�X�FQ���%�"�qW�RMr� ����*�̢���i������	���}�@JK.�[�~�:W._���t�?SGp�t�L3஍�` ��	��s[ޔ�Uh�<���@�8���!}l.ɜ�W^�J�H���9�)�0!�j����b�xS�CC�<π&p�o�,����r��OBX��e;��a'/�^%%n���#:�{�VG?VI�o�xkN�Zb�ra�R}E:�\���9��4L��^c,�����f��<��[5
m�Im����.�����K�x��K�5hq7�>�ɨt��w�C����{��;�p���N�ཅSVī�d����>�_y08y_g��`�bh��|J�r8��Un��Ko�)vJ	u����5/�m�����B��.!�r�}D?%w�ؓ�Zxa���|���I��)��?���@LL��=��ֿ�q�̸AE����K�p�b�$�ڔ��,�a��>�"��,c[��yfz��ߧ(�I���/�%a��G2���x�T@,��;���pwՅ	#E���cN`����\��?S1D��a���=cW�LR�.����ա��p+�[0��s�I�Ȗe*�VU�r{w���W��D��ɚ�d)i����LK8�/!�3ⵤl�֧�.�"T�o'���A���̬^ɛ��|Ǯ/(�J�-��K��z]�z�q�IG��\g�٩���.�������nq<�����k�"I��=�'��Y��Ȁ:�:����<v�[�ւ�4�9 ��� g��� =��"a�M�����o}"������Jۇ���w���3}oB`�C�g+��UÁ��<�T�c�9��;��9r�úU�5�f�j�d1��@b�i�_�u3�F�� C��85��D�"�l\ s$m/�[	E�*\ZI?E�ˍ����k����ZY�nȆ�/�&����ӈ��z�,Ѻ	�I���F*��<�&�~��K�ÝbC��0�m���0��)�ٞ�PR�SGZ3���)����?.V�������q�J?�0"�rVCx�b0V�V�!�Z��cɯ�`�굀��GG�x�D^���� �P�H����9����VS-5�p��s$mw��S���G��v��<���'UR̷����s�$�C�i�kÚe�a��:FF�O�\!������jC�rg��`�&5B�&,�|������H�ړ���a8�V5:8��]�.�B�plve���-Sqa(5:��-5d�T�e[���SAy��<�~۱�P�R퍅c�3�v*)W�Y``d�N�v�C�]��w��$r#�s��t/��+� �u(��R��:�^l̨�~T�%iR|�"�<�%�%ץ��KFjM]Tn���L%���I��^�P8f	E���9"r�������ۣ�p�1_0��7AoڵYv�	
�!��G���#�C��3�"@�+�m�lV� )n�X��Jn>3�A�r����q�&�׺ˎ����ȅ�;�`k��S��x�:	J�Icz�p�y�Q��IdLeb�j��2ZB'5�~�,�omX*D1Sא��c5�t�����_9
�Gؘ(���G{'q��@��X�A�H�b�D��;�����&��5"{��70z��I�G|ȯy�5����p�P���w�U5�|n�%�O
�cY����l
�	ءX!�ၕy����]��!��V��F��L7u���x7���=�������=���SjbB�FԞN�q�.��[��ܭ�בg�����R��*��h_�i0G��lA]��-���0�>k��(�����PN<����P��!ȾS�=�qt��EV� ù��m����^��o[~��a�mY���g�E2�����B���a9sdG��eza�C�doE���]�:���e�J�w��>n<p�-,>*��S/�����'VnpNf�����qܻ<��gW��CҠOF7���T����N&?(�@0X�1�Xp�}(�U�[>�Hh[ �A���K $�E�@JM�T��1<��=7�#:d�������+�t���ؽ��� ��D���a��k�*#]Dbkq�?w�Y�w8 �o����m�>y0�L
���{y��Uޭo�gD�鿺��W+N�#%w��Z�6:�!��� ������	(>׆jz�gdpn�;+1SA!]Y�	̈́wp�TT��C>�<�U�s ��g����h-0v���^25єOJ9�C%b�0݊� �=�2_����v_�Gy���(y��X��B�YPa����hZD1	��v�K�s$���\�	߲J���d[�# �G�gEكr�Bғ�a��@�	G$��͓�ϼ�)`�7vV,S� �b	�����ێ���)��lAP ��>�;���������[g��y�,�$��kMe<�(6C��	�j�WHfؐ�ܺ����X�|��n݃uC�e�v��&�h+̘���K�����3*�_Og��j�9�;x��c�"�QYk|��hx�-|�����o.�`Y��_����Z�L�A;
Y�*����q���W��cL�:u��=��P K�	�<�uM�a8���ײ�]+�i�B�2�0�Dq���X`=&?"n?-5� �2�J-����s����[`�~XB��W/]���{>Ƅ���'}1���?򣏱S�7C��J{��k��2��k/��W ��z���pR�t�)뿽�<�������R?�g?iU�T������s%��w0���7�*�,�&2�!��=+��T/)mԄ]n�6�`��aw��>���[v%A6d�)0,�V"6I�U��v�j�XBU��y��F+����?�YA� ~�I�>�ܝ7���5����zj���ha�Y��*���q���N�2(�9�Rx�
n~s�S�z�W�(��k��'˕K�����|p�NAD�����'��G�Fc_K�ӱ|�LmX� �M��yz(RX@�5����/�bp��!ߣ���a���JM>h�E:���>��F�buS���E��h֜�I�Zwj׮uV�c��T�M�v�M�w��*[�T�l8��,������Mٞ�Se��feOlr�[��φ�߽�N��ʠ�t"?�xRF�G�U�=�l(J�:�����z��wt���TFm��F�9�,k���E��e���W����"A�T(���DXio�y_���+�F��b�yB,C�j� q�a$����/�-,|�U��-�J����|���yҐ�u ]�O�Z��Ű4K�{9K��RW�.�_���Սb�0�)�ڌ�t���.$5	u7wv_�F�䐵<��`&
�b#�*-��7wM��n��u)�b��#�6"R�<�8��ٟi�8دm>CO<����_�X9-M��_���V��m%Dw�&���&km��Y����V6��Ih�*�+G zM2՜�������Y\`�������9����uS�0�L������n��JlyW=�ώ��kZ2=��0=�A}�)ᜎ�u{���|'b��+��a�?e�̈́W��
\���l±�hq�vi�����L{��J�E!_�e���:��A��DI����d�U���W�E$)^�3�$;e���X:ZNi�H þ���rq�+!�IR�� �Ǒ �ÓW�[�(���] �>��E�.��<�]K�bb���gr:����=��eF��m��o�����nw�Պb�	�(F�^��$��ҾP�������ÂB�
��]�sf��G�g;)�*s�.&P�';V�|������ �s�V���[*�Kmʻ
o�bq-=��� �f|�Wq�;��"���3��4;���t.�?m!y��M�*7����P��~��.B��-�L��s��M�3��8��ʗ9QzՄф�j� �bF���u������OU�"yȎ=�v��%/�=�t�Hu�.���C���,��(�(u!�բQeJݟ�Wn�.�4J����-�ϽhS���IC��o�gxӔ2@ ��ɳ��P�s����� ���i�"�v׾~�Bx؃$����!�s/���	���ׯ\s����K���x;1���֣�h�|��eŖ�(t$cW���ڟ&��>,`�h�7�9���v�~!���t ��(LJ��@�&�*���#t��N��F���R�w��~8#Kcܭ9Z'�o.~����E*�m|["�7��+,��(QDcD��1�M� ��W�FQq�����\SM�/l�.	Mxg��?' Xڭثq���B����N�s�÷�'�!;����/�Q5.���� Hp�:]�����t��}�l��*�WM�2)�j�]�zW8(�A��N�?�����d�O��Z�oklcVq��P(�Y�+���U(⦣�Ȥ\-��r}\uYT�9T�y�c'�f���Иa]?�kCNv����-�\���ͩ��c@Ҏn(��Nׁ��&�>^'�H<�n�t���Ug�<��і�����e ���b�+گr�^ ��m�˼Z#.�?^;o���"s�#�����=�rH�P��JT����j�ܠr��ڇ>�4K`v���f��}��5�5��U��bYC��Ю�������Zا�,��?^���F�&�mIQN��WLZS�T�i��~���OK\��*/4GS�V�w�߭Z5����l�򤐋�����<��D�ۅ-lڢo�S�C:#c���	MzR��*�ϭ��_�$D�0��h�:3ym'���	������%ʼJ�R�z�m]����j&�Ժa�;��)?ټ�2�����#8~�נ�)�kX@�@��=0�(�z���gN�^�j�V,|��;&�xU�,�<w�;�A�׏T ���k�A5�il�p���%_�b}�K��䜻�����W,��N`��\,Z�ʛt�HL� �I�B�̥�"�e�N)� ��@��+$g+�S�y�u�]��HJi�!��693��.�bNG��3�Y�۬�����/���&�bx�ۼ%|����\�ZN�*�<���2�d�0>d�I���$��S�Q� ��)Q�J)w�S�
�-��?��{'D���Ħ�� ��vr<_�Ġҭo���?�����v��j<�{��م����k��uɎ���N�j�+�v'��d��)����<�ߗ:��ȿ�Ê!u�_nǒn�q.��� e��Qt�fZ�~ayַ���NF�aBV+�2���OQU<��JgkN�6���B�'�d�K ��'Bi0��%(�x����t�|Q��h�_����1B��ЍD��gP@�Z������i���U٘���^���"�ųӚ����d�H3�����1G�T ��H��7!�/����W!?OEsXG�Y}�@{z�����]����y�	��9ꕖQ.���|�4O��5Wb��/�����BS/SA�H�+d��p�3�8O��ey٭�fo���4�$�-����ݜ�⬔�s��Q3�M��f�)-���~[��G���»a�d�4��ǴN�C�v�(�k]���&|��yr )���ϵ$ʖ�&��Մӎ�hC��jk6��E��}��0�GC0LR�H��r�!ө謦q^��
���D�����\����_W�єh]i��h�^�6����X{��?(M[��`�(*��,�@�ۆ�������2��[)9,�:J�W����Z[S��E��ܗi���x��V&����IAhT�1G5�:~���
C/�i�,7-�Z;׌��H�x��?�Z=�o�|�������?�R�~p1������8�7N��N��m�U߯�|t>�0�<VZ:�����C=����2˰,��a� �h��K���@`.1͗�jS�DU%Z(پ�P���T�*^3}a+lWq���<��V�pFL��IX���Tu����p�s~>i��	_��4��-zjH�ǸKCL�_y�R3�#�c[`r��6�%���QU(3��@��G��N����(���CT� O���+��k�"�3�� �x]�I�*���LݒK�~Wx9�c{%ȸ����Okc׼\z���ce�2R�ɻT��~5���^�*�wU����K����T�>|��>�h H��A�K#R�v�1o�S0]���1�Z�O�	F��(���A����uZ��u�4\���Sbר�7���x���M��,U3�X/�|��܍l�5{B#���X���0�y@O� [TJ�V���>�J�c%�^����gw��`kR˘MC5�����O�H_��f3H������QIܟ���H�7��[�%äȿ������5�r�Ē�}:��)bG ��0�i���o���;Xs���[����顝��i�<��<�jk���n�L�(�Y_A�&&4C�[)��6��΢bo��4	�w�
��o�5w!��xc*��ɲ/ �o`�;I�#�.�`Tc��� �N62���S8e�@B(~��e��m�~�.��-�F��oF������b&>��UM}*y=���I�޵�M�28S�E�S͖� ��(�y"�&�TX3��A{f�iݸVi\!�=A��$PGxS���2�iGC���7�ϵ[TmĆtz|���{�?GN�s�J~��^��� 	�O�aT�Z�@o��Ônc���L�K0J�-���T��>��2	>�]�[�)p���n\_7���GC�8:�Ͻ�p�u�3�z���`�S��y,9K�y�A��I�:n�Y����
׷�IE�/,� Lf���+d�So/P2�s)B	�aItͅ�Q�)��^��sb녆�?��#�!�g���=0\cb��#UTEßS�tsx�T��t�R��9��~�qe�'�}ɋ��T�Ȭ�&��Co�9�~�Aш�8YS�/�ވS�kИ&��_��&�Au9�Ţ���On|�^c�!�a͢��#}XH�T�wˠ��o\���uA7�@��y�ZSb��E�k�$��u�lg��2�&\�\�����[�/ ��[ep7�t{V^ڈ�*}P-���2�b�<R�Coxt����L� K�eѮ���U�7���8&h�^�D��	���:�߬�������)95���Ȍ���!kxV�1p/�x$����7\�@����
;U{�1��e���c2]Y7�t��qf���w=P��:����,��s�Q=T��Я4$#��(mP�O�k��a�C�۸�~-�=O��ne1� P���K��,�o���C������zL؂[e=���2��sp'@ڝ��^D���`q�t�2�_��>zP�t#7�%9����W+0_�	L�gv	���8 ��Z��#��Q�W����1����s�8gb����`�'ԷZؤ�A�n�`e�)��~�o�|-gG�C�ɋ�uf+B�]~�:bIc D�rWةFߗ]�G��z�^t5�v�Ua��ڙF��Hؒ|#�핚C1k!���+f�"���-z��.��Bzh��2�l�=�,̽���Cի��fZH@�V)���;�r2oT�hV��_d9Hz����� ���r�@[���Z��-�����)w�u��ns�����3����|�c��T�0�H� =�M���\+�<�`������{Ot{�ju�e�|4g9���Z1(�����%D$��b����
��l��#K�jq�}�g�xj�Q!�<$���]"�1��3(�Ǎ���W�V�rn�F����E���ېZ�	2 �Q�Ψ���V�C˳	)��F=��������4UUn��G�K�s�_�V�'�>
���j~�F]��mO�[:�E���������	2��WkV�Tb.m��Y�Q�d�K�n��4mi�[�_Bi�Në`�#T��6���� 2�L	�Ęg��_h4�=p��_-�����o�ݦ�d�;[uKԏ2�>�o	�W4^�\�����Z�a*7<��L6*�H�EKB�?XJ��� ���a���ϐ�^�|�U�B��1������6	�L�6�������j
{E�e����7�w�����d����<������)��o�Q��I������8��_� ��<@�47�<vu�ꓴ�B�Zdn�w�#ײ�������ۑ$�>N�G���V�m��<�����W�̀�<�즁���rtU 1m�a�8���E��b��r@"�Nf�w�F�A�	`�CʘT��u`׊���'�4�^�2ӜT/m�ۙj=@�R ,��(.b�z(,��ǝ�a�_M_�����D
ٟa!��<#}�@	�6�ߤ�2�N�����j��ft�@�+�b��L��hr��T�O���R� NV]4���A ̹;�ȋ2p�oÑ�JYx����Dp~ ��0�
��9hC��T-���݉k��1�ժo���*s�B�R��-��F�vNc�)���?�˳�}�|��)_{ؿ8�� ����zzBL����F��.��?-)�=�-C�<��ր�U������HH��W�O;I~�d�ӷ*Fl���(}_�ё.ӤI@7���:q��I��Q^A��^���܄�Y��,:��c�����~����f{a����(�QNE�#�(9jC��ٛ�Db�������a�S���iBdЁ���-�5�Df$� �� M֔;S�� #�z��;�)L���/?<Ld�q��UO���ڽ-��XID�� �o�a�;P��� I$5�䫈�Է�V.����@I&��e}���s��Cn�)��Z̖	��B��R�Ő�&5�)��T�`v�;�J,����4	ֻqU����g}��54���UN�H��Hrw�h��eD#pn!yT�{lM�?� |O�[$�fO����
�,�R��T��hg��&���?�4XI�vSѱ��ʈ4$V�����H��_~s�x�t�`݄Z~ǢS����U��Q*'̣HA����s�f_�!���7빚+�
��i�2i(�hg3.�I�	2{R��[r���tL�#%v�r�?�]%�ö�3�OauL�se�jЖ<���~����p��OARp��v�m�g�'�*�5K��.}z�"��_mF�%�B��܆����(ʱ����`�>�z�co_Vq[br�]�A͇s�ƕ~1ׁ&��d�5�,q���R�z��4�-Џǂ�C��_�7��Sϸ�[�ա���1N�h�E��Bz��5�U�|�dk~���V?��go���*q�o�'��#���D
��M�!���*d���I���F�E7���C$��t��$���1��I;�>Ƌ�'����u,��]g�^�_�%�XCv�����4C�W�����ʊ _"�h����sN�=b���ٲ�NS�~��>�'*�C��v�cV�eG;zo��o?k���KH1�`�����T&_��9�m��t���-6� �}�,-��ɥ��}ˏ�ft�ՐD�`(�����Zt썝� ��ѪM o�^���CG�e?��3q�^x��a�����򀏚,t�n�u�_}*靂«�B�{�'��"ڟ�_| 3��a�I�~�n�ϙ�&k�Xڥ�{.
yg@��F�SPE2���Y��`�0=�Q����K�i�g���L��#��F�ML|A?;��rW�
�,��2k��"��]��I�O��r�I����O@2�^�.���Ww71��hߎD�ɷn�mX�m/d�y�L\vﱸ\�m�;���2��b�+�2�DI�N��,z���8�f�wA_6��t>D��V�s�U*�Y �B��ߵ��#ʲ���٣.�M�\�z\X�+��{�O|r�Z'.ޗ8`p�R��W��h����fu��'�e+8���v�d	�A�
=�v�2��0]��Z{1"N�gB�
n����� Oa?������\����i��u�CL`�q�}f<�}[҅�SyB��0�W�b�_�s{2�uA��Һ2�|o�T.2(���[��<���݊�� �O1� |x,P�c��� :?�s_䛆��Z�d�]��7���__�vj�� 9��J1������5�y�x��)�TJ~&5_�q�~}	^��_�ː�X�e-�	;UbeY��ѥ�bM�j�Sv�D�L�K�y�s��4��_�����u�#�ҕ�M����r�
��kK�~ͪD~�C���8k�+'2,Eu9B��C�4��7�a�o(�:�̠Ou��֦B�*�5J����R&t4Ho�̄��@W!�}3�9~���	fD�*�:qG'�l���z� �'yT����eů�r�� М�ѱ�w-N&��������ۖK{�r�l�"�٨�=@��#����lGp�����QI]�V?��gc=��Z2.34Uf&��ŗy�
�N�9��~+�H�ȓk�U�r�0�h#aSb"8���m����v��t�^�y�=��7��_��z)��"�S^�~4��f�	u��^m�3N�]���y�<ЎL{�j�E<��;�Aҳ��������n���f?�j��RU(V�䏭mC��ScҝV!$Da�j" �-u Ʃ�O�,�w�hL�ڸ�Or5Y�HS(��	#��{ Z�DD%��Ҫқ����5AҺ6E"�:r�M'� p~κ7�"�AYE���in�9=�d���a`]pa<�}^"��a:ܖZ�#���tY3�`aҶ<~��M�3��nl�G)|)?-�yN=��
�L�G�"�{��8D'q03���LP��%_���.��ia�P�.�w�b��S��j�M�;��q(������/2��^�vΐ*�h�xSJ�q�<������U$B�Gj��;s���8K=&����m@���L�z���{�a�9z� cJ���T3�/���V��a3w%i���yH�-��>��!�Y{:&���Q�Z��f�&�%ѝ�)�\A�����`^��\�T�%��!U"iP�����^�>��M��m�2/�i���9�=Ɠ������"}�T�@�ؘ�9f\�����W�zh1*�Y	?�!�c�<pA]���KPh�Ԁ�%���1��<��OΦ��w^���NF�L7���n$�
	�c �0��w9�����}��@�=�x��~����1:�~�s﹁j𽒨�����YK��/��_jΞ�ca��ŨH�­GY����? �[��	fiz,�C 8�T1D�^/&�'����VTLT����e
�5a♆�������(x~C��rP���_��d %���&���,^d�>k�E������˟{z{�:����Ws���f�#Մ���ccL	>�� ��'|�q�i�=�B�5jp���?,Դ�x$��Yx�1��;�8��Ic�y�-����d�N�U3�Y����+`I�\���_�7r'*�>�Mr��X���U�#���V�T�/�l������P��Նf��H�}��6~y���X�TX&�zp�	��T'��u�ߌs}ʔ`���ߒ��	���eyp���&���9-�h��j-��S+�c&{��d��At[���4T�I���7&~�}��i�a���W��r�5> �LO�K���´KM̻qQ*{���LS�<%s>������:�M��$��0�\���c<���nD�
�i2����?Wp��QQǺ�}\k�/�E�"_�k�� ��������"R�)$M6:��QJ5%@�V�75�L�f�i�^���9���Z\��EO`g��	c�p
�"i��}I���^�9_�񢞗�|���Z4S����	^�8�(]g��E�J��$n��{�	�Ao�vp6�KW�Tw���f+�G���
�^��	�(l5�0H�E�KC����;� �{��3\�H*�ga�>�J�e\-RGP�˩;^p�kٷ��`��Q���h%�w>6(�L�ݗSt����9��XR
KA�y�����=�� ��;�h�a��n�fju�
Ew��J��C�`���5������.?�YotYޖ\���!'6��4�j�V9��"��%k��R��Z9�uҮ��!�
��v3s@o��s ��:}[ü6G�TT�d��5�@1{�ш���f�R���~��c|��|�i;#*"���1�3�ub����$K��e�z���b�} �-B�i���Z�%1����y���d/m����{��$�R�A5%�m�	 �V0�ȳcXB�RH�:��/�*�i�B��L�L1��⾈}�x��v�RO�@Y&���e��0��L8
']A=5ӵ���/�t ��~`��H>$dz�y�q�/g9� �H�'���L��Z��`���	���?�<*���sS����j?"x1���y�<`8���"��ʭZ�E����b�m<���; rv4	i���鵏���ȊT�WQ?W�s��WSĪ��r"��(m�Ժ�W�����'�kS����w!�Yp
�d�:ǂC�E��~2��OB.���|�t�A38��M��?�N�U�?�!Ca�ગ�2��(�X@���v�g�3SM���C_��Ȁ�y7��.I%������K��_�>��g���K��"����k Q:�8^ʂ�z�� �-��tzk�m���<Z�lLW�}�����f�ػ�dͥ�m�)��0s�媇_��Vnj�ͭO-�_��0�q6�۲x�M;5�eT��;˩�����C�$T�C�9�b�6�+d��` ��;���Rʞ�ۣF�eT�pH�#��|QP��4EJ�z;���UB��Y����f�B��J�fC��,�q%|O��`YAA�s]%�*�q��v��H��ZC`�O���(��͖�|�&j�q���j���J-1Tl������8p�����K��h
�m���Gk���̷�w����:�A��� ~�Q���S2x.��1|4YQ�T�f$�.�&�ĸy�oy��,|d�-`޲h��B����b|����4�Pw0��i�w�Ik�#���c��$N�2�텶(���хS��I��F7f�OUW&T&��׷���k%3��K�R#ile��P�{�^fx�n�l����ٔ�V;���O�2��a^�J��.3�*��y��ð��Gy';T�b��@#'���_�0�)w�<�۸-��Jߧ\���4o�*��!�Vk����R1�<�I�z�V�)��P���r�����_���m,p�5��۫.�	J��خ��2EGV"r��M�X��8�O�xU��<��,v��a*�5�E��xj���ԏ�𩱖~.d�����zZO��kW�!�_�ͬ��/�P��屩Ú�/z5��O�}�������ȩI�	?��@���B
���S�������>%MHJ�%*�7r3��=;��s�BT�U�a[��<����O�j�N9ԳOxOڮ����b5�=�%�xɶ��tj4�`�ˀ��$���Pi;M˃I��	_,/<"޲�q�� Kb=:Ҫ�����;p Tw ��s�^,��3�-j'�Xq��D��S��n�o��˜�(��Y��c�Ϳ�vJ�]N �0��Id���IQ�E��N �^=/��?R�}��M�}�V�uPͳ1!|��YD�_ 2�E��"��\��������ئHtYF�����s�%���ip�v�ߟ�ewVqq
��29.0��
̒a���>Sx�5���K�Gi,TW��SMZ{N^�5<n��`j�[�1�3O��0�9�i<����7�y�k��IuR����@rj�a�5�I���l�h��s��/��;Rm���'Q����P�\h�ĥ��}!v���Y�-���Vȩq����=��&L���o�H�ˍE�j	ԂI8V;��}�Ş��j4���G�*�P}��lW�n��
n'B�v�/��nq�A	宸��(г\~O�@F�k9�LoZuvN��@eG�sH�>(���_��bE�X6&�k�aƞ�w兪�蟏�غ�[$%Ռ�֢�>�������O��ނ�S�E������۾�'�A�o�
q��ͦ�0�hש�H����@��B}�r���$�\!���@f��wc`�mY��)��d|��1�ϭ�F�f|�eo��W��*� {�z�B�hd��l�,�'~��2U���w�jr���q&�#ђ)��褳�YCz��1��p�7O�{%��&NV,��בt]"1�r��*F��V��ri�t�D���Y��}���޵BR���)�����:߲8?�ߨC�1�Ǌ8v�߼�8����G�H�'�­)ɽ�;���L��I�E�w-�"�}��U@h6�p!�_�?TJ/Dƚ����syf��A�~Ԁd��U��5��&h��:����ц�?d&�E��*�I���3�nr�1$t�GSx��D�/M�^Ou'�X��~�� �}I\�~NhP�Y䛁;i6̂��{!;��20�xU5���^h\�0���?ȬƁɩ�C�<|�e(o�: �>}�:��Cs�7�`�S�ůw��D�8�Qu��5I���.F�c�D��S���+te�d��Z��3x��=����ٟ]u�og�Z+b�6��1=u��C� ��j3ʵF�V��x��0�3n�:Ii��qg$�$��E���O�Z�0�u�`X/�"��4��fw~��^V���������[T��NNw�@�0ͮ0��e/�.n�$nfi'�LXf�8�*����8�X8s�"��Bʎ�ј�OcjY?N������#$Eb�b�#���fjƌ�V܉>q����
�n]4�?`m;Bd�t�!Hk�_
w�Dl2J�\#�y�=�*�idm�Q��vu���ʃ#MO��>յ�^�ʂu���\ڏ,Cr� ��[��w�U ��]N�Q�OB�VZzl=�!�B�x�Y��n�W>!�_�wJ"�9���N�?�����|��+K���/�ژ	��D[�b�$��~�Q��}��K�� �Q��#W���`�+},w�NQ��沒E}���c�D'�V�x���hay�?R�6���P�KX��8YDA��J��ylo|3xJ�朢<��	fŸ����
Os�3��N��R�	ަ��Y{�3��!֪$2 ^�ڥK+�پ e��w�x�eL���RH�8���-$�3߉�4�`i5�C���1�_���!�dg�w����D�	Ia!��aC�ЎG��e�~ӵH�j����h����Ův���8�e��a�RҘ/��J��6}�<�c&}��ug�T�k�?�Q��Gv����K��x��"(t|���8A�+���7+�s�&���}:�1�N�t�����m��矗����#B��L�i���uB���d��\:�M�Y|����k�ڼS&�����P���g�+}`_3��M[]w�n�|�+6�f�#���Z�:��ь0~?J�d��Zk�R`3rk�V�h�����Yǿ���{˘�����K�G9��2uG�ſڢ�U���@aZ�Q^zv��u����о�_�^�]�oќ<y��X��W���x����Q��F ��g��5Jm�q�.O0/��X���J����ex��u�i3(�>��U�c�ZM%�{��1�a m� ^���h$^�ߞ���ep��]��F��<�͊�O�*��&��ב�����shNHj!�Ԝi��6<�J��d�)�tqT�&H$I���
3�5�Z�٭Yr�fϏ�;3�S����c�� l���K�C�L�T�tx����Hv��]��^w�u5H����:�&:i99�dL�s��5��Z��j�+~&d��f��<N�K=�Li�Ɖ0Bc�X�Q�i! ��T$y<���8�K"�}	=r�z�hB�wd#0����Xd.��8��i�}�1�;gfV���}��d�3Ƚ�o���h�4�W�uE!R�L�K�����퇯���b�0�d�ܝvc�()3���Bҏ��eH����&�o}>Lf��=r�t(K�'W��Nx���R�R6���S����lbl!�,��
��gL|,����\��M�s*uZ�A�Һ⌁4�_��,5m����w��x<����R��=Ρ���	q	����A{���4��k0`:��R��%3;��QX�i��#҄+o%U�~�+�G���V�m�I�O82V�οЭo�2�p*Q�؁��=�^l����zו��>��������@���p�R�Ee��o��U�C��9~�O~t��ݿ\6b�?3 ,k�\5DW]���y2�#ͫ��,K~�v��"NNKdj�֭V�U�D]n������?[BM�RM�(��H��,*&l��S�!]鵘��}2K�yEh�+mW^N����Ek$���	=xt�ت2�pE�IPL���.Q9�V"4Zl ���c��Ԛvm�X²SyT��p���Lļ�st�]���wP�i���v����*�^��N����8Rv�u57h�`�'9�r9�S�Gq��+��e^	���CR���X����6�Gڒ�'�4G��4A�5 4�v(tx�<U<e�"J	�Y�2]4A��_6����'\jɶ>�Sy���� ��'��X�}.m�t���fV+��jm���\����'f/�Ρ�����y\o������Lro�&q����S���X�.d�1�R�o�8��^�Z���7^�u�F6�+�!�st�J#w�&s�����jl�Ä��i[+l�kC:#��G�`B�a�rG��@e���ʮ畠+C����N|�~����F��HA��i���k�5A�=����Ѫ��J6����(�>�؇��Ε������ܝ�w�.�6�W"؇ߛ*�JB"�t�+�>?��~�����݁>#5�=C�U�Cʹ8���:�ւ��lX�@Cxӌk��^n]Ы�%����|~
e#����а,�t~0�'Q2����2'�/e�/��O ���d�X���'ώ��;�Ρ~
���{~��6����a���{M^�[	����3���B��K���^�9F�%�I@v�o�߻%�ε���z��C��~��z�,د�p�Լ�`�g��5̸mt�N�,����'��&�(��&_�j�5#��!a�T~s����8~<�L�y�P�e���1�O>�sj^����Н<�q��M�i>pXy�\}��_��*�j˦ﰸ�]k�z}���G�}kZ8���͙�b�d2��A�h����'���E�;���4iM���*��Tf���:���]oK�o>�}����}���ɟG�Lä�}O@�"�P�5(����U�V֖zOΏ�N�-F\is2]j9�Uz����7r�5�0nK�ri�Z`o�Y� �]�� �zO �����|S��T�Sۇ�H깽v����I嚓.�26&�v��vi��$�B��y�ba����պ��`�:������J0�;^<;2	����#%��(g����
)ȑ��ۣ|��ӎ7�,?y󃽻���*�U�9�ۮ}s�P��H����p����M*�;#�nOY�h+l4?�M<B3*�hSd������y��%��v��ɘ>~��4L <��&�QwX`9ׁ��9��{D�wDAI�x��g�gB)�@./n6vW5�QU��`����}��F�I��Dg���5B*��	��UiQ{%㳑��s/҂�rJ깽����Y����mdkE1�e�ɞ/!0�
J���$m������?f�.NC�:-[��{3UJ����º���i�D�BH�X{
���ת{��'v I+6M��"�,��=#��1Tb� �'�4��n��fz� ��;�	˶��� ��p~�,>9�X�23��E����a�`�)t�['P(�r5�y�#���;E����{�����a��\T��Iۿ(�&"~V
I*�Գ	x�!%UMX��lpf�aķh�7X	dV �	B��,�6�<�ʆ��J�SRzEJ��:z9�o���?��í�2�ە��o۳M�������zg�x�y�J�4�/��ll#?x��پdUyOfXs��c�Ob�yw�3X !��`�?�Fr״0�O%�]��6�a�Tmd�u/F
�g*��#-2���|g�fr��-�V�,����#e�,�@Ns`[+JQ8�H�ɜ���s��)���%�:tMx�������}f8�G��퐆A+??�@{i�_XU`�G�޴49�C*��E�Ha���s!yٳ
��;�O\��(�xti�B���i�/�������c��|�y��[P9����<{W	�\�^4�,���RL+�0�w�/�iQ{T�ˁ����Md 0�jq�h��]>�Ew��#�����!�������S�Ԓlz��e��S�&<8/n�B6���9��j�� ��b����8Ji�j�W��A���=�4��G�|�Z���/k�}�hϬ�"�Gn�[PVu��Dq	-j���1�����62Z�o�%1�𬶈���2�t�
�a����ː1�:zo���ł#���P���=�~."3�u��.��t�W٭�����Y�5�����Q��CsE�,kv�L-�Y�����L� �Ii��Bl�_�U���ďW�����6 GF&v�i;��V�H,�'�ϼfт��^zf�GY���~T�+��(9Z�JDp�s��f;��f48J��ct#̑N���P��R��R�h��2��xOxgf��Y��Q��̿���I�7f�y���b�T����܉�q�D���i��B�O{?��澾�Jl�H�tãe���q�Õ��v��ǈ=ZSr�}��,kU�m)���e��x����O�UV��W�
7=����]
.4�*��}f��z�mm�"��9�'�f�[���!�nT�̂U8ϖ���Y�ȡ-c�9�H!aV�X��/߉o��?p,��n�3������U�@�z��*%�Q4�3>�����	`�.O���a�fa�(j�6�P�ǻ�4�o�m���Q� r�[�+���KoG�!�[Ӯ���2@�H\����C��F���Ƨ�Z�Tv�:��9}��~��g��)Y����d��S��@+{�����^�&�o�Mˊ���A-nnT_\Ɖ*<O��
~�3���}2i���ɝUU*��i=����Z��dIM$\$�1G�-t6і���m7��&z�Hq�v�eG ����O���?�~��l�&�&�8�nW>�c|���vU`���z2��o[�NH�؅SHG�@�<������>+�Lz�Y&P�l�2�#u���7N�nNC<�^� ~�g39@���&^�-_��P	gnv��
����;�7�&�:��*>��U:�m����:��g��i����)xؽ2�{f�'ë�4��Ɋ9� �jN�z��̭<?H-�>着@����OE�Sd�L��_v��r��s&
 �f�����=�p�ƾ��ϕ7	\�n�F?7覰!��W|�,O$��¼���Ǡҿ�P#�,��q���ep��(&F�ى��G�I��g�5����]����m�"�X�|W�G�,��
�t���ժ�a�PU`5�;�Bҙ�C��C8/�'��Su��#��U������B� l�-)����,�*���բ�����Y#n�z8���g?v��˓�`�������o�� ��;Zi��5�n;�x�Sl��-��W_d����В`�P�Y���0�|����.6z룫o5��W��˩ǒ��BM3O��hK4�\���S�	��:���5���B�/ū�Z�X�Q2��4WDQ[@�;A{_�C�L��3��|��ܳ�5�Fkw��8�Xk�����@��-�q�An��MPn�86o����V�-�C�*ze�����Z�z$�@nz�o�A��_�i�g��YQ�/	M��=K<�\�lt �� ��k�]�Gk�v"c*�nQ�[U�JȄ���y6�[���].��6�����3�W��ğ�ܞGaذ��TA��e�w�d����B�d3ۥ���5�Hf@��uժ����hh���x�,�4��'7N�V�R�mZ<Ii
�VIn�N+���'�	���Ss���4u<���Y;��$���DZ��y����	D8�k^ɵ�*�H�	2������y^c�EcP)��H��;YggÑY��|�b���L^j����
?��*c#Dh�R�C���;Q��8�WGk\�ۄm��y�hǫ���R^���{�A���6հ�o	�Ќp��M�Ԅ�k�Z�`�=pT�U_����^�P��Q���Q�p�c{��<z�pL`t1���oDV�u���#p�����K��Q����ҏ=�%yz�H��ϬL�Ì @��ÓEf�,9A�2�?��3(�k����o����7���Y鍣S��<	�q�S���%A���R�x�"7��n=:��Y�%�GX�G����gz��_[�4��i��ś��t��"a79(J�����kٜ�Mm����H%y�i�N�q���H��C�~b R�p����~r�{�N%�������ܢ��˔2t���:��8�����@I,����;�U*�B�h��ː���	~���$wI�ә=H���(e�G��;�ںK�*]s��}��$�8�X`�1�v[�5��t�m���bZ���V���
�[ ��Ǌ1q�U)ܮ��+��wS��.G�Ff%B˘�"��C��&0�� +�U,���qsjz4Tetha�f�������n�{��G0o��5tħr�5nKF�m��Pm�O��]�ؖ)3:kU��ş�~L���nrMru��*���{�������bP�]���I��BSZT���i;P�&Ϧ��\��uB���?���kj6r���{�Z{x�;⴦KͫL�����^0�W^�!|b�2C�{��ۃ�:��K��Xq��m�]X|���e(DM(����}�^���TD��$�%� �?� �������覰�B�n�A�����fDp�I^,�D�d�A�J����_pI�N�Lehpk�S�f��>��])�xl�Ń'V>X)������+�Gmpf��N��t��-���Գ�Gu��c�����c��ݯ�R�q�r���^ք}�,�퐪a~�䑙k�O���%D�_6�l~M��+3|B]rS'1�3�H����y"	�wGP��W������"����0�ԅ�pz�$�dr�٪:��1C����Ґd����Oij�.� =��O��|`@������QjY�Ll�����Ɗ��*����7e����Դ�8j������)e�G�
�v����n�r5��d{�1t����N�n6e���l��LMS^;��e�*5�J.����c���b�m����u8�1�EIG�60���dͧKƫ�Ʉ��,-���K0���;hX�hׁ���\)HJ<@A�\~9����UO�=����u"'����>yr��=AH�R����	�uU^�:wނ���7���������ۺu�i��?�
ϰb����:5W�ȟ3��7<=L��B��n@�U�}��Z��ky��uς��p�A��#�żaD��t֩"�y�6�득�����'$͐a>�`:O����-���<w@k���*-���U�ڏ;\����]6�(�]W��דM_Ks�2׻lG��I¤���R����P�s�Aԯ�;F�V��S����G��_�G ��జ�Mc�ވ�h[�nN���!�A53�(~��ۦM�=��f�㴣�J�9.�>����b7J
���`���S�ߴ�!����>�-�˃dcԓ��!�u
��g��R��J�3'l��-�y\ٳ�!.��zyQE��0��E����zЭ��DB2^��+q)ܩ�iH$Ō@AE���#b�/��u�u�Mr� �uW�&�U�6�(@�A����}�C���F�:�H�) ��^��'���ߥ3�1TE�����-EL�����ժ��oJn��ݐ}[�!�j�sٮ&�ʈX9E͎�IXe�Bެhp��Hf�"!���wP�8iV�HM��շ�n��],��XeXލ���ҕ��t�9Kƕ	��<N��}�(���dL��+'+���X��P?�Y�N�:����k�2��T�X��%p��3���Cg4�Ȕs�w�� |��@L��(�ǂ3~ �,��J�����SO%�wp&������������2x�����W����ׄ��S#�n����N�""�0�����|+i"�9'�_�X��}�b�\A}<k�G�!^� �Me[|Y�]�o�<w0�0�KL���V{i��_U8����"$`a�<��Ǘ�JqQ����Z�d۪��}�e��>�F0+]�F�3�X25��q.c{0&��*���F�1����I]p5�Դ�g$�J�:�N�����+T��a�ֶ�[���*����^���c���9h��sϫ��S�/Sy��$��T8-7����÷���m�xܗy���E�>r����U��r�q�!B�U�&C�X�*s��1�R�Ʀ�0���'�#Xn-��b��}^y��wAfQ:.���&����%BqJK�$>��v0�%2���z@}���U�GK��R==��ٔ޵-��޸lwD����}��ȿ~y�Z�L:/�B#��W�N��**f7&��Oԇ=�aM���@�C����u��:���B��UZ4'�ȹ*?E>u��5���OH��Vu�Ӎ4�Y:��:Yv�o$�݀��X��/t�!��c���^�@W��m8�D͔��꤅rM�����x̆7�P����!lҝnJH/}�#i��a�
ތӖ�=�c��hN�%�Zj"J�Y��ם��S���!['F %����}��pkDcl^���V‥yr`s���2�u��	�O��>�U8鰥�����w���)����ȫ�C���MR�C�^��a� �ԝ�r�+�
�t�t�R&���JWDm�q:o��iw͡RJ�"-B��|��t�� �i$DvX:t��>u0t��;�Jev��	�;@�ޔ�v��S�臆�r�kZ	�]wȆ���o�x�������������J�$<��sk��{��Yx]���{.��F
�\��z?��"��sO'�j?�~�iz}�맥�Fc([�U��mk! ��y}�A�{7"��7�#�$���;	�	u���M.�����:�o[��V2L�>R�&����dY�i�B�u�P�}
K��?0�i��`�i�p�JR�ѧ��$����'�}c܍���������O�!�3����b0����]Ff�`ljʬ;��
X��BG����i�dM�s��A��ds�Y₎X��0a�RGq���|����
ܢ���M��}���q�Gbphlp+T3�=�U�K������͡r,�곋ǯ��\:���!��UHs5��K
X���E�Aғ��Bky)G�Wq��+E�"|T͖W\���u�uЍT��pr�3�o�_1���
ahLy�R5��˺�H��
M�>� %��>��G�'���'���l��!��~Q���C���n�%����H�>�\fs���;Ղui�´��ƞ���E�Ҳ�W��G0)�m��?@lǴܞW�JCX�g�6���x|y����)�-�<�#/5.b�isoS���m�h��/T}� o�*R���I��
����o�������ߐ�v�ిe��VC�(��D�Ĝ���ͦ^�� }z�6�=����S��Fl��FP��z���@���jH�	T!~����ʢ	@$�e�I(ք�삤"��Vؔ�_y�"nU��#�y����xL���դ����j��zb�$��ى��P�����E��B}���NѺ^���!Vx��qf"���٥���'0�$�L�X�a
	aWVL'��S���F�bp^�S���\���2���Ω�Ě��6"�bx>��Rc~���p�U+��s��$Ȅڈ@r��sx�(����'h"lv��'�^E�U�t[�R!�TxG<J]	���[q�|�,�~���A�v;��f��慇���x4K��F�w8y>L�Ta��/��kn��i����Oץ.a� �0�_sN������c��S��nƧ۳U�
8b�0l3` )n�=2D�.]SRI?kB���[�Lw&�򓀧P7�?���î����Sv�)[�G_r(��"��׆����krdTĦ1�E�� �R� ��P����$�=����1�U �Y���+ۂ�`�\It;�+���g�U{��#�c����\C��;��^������ߋ�=J��χЋ]��݊����.���w�(�Q�79�A�?�F�ǱZ}�ǒ�����p�oO3k�v�NH̝����l�B�+�#��u�#�<�4����ȕ�5��Q=�Ca�!J��G���T��RdF�{�6"|�~l�҈�3g]�\����b�RVpQ����b��F��A�&��]q��EF�]��+��^]����3k�l�{��Vr̬�l��p@�	A/\J��~f�R�I�H/���/�c������<� ��ww�3+���n6�5����M8n6�'{,���k�J�s���e�y�����"($to�:�-K1�[z�ˉ��/�r��U�l��v	y�`��}�"���%�9��R�/^p%�G�I�[k�/>gO���l���X�`���(�����V��TG"G��+�I��5���Nhځm��oߏ.�}��p�q����)Q��oɗ5����䲿>ZO�g�~���J�|,�w�������[@�3���F��Bd�A$�6�0G5B����?em�Oo�{�<�G㦇�\S8�b׏6H���r%��E\���=>���v\��B[*��׹�_6�u$$	��LU,m�������z'�B�<,"k.ǆ��#7s���(-��/&N��:�y�z)M���4i*S<�K����~9�n���l���VSQ�Q��W�).5y_l�;=�DXL�z0�����,���Y!B��e49�)�l�!(>�w�"���ب��?߹~��}���3��H@��b���X��Ys�r�~Qpॗ�����޼�Z������m�K��t�u,��D����?������i��&�@��THL�\��6���͌+��WM+�.�nd�t�����k�Y�%O�RITZ{��j&b�e;�������C� ���؎\� ۑ�`fvO��֭�W�#��@�KM�M����;'�Q�?F=��K>�c��oSM%����`�(7[�A��g�ەHq'w�`H^���U����~	����5,�a��O�ޓ�0C�
��W�:Rh�����S�苸
m5�=�ݡ_v/%���蛽�=�t��k�}�$�Ǝ�z�EOi�@��Z�м7�_�Gf�1pf%�(!.Q�z�F2�;�gI�󶫸v-+p�F�t����:�[U}��J��zS�Sp�d�^CLʏ��D����`P��9�\�W�sW�W��l�B`1���h�9LO�z%��`i�&��}�=!}]=��@��o���o��E+����7�\���L�z<����=�ڙ5J�*�.�	��O�љ�!��9��d\��$��	=Jv��!3�!�/x��%f��P���~{�T�N�'f4�;v�=���kv���P�|3y�b2G8.DF�������}v�W	��cm��j`�b�ķ_�U�cxxo��V��mT�O�@Ge������[M(yG��M*
HU��y�_�%��_OV�ďo�բ?r�;�k����4c|��*��=�o�,73��!�Q�kz(:#+P~����DA����(�;���)�W�o���|)�yyص���j�AQ>�lOE��=K�Hχ�y?�wZ����Է�}�)���m0wo*���HPR��ㅛQZM��67r�Vۖu�ɾ�׹�4:�s'Q���AWR�[h���T	I�	�Y����M�fܛ��:�񳠡-�x����[� +�7���ܐ�}���O�N�qS:���騩	��8Z�/t��ECU��@�z4/��-��wo�'{�m��^b�B	�
$1w�Oy>�x�5��jx�re��|<ݐ�)V�ӗ"[���,�^�����Fj��BÅ���Sp��S�O[����v�~d=<�N$�Py���7j�J Y�w=����a/ n��0���Ks;B�NuX�"�Y�z-���Q |�S��H =��r�Zh����؃9��e����1�ۀꤩ�}il?"�_���"܎�w�G/�.���O���HD��z��ˬ��u��G�@p�s!�ȼ��h�W�`(�Tm���*i��x��n��җ%�e��A�