��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d��p89��N������Dacf�o��!$��Y���*�#�`b�[2������T��Y�c��iN�g`���	��x�-�/x�@�m�Nyxf�G?�a��a�)�*��A@uY9�u��̨�y��@�`|�����ؙ�v�H��*�KAe��D5�Uٹn~q���:�f:b	 ���5��G��r>��T�CFQ7hQ�fr�|��H9^(�K�L��5�_w��O�R���ƃ\)����t~Gf�;�x���<R4�O�槑s8X�z.��DC���o؅�>��,f�n��4����-��#hp�&�1��ES|��<�����U�o���%/P��Oҳ�VzӕrC��p|δ�t�^Ы��X��o~D*5�m/��+W���V	��_���;���������9NX��h4w/2h�c�4��>�Z�0u�I����c"�B�:Y��.�Z�Y9��w;�	���X��IU+�V�Կ�}pP�;t�X�])�rPE?1�??��L	U&�~�H��_֒�#v�j��Ls��B���d���h��!͆�휸��GЇ6���qŚ�dY՝�?�ϰi^n�=�$�t
��p�hc}��8w� |�����m���:��\���{	��Xl��&���T��Nh��M?
�F�&lh����y�$T���Sh#_�$f��t�b)e�4����s�����h����ߌ]���.;N'�Gޚ�Q�k�������'�'�r�c;�N&D��P����q8��5�G��`K�!�p��AA���H��|��}�}Y{��c�x\ ОU6Ж���1[����P��TF��D�ҊNv:����I;-��I(��S�Q5g� ���W;F��:)��nJ�C4���P����[��"�	�.����Bc�q�V/O�ui�Xxߓ�Yz��m����ѩ��@���O�:T�2ersS�$d�ut�V(�Lȏ����u�bdӉPu8�@��wlK���$"� @���$m*n���t��w������óЧ3��|��g1w�҈��r�l�� �Yk\yn$��{m�����m�n����:��XOC/�g(w_l������r�;�~C��W}7�4��o�x�-������@WG����6Ә4&�m+:�
:�Hx���Ya���0�4�(QO�.���D�$��%&��!Cî*
�����G]��/�d�7ov<���-����#n�'٥�/J��(�{G(	��f]U�K�8����@�FX8gSfO���a�(A��TU�K�58��Fd|�)ff5��<.37�ԢzY�5��fc�Im��sF1��H����&=�hN��~�)^Ep����te�U`Q���O�7��J�T�_��#l�S.^p4�Ϡ�m!~��F����iӃ�?'T� O�"#����jۅCΎ:�?b�r���~�^�����P��9�<f�c,�(�M�Fï��\��R�������'�q�(j��O�j�nW�\C7���K���K\�K^�W]e=���<ΆF��� �*����k�[����p/�efa�"���v����z�}ʕ����n$�!��G�o��~�!��N՘�	t��V��B0�=�d8Nf�5i��_u��x�SӐz�R�:7������Ǳ�����h���I��jM_{�S�pl/��b+��E� ���忌RY#﹃�����5�*�'R�c͏����՞�X{[��˪ꆭ~�5,yOF��L
ϐb��6Be�V�����H''=Ԉ\~�tԥ����g�L��w���ʞ���5={Va�¡T�0X�Y�;����q�ȹV��������|���V�fRc�J�9A�@ZzD~�t���І�:PX�������꤭ J��[L��u��ŊA��@�:#�bB�����S��H��2y
��4��k��͌'�ڱP�"�1��8ܮ�c�@�sQ���c����ކg���y��9�$�B�B��۵���9$��t�)��J/eu�
pn��ɍ�	�%��Q��׀���f�8{_ڝ:Ѣ\蠍�G!p�0�;�]d����:Vy4R\���]q��o��S��p�M��$������!)��旧�H�Uk���E1�Bl�l�?��L� �0�e�lJSێ�H�x?.�rԉ�.M1�C�ܛ��5����9Wd�?i��h�j����b������6�VG�<�`d�wɜ�yn�^�����[�	�zV��K�I��O'����ͱz�����P���P�_w��@cjd|����<�,\��m�5�;!U�k�.I��w+�����������{<y�|W,��1L��߲P'�����Y7E��^h�k�2.@��YP�]Tp��*Z^���6.����F��߭� ��t��h�W�����=(�X����!�]Ʋ��$8����i�Z<(���s�\�=��8���`��\�UD$5��C�W�x��|I������K�A��ޏ8~��=�y��HJ��uc!�qF��m�g�$�!�cOx� �=I�C���p4
n-�^��`�!=���[�*I�A��;'��/�S� |��j���&~�
Y}�jW�`4 ��CaA"*VkPu�<��O�Л����r�]�ۈ�垂���=^����#��q~U��H�YS�}��r)���Eφ�5�ԫ�?���):l���刕�Q5L �� u�Y1Z��@Hū��-�4=i_CE�?d�]�[�����p�2;��Y��n��>ƨ�?<�E�nJ����m�鏭��R��1B?��v��B�������%��>عb+.5@.��l��jGف"�:`�M�n{��՞��}Á�����挄y^[�+�IRz�m"J����=�ѕgM7��~�_++�L0�ų�������S8Y�l�A�̸�\�����O��rm��1}���m�]��p�=�O�m���{������p݆7�kq�Z�/��_�=�n��\;^y���|>d�"��w�\�w���2���C�}�c%��'<w��HF��F%�%"
o�v�����b���=$h&<��#w���Ӆ�Z 5��$ڜ�7WL�ϛ:�Ro�Sx���K伂�	,����C'���s�c�y��d5�_��?���`�=h�XƖ	�.��R�#��	�3�7פ���Y)A�C�����:1V���? ��O��J�-����<��F�!�m�vP��h^�,���Ǟ� ��AWG����(��Q���]^0������Vt�}���]�(�%%1���SȲە�y�:b�R�"P'���,���U���Ps>��~������VU�]�WX�=^P'����s-���d0�t�Hh�5��4�>?b��u�Nۂ��~D0	|]�������P�膀a1Ĝ�7W�3O�2�p�aU��s�~`�K�+,(S����id�x�x��|3cȫ�n���ȺO�.<�����Q��dGx���]yc7�����������!*�:���e̝�(̾��U5;���X�l�!���&1t��O��n�rs�y�7�)��������<)M?�L^�Sx))(���K��[y'y��]��"���d:?���fD�!X�{����s&T����3 ��l򽡢j���i�B�S�p�o8���-�� ��md%���;	��Ar���e�J��|4��`��ⱔ�$�43� �9���u,�уiQ��Ȭ�#.>��Xu�E�5���4 �Eϧׂ�Q���]�m����%K�-������K�5�Ϻ?�CT�-@܇��5;Uö$( �����b�Ѝ�<��>�e'�$�Q�����3��n������4�k윎�O8,Y�:$/��DYd�^��.E	sp>V��N��ꈽ�ٶ�d(���A���Ϲ�"߲��&��2D�s �6</���<_0x�"�_�/e��W*=���n��bz��%]�C�?Ч����"n�G�L`�v��dUr݃e�I;�o��Pi܀��u�T����P��fܮZF��I������w2("�jf���XVe��ݶ���F��,�*���^f���w� ��'��a�{�0.3Z
���1 �;bm};�+���]:IhB��u�В'�w��e7��ɹ���Pyl7�x���D���7�嗟9�N#��	�����V�Rk�%�SGp�sZ��SӮ(3qD�J���y ���D���a��w��S��,�|c(p3����'4�lH�(Q]n��	�Өo���F�bH���`��X!T����Z�$��.�"�C<W��7��9�(�Gŋ2y!{
�7�̃�T��+��"�p���!�R�X[�u�ޢ��f��%h������M�(*ۙ,�ノ6�^��ޑ�܂�FH��B��
��b~���N���|�Z�ǌ=w��N�˻���p��~ ��Y��3��T��F@�|Y^��A���=�-5��M�\M��8�n����g����)��R6�p�TS05�a�բݰt��pM|���� ��ӆ"�����GƝ ����r�hY�f�\ O0���E�=�����r���߿Pyu74�fv�� v�/˨���A'��j�i�n��ǬR�6I�[�+�h4������/N�?"�dQ�-�l�^<r�2f��A0b�9�t���卶Ȗ���>BF��d���H�f i�1�<�4��]���0��&ڗ�S.���bt�:6�%zɮ��|]2~T���;M�x��Yx���&�5�$�0�а��'T��I)EB,�|8�!����׮���+��38@m�WdqC��`67,k۰=��=��>��Ki!��J�U=�~�Ps�9ҕ�
���A[Z�F�� ݓI�<�ZE�
��%�}��,L����*!L��h�]�oA?�t0��U�됓����"B����jؐ����w�#휱⾮�),34��U�� )���p�{��r��;��]U݃-�?ـS��c��*�%�A�%c,쀙T58�t�h�*L�[[.O)��O8��c��\��	�F4�#�>�t{���7�������d��z�B�x-������s�=c�=��y#CR�t�s&1;ۖ�)�Eɣ���. ��g8��Ǌjlh:�G������_|�ŷDB�s��^|ʿj�ʠ��I�M���txw�D�����Ԯ_��e�^(����.��/���/��C�	X�*;�`rB2�$��10+��i0V��"�c�s�D����w���'�»�m�0f��LM��L'�և���U�ȉ��_L�Pf�jk�В�����'�.ն&Zƿ� �ҹ�`�HU�2TP0���K<t 89��p>��������ʋ��˥�������q���r��������{��Q��Y��"��O.��
��tj[c�ݜ�y�DGn�$�}."�2P�����vr]`�4b�U�FJ���t&jA�4��__��S��;���u�4����>��3~�<��-�X� x���U��v���*55� ��8/���?�TH���(๾(B�� E��H6PQ`]�ԕA��}<~�hMHٟ�+����n'F@o��� A�=�2�g8t�E��x�(Z��������N����q���!4���_��T5�������c^T#{��6�w�Qf�,�L]���%p�~��%D�x`B��[o��ӏu(�[���[x?`�,z�U�$Ql�W0MB�*��ӳp��v66��❷��F��C�>�:"�����a�@MD�u���r������6�|wu�s�S�d�
L�U�r�:�N��B�fPCo��j�U��
�d����#U΄���򴰥�&^Kz�ǰ��/_��aF�i�79�LƳ��YV\�ހ�����>����S>�&ψ ��)
��N��(�%8��&9�D#�Dq&[����N:����D&=��1����8���zq�3&̮ W��&$`��zRf���8��FxV�>�2B*��pnɗ|�{ԡ�����L��UF��+�I�m�`���2�����@�â�+�o+�	9��JqK}�υ!v�0�.`�sc�_-�����^����K\"тkK�JX9�_���BG������C��u��%��e��5��r_�<���\\7�$�;��R���{���#�&�É4�pP��^yB�s_�-�Q���)jl���<�h�`��Ǆ;@�KxO���o��:#�R�&�,�>��T�Hf.�as��v|e:�����Zy�A*�*���WX*��ɢH�O���_�Ю��Ǽ�}�t͉��0�
j���4>�U�e��?��	�!}-�(y/��_r6(iaxҳ�0�A�qZh��vN`c=���/#� ���`cм����x�>��}8�К�˾���%G�
͡%��:D@}�a5���daQ�h0+�a/@��0A�RV'I���9�����_���=��{��7��LU��tXD���+ۇl��خI���F��_�GrPF����LR�`��[���X|�}���ʒ]r9�<r5xxL�������q�@U�d��@���a��Fq$V�j�&��ox0u�^�n&ZB t�l��Y�7��!=~��
��y�Y?d`M�*>SP'�I���!2�fF�Ȅ,�Yb�C������#�K��"BJL��]<�9�yV�)���E��k�b"����T��P���JZ�lpĎ���|/P}w#h��x�l˓I։�,��G�WW��u�$���q�o��v�YK�d����ߧ��5v�]|�����ٷs���zo�䳛<���q����6~���]ݾ��4aqG�����@$<@n5��G��d�c��U�Y�p���1��VB����)H|�~b)M*�t�����q�R���I����<�Jk�&jHr-�����R��0���:՛Ґ�4�$�9�)3�P�[?�&:��K-m�1,��Ka?9r���������a���� Y����{K2tx��N��f5�m�-���J;��P�i`9e���&>j����Z��v`r@Y��$���ǰI�~��&)L7٦;��1̄�}�g�@���u�"��":���y���@�����Zf���&[a�A��y=<K_c���]R���yIY��kq��	B$��U���x��[��NA �Ú�a�:_/�sj�-8�}4S�5�K���x��������#�٤���{9�]2:��3�xش�ҥO!�|���@�/C�����i�f�2�N����^J��{'V�=��a��4�v�Y4m^���N䥠�ix�J�{0q�s��}�B����"�*�e�2�_OM��j�5������#8�ͥ[j-�e��0�lB\��� �[�^��~�f�_<�k�4֢W.�[Y\��bfX��s�[b�ʓ��;��*�
FA�\ }��I�R��P�4�uUh�x���ד���J���7���Mp��a��/^��LN�ϗ�Y<R�����d��g�`d;�R)��!���!�f�ӛ%E�m̔�� �FNCG�_`���Tmf��F:e6Qi�v$	�l�AB����J��i��9u.g�����fjؚz��{2#���N��q!_�˾����}���r��u�r)�ﴓg�,��Ò����q�n->�n�C�y�ҩDG���=y�a١�I���q����g�����B����e���%�#X�nufa���I���Œ��J\mH�����k5�uE��%�<�08b8g����K�$���<��,E@m��<�?,2 �����7�G�e��'��!�Ty�Í0=( x�17C�@>���J"��^o:����D��������g���˻��MSh-9���(����%0�s:%����sU~�$��bB��L(���c��mC�Z�e%	C�H��j:4��5���B[r�����Δ�i���UZ��kw%�ฃ`����]
�r��g4� /�s'��Dr��(oٺ���Mj��Q[[��8$�.B)����-xn��d��C���ї聏	^��iZb�:�vY�T/I�oJ5����@
&y��!���쐮s�C#�EHa+�_�b6҃�dK���H��2]��"�_�u��J�1.GM}�1�a�qTM��r���M��+���wV�P67-_�{�5��Yl��h�܋�X�ۍ�ݗv���0���M��AR2�+5�r��I���uυ��ݰ�Q�m���M��#7���m^?�T���z��@Y�0����}}�w̨�,���	.c�m��_ċ�-�ߛ��.�.�|Sx�^]4ZE����}���x� ܑ�2��s��ٱTh���I;�]^��@��U"�`r� ��r^	G9��~C�w�%ރ��x"aȴ�`VO�!�ҁ��B�YQ��Z�[�s|�._t�m�<i����9�J�w�Iտ�r!T	��Sڀ������NY���n��]����W��D^�1�]]���1b����ڷq$CG]�ka��ye�o��Y~}��s�6��_�2���yD��Sl�	{��P�RF9���NS�\�;y��(i��� [ �l�'��K��ϲ������T"e�FB�C_�1`���h�Q���֗����i'"�.��P����C�Y��Q�7��tB<�\�� h�C��C����7u]/uf��kv���\W}~�r�%L<5�	}'�P���|��8����y�t���M����v ���.�Ȝx�3�_���o����0�5�|Y뜏�%������������R���V��������v��G�Sl�Yu�ᶒ�3S&�L�� :R^��2��&{���˘[����_����ܳ�0cTi]�_+`�'M�?W4a�&��f/w�ػ��|�&�%�U�^AE��L`�T�`�LxĨo�Z*S�+�j��E�����ws�6`�ֽ�����v�i��������QB��LH2%ږʛ�}-����Qs�̔0h�8�+-��B.��u��	e�-)�hq30��1��������k����|�)l�z�Z�CU�b�T�6,�JXʌD{`�U�:G�\�XX[Gub��2��35�k��z���C���e��FD��F\�D��� �K�g�3�GvKJ��܄�,�������w�%�
Z�
&ҳ7.��/���4�>��hO���\� �"�b��)G��K�*:�;��gJVtN�$����x��dyKW�d��2R�j�$��Y�@[�D�I�z�Ҩv��\i��B��^�p�+�&��)=���JT��M����gk�����n<����l�?G� 9~y��_�l�I�(����9��AH �eN��\��j�:3&�����ͻ�/��D��Sy�����!���S�.��>��d�4�����C��lo�]~2;}dsF�������t��;��� _��e(z)l��҆Ld�ZW�H� ��S��*�U� ��������0��&�W'���G$#�0��Z�-�1n{����Ԗ(�5�}bG�M�Z�2�\���o�=61��C[��/�?��u����`Ӿ��e+���$;{�F�"S��n�� �$:P�:������3���bcyq>��Ѱ�c�,��'/'�7��P�`-
V6�_s�	,� 5� �D	�2��H״P�=����Ƙ��;n����u_�Hm]����)N���Y�r��PlE�i��/�,}��Z���.l�'�χ�Nr�NH��q>#�ۣ��ʨ&�I�l1���C�`,};��g=����wHd@}��g��4P����h.d��}����2��S(�S��p�� !��҉�M�@�L�U��pLUb��X���_��C7�_�E�/㎞T�S�5f .�ɾ�Bw��U%;��2K�D(�}�.��r�`ӡ��"�C眪��(o�O�y�R��	2��v��GQ�z�~!t��^��	��ߎs4=�d�Z��[��[��9K���5m��@M��;@���f[��Uݐw�֛�ђ�-���a��F�1��9}��y������|��^)���f��l��`J�*lAP�,��ouX�� �nS[X? �1Sn(t�J֑�z9����7=P�{�뗙�gd�Z�b�X� ��>��SQ�K�m9��������\-դsZ�\4y����tm;΅�$��J9�R��$dF�����r3���|��5$-4:ë`W �X��d� j��S�İ�pP�M�����I~ȩ"_ �ձ2����;�������f��'���[Q@Ư������7�ɧ؆Y8�Me�)4��L#"x4��Y�� 
4�X���ϩ�n����Vܱ�ŻD��8q�����!m{����xj�бapb�_0�C�~��pf�/yp&�� �I�����/W�� L%��ޏ�6;��Y����T��~��QO��|Ĉ�)����`�l�G�/B�Jn/OW�R�{�|h�I3�&W�Һr	Ա�}"�=�7�+y�V?I��T���Wv�g�4{Q�S{�nő�h@�u����Z%&т8��en���\a�lb-��kx<���O����V�8��@��hbxR�m���x ��CGmQ^IګxmsSa�A�!�rS�w��`�F�$0WzC*����#(�:��Cj��n��-����OAv[���l�@��t���Q�r�.�/����a9��o�z�5�"�9��T�o4�O+���l]}�R6˯�Ƈ��Ό#J"E\i>�T!��$R
��¤��$G&h�?�ϓ�":�C��d���Q:�IՓL��Sȏ0p@"�x�� �Jƈ��3�'����B���D`�����������$\�3w�T:nC�J�a&�>�z����'L�����]7�tl;V2��]�lǽ�am$��|z-B�ӄ�8>�t15��,i%ݨvNR>��1^^B��'M�߫�׍<x>�GJ�������8����H��P���h��v H��MƏ=�3aĥK� �f�*������8��Mb�"Z��F�����4(���Ý��m�-2�����_b�$�5
�����w&��h='�~A����$yVKd��!s���<!���e�:��c�D� '���+��$�9F���u�=c��B ��&Xlҩ���qD�w7I߶'c"b�QvI��ܗJl�:`�Z�*kJ���o,�ssP)���3�K���Y�}s ���-0ׂn��h�ϋ}���P�����dT3�'���1	�.�I=�v��ۧ🲌!ԭ8.#����`n���]��G��\wu�v�!A�ׄ�D��ڶ~!�K���3��Dܒl*��S���pwQ�8������օ<�^ޑ���7�T���iq�5��\�ۼe��`91*��e��|���#�Ҹ��f�!C�0B���@"�U{4�f�--���{S*(X��'�%7�ly����h����>ʗ��	����x&�f�q�ڡ�o�6B�C[9_� f���ˮ�qI:��
����oh�� �ِ�������~�JP���:�q;���6܆���^���M��Y��E�pQ/+1%oŘt�ی��	'c�P~ AG�Q1+7����S_�e���_�}�P2X���>�#��<Ʋ7금ܡ�0���B\�����){MS�p0�0���*�LQ��w��#Őڃ�E���1��B�� �%��.�jp4Yb"�JP�_��iP��j��
]n�$���FwSKh�/�>C$�j���&j�A��M�y>Cq�M`g,}T�ҦZ�E��̅n ��4�:pwm$|��1Fk�!h9��ZD?�<�;Wg���h�/�H�󱶰I:���,����B)�c\뾲m,�5���4�J1��<�6��� ��i��O�[�:����׵�Ԛe�3A�u���R��A	�ز�jAO�h��$GS�d�4g�ͧ[��=����&ɭ�IOH]��Ľн}����W|i7��l�����˿^��
/�N�7�$�)���x-��O�O���ュ��C�ߠ"2�OFZ.����z;��ά���&'Jt	g_HN��z8�]���Z��d�G��y����Bj��'��!�q�b�z�����ѐc�_tw�V�����t�M��n\�}��(��`b%݃d��/"R�s���Do�m�C���4s#�)����`��|��Cx�Ff�9`���T�n��p�v�yY�vd��"��2u��j����t%��i�`����š�l��2��]�TY�W�F�We;x#7�'J�/�*��Er~���=R;��sfq�[�)�"����^V��b�$��uz*c��ːm7l��z�|��^��c�"U}�Ho��ML���H��M�������\(P/D�1HߒK�*>�n�.�LVZ<�K�M�ye�TpƤ+��N�G�c�|�sX�xVuS� �<p&|��6m���!z�
��<�������g�mH/opNHg���&З�b�l#>�x�j=��bvn��^��6�sa"�am�jyz�C���*�4���zl�،$�IBd�d�_�;���F2��5��Qq�7�N_z��E6�Wx�P��v����w����\�;)D�g����߳΂��d�H3{��ד��zӌ�f�S�%�OEMA��F،�, �n��C+wUv�8��w�
��?���mĺ_h��d|xb.s�HđxP��%a�朒����hM�E������OO�bs�$�{ß8��IV�������w��-�R* ��o���m��3f��[0��������(�9Ø�DB;r��	��vx�G�a����Ⱈs^��48�!E&@x�����7w�%*���6����a��ߕ�_ؽ;4�h\�Rn�ؖ���8��"�k���������e�t�dJI�Z,���b�9ķ����R�1����W�\:sѼ֯NV�^a�W��(��M����0�_���\�+0�fe�ɲY��ǜ:�n�{���n�[������@�(�W�0�(��/hT� �/e�"geMg�r�ZҨ����::���R&��֌�#�� ^��m��\cT�����D�I���}I�FZZq�@�d�t�`��'�����#�'��/�쨻9Ԋ2�Z�� B$e�.���Y�Z�CJb�t�*�M&��o���z�`8�]�Z��V�T��Y���Z�ו�X�m�"�wʹ|<�=M�mҬ����x�}��S�)�'�ݱ$\Ϫ~W���Ύ�cB)��EE&�dsj�h׀NQ���:��c�R&��;2��-P^� 8��y����m������`���G+����CE+L7 8O�#N��v�LY�\���6�]2C��c��Y?�ٶ<Vְ�r�����N�� �^�᫔���ɰy?���L�!�}[Y���Ҷx*<�H�%黴<�O�[)j#b~���̑e�U���7#�XL�2ff��b�/�+�(w��#k�?E�|��%���&�4�,�ٞ��N�4s��?p�i���s����A���`�V�}������c�}��V��?Y�Ȣu�mP+�iG�C���򌇚IH���:�U�
�	Ce�-��>鱋��q�ϳ���,��X� ���*dx-�q��M��Ru� Y�?���\s��Nj������5��$�����W����iO�AU@1l6]u���Fot]>4g�K���N�5�L����'Ɛ��(�����KcA�4�^���)��	����t&=�|�� 9_}�[Pd���h*�(pR㝁7�LX��Т,	w��HЅ*��B3 ǲ���-.��!��}'$؂�O6p���>S^9�[0�
4��lzm����P�� A�,g^���dl��Uض�࢞��3����D������ކ�>g�wK���Q@R;Qx"������j�S��zSO�Ұ�I��N�m�T>�ە�KH����Adv8I�{_t� �Ӆ�M��WZR��Ӷ'��X�au8sibP`�����͏�:���0Z&��"��)��(5��*E�/b�P\Y�{p8j`�K�v��L�<y�!0�f|�)K�r�K�.�O,y��o�D;�۱�\X�4�͹f����<���sv���d)b�F���1%1��E��l��-q�c�X�a��n�ֿ���p�ѮmCUo`�ʲ�C>;�<S}�C}|x)��ю֊��2��CS�z.���g��j�h��_�s�p$��L�S?HD�i#߱i�*i?�԰p�����!㐵���+���|�s�#f���]W]sVS�(u��i�#"k|����r�>��*����q�b���Sh����ɂ}#�������Cs]<[%�����&�Y�+	�Im�j�y�r�J��ĥ�'H�2�j���p�{`/��P5#����7d�k�N�O4� �!F��P�~�1sdF�S�˧���[6__�7k���Qz�Xt���hsˬ�Ņ}"�_n}zj�ۏ��P���gѴ
���~�B {���aګnk�@�hż$�����t�Z��B<�$[e���߾(ŕ
������{��m��r�q�	���l����Dn/xn�����ӏ<ؗOӄ>����bͼ�W�eA�_d��7���֢��s$����ާSPb��G(��n>�?م�#�]y�8	�s��s@T6 &^�؋n���D�p�j��A֍������R⚑k�K��Pɛ�.��*j:\<�ź.��1��*�Ć��6����w��1��p�*�?�Z��.��#���|Lt�/z�a3?W��,>�o̮\¬ƨYV��ɲ��|��5���o8�y6m1������Kc����[�����zn�E��#/�B1��0`Yr� _�& K�58�m���X�I��q~s�?�)� �:�$�Uو90�y8���a������?����SA{UV�8/�o��/k.��Lb��t����fV%��h�3yj��I��׮�"���`,_�`g�q4�5Zt�4�.Gij�M�1��N*"��o�I�^;ޘ�������^Ԫa�����	���7�-�Y�Z�z�yϨh�����g��ӭ�T�,�48*�fOl�4��v����.�G�ȋ�����B	e#bҿ�p;�ȟ� ������f㳖N�$��G�(!�]y)���%�e��z�SO�����s���Td�����^^�}�1��x��z��a�v���N��`�K���^ې�V�aa�A{����[�ڦ�LD��`u|?"�k������	<O��� ���/7���k�<��3�Y>Y+�U���#�� ���VE"�%��Q��̫_,�'��%ʭ�i�"�{���/����2�!
��a����d�k�Z�dޑ���(v|Sa8'�L�^����q*|p���.�7��r@s*/,��;v�������D.|C�,ݐ�vs���H��csfnz?��WK6��K(;:m�?"u)q`��=M��F% �v���VQ�*M��k&vUAIZ#2��É����k�T?���:�@�#ĥ�+����?�$,e�����[�<�#��^���]�Ww�.%��O�Z	�՘����ݴ]���܎C�.�/ݹ�`��{�'�v 4�u�D�֧�>������:������I���e�$��K'T�Y�ZB�7T��/�g��$�mQ��;$�9�F>����1'�a�?]@FKALl�����>��F�c[\�B��n0���r�$%�D�q^V�����䎊�|C��PZ�yn*��vx��\�|���տ��7$e��#�"h���Ɖ�ϋ՜V��v��>�c~59�z	/*;g�9N�Vҫ�h��h�B/ǹ�o`���J�On�N7�*C����g�C��g�l����i��q��������<���U���C\d�M�DJ�e
��P�v����A+��%�g��L4ƱJ���N�ec��^��o'�v��1�P��-�e�����{���O������R�ʪ�B��yV����Df�Ql����WVujYxIX~e��C$/��d2���iz�`I �X�d�+�zWT'?0s�y�j�������+\>Nu���/��ؔ�5XJ~�\9�2�e(�f�蠹1��Y)l��X}�\U�\o��!nܓ��et9�I/:9��n�d�w;����3�!�瑳0��Y�;2��U=�����W&���Q�	Uh���@v�h���L�N���2���Z�ܐ5���ߒg���ߖA�H���Z>��>�d}Π��\�6�"y3�sl�R/f�l��MQ�ưr�o����%��9�D�=���#������	g"AR4k���,c�̔�>�]9*��hi�w����dQ�,!(���V���9d�}��nA��/*��o �h9��
�mٻ#N�t��ԂR��UG[�T��_����A�9�?������)F%��?y�l�S�gf�E~SX���mxRt��8U��;�O�� G\4��<���d���7Pjs.�uQd�#<��D6I|ԵgC�{'b]&�{�}Y���0� ]���{���+}�q�2U'��bNt��ʒ����6q^{?/W�k<0�� 
�W��/��\���e� ��ڮ�W�n��lI�.�)F~�ٜÎ����+����~q��馋�m���S��&��;:�*U ��U<�e ix#p>�i�Y#�]� ���v���m�N���Ë�d4����7]LD�li4"Z9y�ʰ�D��g��r]���j�t�=fs�I�sdN1�'x+E��(V%��_*�p��y᝗�c�d���^�Mc�s�d<�(�Tz��b��R�,���K��/����ͅǚ���#����Y�~_�*�w򩄻�����I<�������� Q�R#����`X�V4m�`bA�c�K�u�L�H}Y-��~GԂ9ZT�E�7]���� ����`<*-�9hG���K�!%&�.��͋g�e{���?&�r|0��7�v#��J�i�>�~!�kB��# ��?T�����	��EXQO �Z`���]�͒ ���-���ٯcu�!�k4񔩇����)��l�`�,c����s�F�n���~��%���iM=��!��h�Ky�jOשM��ke>tvXnF�9���g(�L}v�̒�9>=�?�H�lH���,8��	6HAv��Ӷ&y���٘��i��X��4�k?�j-�j���B�����������q�bq
��!��{��`���$�g����(*����=���ur��]H�X��x�G�'��G�ݛRC	�5��:⼽���qJ�[E�C�T�G��R�'y���<d-@������!�5Xr���ؖ��w��/��Y8|f�^D`ţ�^�v�l`������q��b#!!���g��Ò�~�xH$i��O�]6�%��-�fJn�
���L�ۺ�ĸ��
3��Vk�`�3��C�$��'x�<w(�^"�H���e���S(M�-z�l�%;=��2a�L(�pd�P�Ɏ^���B	�|���GeF�D�mA��C��Զ�9�[��Y�{1݁��߮A�N�R�����~7����M�(�z}�w� b�����9�t� ����زT�o4CǔQ�M���şc(����B�g��?`��
�Q��/� �?�6�~3?���>��@�;h��
1F��/2�y�U�ɞ1���,D3:������LOII
4[� 	�%��Z���1Y�E�:�7��C����_�5NLm�Ք$	�'6@gy�%$����'��*0����O�a�l�l���@�k�A�xZ�)���$54�m�t��P��[a���e���5�H���Ɗ�(�|V܃���a�yST�R�匝%h��Qƚ�Ѷ��X�e�b��mv�3
x�
�.�gD���O)\=X���^ʣI7@�_�k�蕒�n�Jr.����X=+�L�iM�8�	&�nS��βR�y�51*�~��tħ����,�gؖ�<����]��b�M����J ������eO��id�H=�ku��9�z���}��x%y��\k� � �\͸Q\R�:�)����u�, 7x-��P�P22�^ч���{�oYkA�	�(�Aa�w�!G��f{�3:�q�/y�=_h��&,ޠ�㦻;S���T�b��X�@ZнϷ���C�@5<���NV��~�+ǱD�iջ�{��q�"��A�Z��2ǲ4\v�ɺM%���tķ����!��hRQ攕¡��^�6:`��*%"������s��+�b@��L�'���;:P��-R�0È���o�� {9�DU
���[�%�)��:��~��@���1�Pl����*� �I8��	��{�Rj\����[�ґ.��k�׽V%Ôz���8x�/��R�.����P<+�Uol�J��<}�k�(t�Ǌ�9ز�������609\s�Q��GĩM���O� �G���Q��H���Z@�,��,`��{>�����J�b)�Ci</,~+�[��$�I�ვ1��Y���3-%K�Q�� �	�6Lo�kJH9.�����*c�e��|/�2Eи�Kh0���5��~i��Y�5��`|���T�1�ڳ��|%_��K�{I��U�>h�� n�����>A�X�E��J+-E��O�M������)#�&���Cc�MmR�ג���2�3�^�o�a������-t9q�Y��q�3R��/����o@���]w�r�1=3�j�k�B*?�E���������Z9���9�W�G������}�2�L1�L�7@ӔX�d5x��O�gUkg���n�5��Q��NaҐ�.f�A0�-��tMdI��Z�_���f๒���U8�Q�~��[@�/��G�_�z��=��E*�%��u"�U���0���& F�������s�Q����|$��ԣ+�N���3br͔�b}i������p�N�F^l��'fk��q���zzZ�3�������!&�����u��N)$�B��\�q������O��qQR����uq5�ϔ�Y ��螸�����,%/LXk���e�A����)��2���漣X�j��ޘ��[�-y����]�Uf�'8Թ!�nFuoK��]�N�l�v��{ß�!�3c�����]��4��E�*�* �6�>k-�:TA�~���I��P;e���h���nT 8ˁ�}��M,a�b���^�P��#���`��2�4}��|H��yΉ��f�q��i7}ΰ�	I��h�z��#'�fQ�T��Ӛ+��]g�-��fQ�u��,�����ަA�h���1���0����S1��RY��Q@�J����UP�¶}���`-�z9wSTiZ���!��:�\�6����1���4�50hBNGE�_O%t��1f����Wm��"�S�nђJ�����X�+�2Ka
�}8�Ɗu%�s8ᚇ�wh��Z�߿�_�-К�h�6/t������̌4��D.q`G@l�́�����6�{�D/ ��{n��0�29���ɳD7��#t�;H]�i8(<�3}�^��D.ѷ�z905�yI�E�>䈌�Z��S�����O.�|%���ɭ��Z�x*�AH�͕����ݓq1'��t�r�&��Ux[է�EnD���s/���C��To���������	����>(
�:���6,-��]��r��ё01�w7�&���vO�-�#�q&���	�z*�Vg��U(7�̡cDi�U�Q2a�Ҝ�e�c��e@� �����a /��9���~e��6�vOQNtc�r�A�ӿ�<��e�OT$	J�BB���7-�H���è�A9�sk��$$�&ш2՟�d^ZV'O����O�����:�`
���΂r��g�R���p�=E��D�q��-r���KO���B��A+��A��u��rsA/{��A�
��'m�E��ڃ�[��L�L�n��j$�ة@X�a����)���c�1��P�C�}�^R>`̷,!����+˕B�㩾X�����X�	c�wR���l�a�ڀ!�N���N�)#.�us\ ˄���;��� �}�=���Io~>cХ;+9�<����)��Mm/��z��YL-3X2/*2#�ja.3���pwV�0�V�'�rhñm?��7�)��L�a�9R�D��4T�4����u�l+'t�Z r0�(T�;f@G�P< o�����뮿3��ro%�b/�L_$B� ���,Μ��ssj��]Lif���M!�����,3OZ)&���P&�ae���OT$"*EZ��VV�ub}�8Ad�� ���T(��|a9h���{�7{�_�+[���-'s��<E���TC�qj�R�#(Vg2�d7{���,^'�kR8����I�H�֎�8x���U?eI#ς������f��e��03:��B�M���՞	y���+u�Tp���E����e�DhN2XM�� m�5�y���&|(zt���>؂a�B_�9sn9�m>�}]�n��j�feߴ��M
����}�Yd��!F�ѓ.��71�b	��[���9��m�M��)�x9wڒ29F��uW=���s���.4cU�NMp���!�mx���x*ЀUK	�ny�(;�7�S�ʆ���F�ឍı��lA�mD�k�M�72�aۛ;���L�F;�������%���N�>��֛�ԙ�X���~|�;��� D�(�:Aw�b�fq�@�Sp�T��J���fS��.���3J�:'��V�)w~��0�xo��iϠ ����G��H
"��=�i{����L�� ���j���@\eV{O��P���qE�w#��ZRS��5�E�E�` H;4�g���b��E�߱�g*�Ch�@��J�B�LvI_���.cp̃}� ���<�8S�D�}�F��]xw�V��缓��A�[���fy}:m�d7���3�]��b�ef��:|�C�q���ױ��E'��Ə�}F���3�L��RyB�+�5C@��"����)Fr��8��3~/\8��g4��@8���u��\��)�s�XQ�4E��q:�kS����f,G��rѥl��-����C�eSGK�w�We,GX�/�06����rSK��9��)\���?Ċ;(X���b��ëlI݅��6YK�.	��j�NJ:��d�l��4z�(h���\�u-.�>C/����eI�V*���h��r�􆢖$3���L�Y_�D�^���
�@��F�y�V2�Qʹ;4w�@*��H�B�8%-���Q�Q�{�}d?%��~y�	��qrEA/$0=;�����Ӂ�����BGO?zHA((.P D��d�S�n{�u=�2a֞>�aH�3u�9�w�B�طs4%Rtb�m_�L������8hG�v�ل��;V�=L�F��mg��
L< �O�1�@�1
o��|�W��tR��:�H���{�R�x5DB5�@؅����}F�	2��m�	3�c�he��iڧ��fF�׬'�F��_'�x8K>I�LyI�ϣ�ٓQe�#t��%���k��i�ZPS���
Z����o��F�nb���β�� '��Z�b�6&�b��V�E��Z��H� 
+n�"��ꠋno]*�=�`�A����]�+��"������4���ke�Q��W��,X�st�o��[q��N�P�Q}�B49�^/޲tb/r-B7AU���\r�w�Yf�-t��b�������E��A��y.7r�0Ƞ{�p��D���;)��q��o_3�%z�Ǻ���C$�;��Z}���TY�>�.��,���y.둖(���k�u�5V$��+O6������źu�Q�g�����:�OJSҐ��o�Y:�+��[
B�H�briv���q�=�)���~�:�;]�أɷ���!���ŏF]�D0���l���m�����shڕ���΢�,�v��`l�7a�hftp��t�i�`��5��"�ˣ?��/�T��Y=p�R�܌>����
��MHt���}�����5��]�\l�"�k~cJ�͖ �0��6�r� �A��GWQ�����jS$�N�pׁw3�#�Vk�q
1���2�tvK���ʹ1M-ąF�п�>�q�$����'�ֹ���(@���[�B֍�~����V(󨿊"�?Pi���޼11�N���^;M=kL�������6�v�6���-i'mRO?�\�kr?��(�m�T.��H&z.|F̵��'����S��}-M�ݐ7���Us��,L�-1P���&U �+X�>q�.΄aMW�&�������3N���U9�+����G�W"o���I�t�Rp�X��>�����^ӏ�(AШm9�7_2 V��#���R̴����`�@��΁��;H
����E��D5
�}m�N!+4�j�m���A���ǵk���H���:��Æ���Z�-�柟#S �BLߨb��vR'B���c�e�6@52�ː�.)�A�>�6h h[Od�q�9��90�N�͇�aܗ� :Y�����o��Ƹֆ��� ��4A/� �\�.%�(������������92���W�-���=�F���v��ܛ���6�D��0D3�~�<��$�/l��;���v�.����Ѐ�FXaK�ZօSш,��~���A����L�[�^B��(x^,
��\#��M3�q�����IL�ۛ��I����[+up=P���ؚƉ��.��f.�i���x"(u��:s&9e�k|���!)�w࢕ ���P|_]	� �9��W
�6_T)���sD��&'�[�a� �����:+_���RĈ�MgyJR������hG�;�ɪhQxP���A�=��K����'P(�'����+ѻ� ��Z�aD�v[�k_���D�[u?*9�ln�����)���S�UC"3�
C�<R���Y��5U'�����]/`q�硷}�n�Ƥ��h�+��_I�p(�+7C��
��]��h�:�p��d���Hl��e��z��mN���]-�؞�t�W���h���T��Ih�����\��P�kf�m��}�5��(U��&J�C�
iXʉ�5"�t�?0l� ��3�$�	?�F%vZ}��<s�����+6S;E�G�NV<������9D)p�Nz�b$�a9���ǳ�/N��Z���N��2`��Y��8�{%�7*����2~�����vh9LQ�Mqh?3z&��6Nb��qvG��~q���ۄn)G�ś�W�w� n/O�q�i�x�\oe�1}e =q�6�aV������tt7�6
�̯v�-�*��Gc�-'˜B0r���	J8 �J��[�H�Ϣޮp3S�����K�?���T}��$J�ƃ���?� x�v��%�e���+�-���t�f�"���6�ho�u��7)o[2��ք���oڳ~i5
ǣ�eR�m ­
�,[�va�����Z��e�ChR�M���2x����>m�G�U�i���"t��*��ɫ��W�tz���\�Fx�F��� 4vX�vN����Ud!���q�J�Ô�޴u7�@���*)\PX�Z��H��_ ��ز�`�sU����/ӊLao!Ŭ�e]�g��u��}Ʀ�~W'ո�����Sˑ�'��@�`ٿ�l�w����F��/)Q�\[{kž@7u���KIqB5�813y �I�jg?�Z0�S1�Z����eԾ�%_��1����LJN��sp80�c�C5�t��>�s-�6�^H��
������k�|�=T+�-(�O�����h6�U�c�Gϓ��~�'|��+�@q�p�ג3!�=}�^JT�������6g�����ѷ�'��_\l)���|��!!�
L�m�c�՟
�g��a}̛�Ŗ���/�2�T`�d���=�����{w�3L])��2����:��2m��P"rJdk�T�bz_J�Ic>���x��yH�ǋd;^90����֭�e��4M���Qȷ��o�#�����q5����J'����x+�b����C*�͢�J�l�iٴ\,v�W(Ώ�"�<��8�.�y�O}��R�����6;�e4e(j�'��]��B�3�Dz<��ه��+���?g� ��]<˜�����r�2#I/��Q+��#�:Ol4��iה����Ћ��cx�{+�"�W=�Y���x�
 ���T�婾#-;d\�-������m�����*��=C�M^7�~������v�D�� ���@�r���Scw�hS��2*ս3���I!�����Ⱥz%Q��'�8��j_�~.�=3�5|��%�$���j�H�gyN\F� A�z���tZ�K4o�~��F�n�Q����h���Q��/���H4��b���8@�����Ǘ��?��%]�iŘ^�~����F! Z�ʏ<g��<�Q�Λ��C�Q;�ُB�p�ޔ���4��X~�XF��������C������w]�6�P՗*���&�,��E:�*UV�DJj��Z��cQ�/�X�ߖ�v��:��[~��%ݥ��_\����UU_��}�[U��V��ڢ���nCqu�l�Ab����C�K�:�~�K�T'�i�`E��Q���db�"^�hթ}��p��O�ѭ�k�'��-JL��ڪ��:�]������h���Qs�c��n�����	��F �c*�d�8�q��&o)�/���H��'��A��ѫ�����с��G���"$�/V�IC�`櫼0&��ib>�x���Om����d�Z�!o��z�,�\�ǋ;`K��#@� ���2�9���Ӡ�qKF��|A3&ʫ����UW�����t��&�6C�5��²���o�;��J�2�by��c��"�_��wN�m8j[��1�و}��[#�yҐ�cY��m?�Ř�,Mz��H}H��k���!�I�>-�~�b���JL�a��z�EU��c�Q݇W�;�Tfc�a�6�xҶ���&�ly�~�5_��ʷVj a;gUL� ן���fq���İ�_R_��*�5k��Z�:Ή��=ōQ]�|A�<����%��9ڑ��	�O
;�[���/J���l�Kb>zG�i����ۛ���o��kc0;l�W��֥����D�$*�U�˘�!�% ӆT.��u��ܔM���Enz��ҧit�?Ja&F�?�&�+3:15���n�=I�i����5D}�{��(�����CcHY9j���dHIo��T�~#*kK��9lX�@�,��q�ѤaB�������|����L�,'��3˖%��M�H�v=D�hاk�HV��D�����1�k�HuA>S6}���������I�Jq#y�CpT��b�"���T�U��-�K��@�7�x���8�ZO�}-�X���=7�Z�z�K��mJ/�V$��?$̳Ʌt�<W���"��G��F��z%��������=|V�a��壨�:���"��XgW��r��!!Q	��G���RO*���;C�>����|E�:}�o�*Ur1���rڜ �I��ңB�!����0�Ӄ�b�c��������H���G�R-Ǽ�u�:���f�w>`[1^���&�茗�?5���� ��fؐ���������2�*�r�#����7�W�=8e1��g�v���w4�ZG���(ِ%�)4�iZ��<���y�c����R�Ʉ��|TW�4�$V��.�t�_x�'h�\�P^oj1�X�������{��V�nO>�"ITOA����*������BV��U�_����IB�+l{�x3ԑ�iC\�M&��T�(��t*Io���s���)ř��y�_���Ġ,o%��i儥0i��F�&#G�|�󃻇]<d�MK�nU���{}���/�7�'5��1>'��(t�@��#�iF��2k&�I� ���G��	�TzjD��F�q�eZw ���O��GO<�E��l��Eg|}�������ب M����5b:^E�P
�����u���>�G0��ԿW.)�|�>w�W���J��o�QkWjk�q���r�gI㊌1�,�o����@�d�,T9�����L	�w��K�ϰ:0;���	����5��s�
v�l�6a�PL��m���CRz�����<����}*����\^�4>�iL��͇���ë��T)���~A?�ZY�����]��Pn&��Sp@��B+F?U�N����ӍM$ި��W�j��&��/�G"j��h���gX�3��0�Ƥ@v�D���s�Z�b�����Y���j������퀃1���S��� 6��h���-�d��h�ZT �GsBa��A�XWx��fdϠ�wg�_�X�-�s�gQ�(R������|�i��eE�?�^.�S���u �'�ax���mj�.ե$�ۜ����4�oADBN�E�a���/'�&�w�Bߡ�<�t��^��T�P�)��2��� a9ۏ9Ȫc{�uE�[�1X��'���*����ᛦC��/3G�Qm��{�J��� ��^P�Ԡ�����BLӂe���M����C$�-xؾd��'C���Bd���y7���0��� 66�CGty�5�l�Ӹ>d���V��ɷ�G8L��K
I�ǆ	� r�.�N�{�h�J��b�
I)q�@t"Y���צ%,��Y��N\g��2�d�������1;���V��V���!U���M�>V�pF��b�e����wR��H��|<Sz]��Ek�1�H`L�Z{t��R�����G�����&Y���S,���-�e��V����.�Q��s~�V+)��aww��J��C���\9͎鶹B�x���S~`��IN&�L���u�˒��;��`��p�m�W+�o����)��Ɨr���h=�˸b��\T��UE�[�>�ׂ[2���		#�e�1M%�Is&��W�()��C�I�Xub �)?��<���@��\R-0i���}���i^�n=Kz�v-�
��^�~\V����2��ݦ�ԭ��"�oY����!hx'-o@D�\�>�c�E6y煍<�޾ԣҳ�D��¸�$If4O��\=5�|��O�8,ҍu�6c��T��?���o��WY]� �|��;R���#�Y��]m}�=�FG�Q&�D�k�@'�x�v��$����)6W"�O�-`��q����v�6����
��u�������G��v��\�u�0�M�f�����~�Q��g�@rP�֐�W�5�V"�L���@�e:���(��N�"�Q�;�Meƈf��XZ4hF�~%��B�e���C���hM�BDܸI����������_y1�c�!�Ivmt��w��|S�F�����cц���4�\E �]��ac���+�!bӆ8����0����
��b�39�\@���QbhTw��f!���ӣ2�'�����B��������,�
m>�Q/ ��F�F��Ta���N̥����@�j�֌��������(��B�&�J-r�P���_�r	,�8��ؿL9	�;9$7�@V
K�աu��Ҁ���dJT�Q�J����@���";�Z�	�!M|����D
�����4����������9lN�@;�y�Wl.��}�j��|و���-ڡ&jR�w}�?��i��2)��fN�<떻7�����I됝Z+)6���t|���h�v�z��K�fW#����Ju(�$� \��a���xG\����Y�X^�&�k�6�ނO�t$��4�^̚�ݷ�^n%��r�ψ�W� �/��wʑ�M�A���[��V��;�(� 蘻�<��aD
uSy���?��z]>)�����̉����b|��Tm,0ZeϾu���g:z�TZ�T������)��rL�\uք������AD"!y%�Uؼ���V(�� ��[���턟� t��Ij)�'"/�2� �L!�p;�+�%Oka}�k��uI��yI}W�m3�;ZV�=��G�Ђ�r<�ߜ���^������h��� V�K.p�ˆٴ0V���� �_f����9�<��|�c�F	��ǜ���ij��l!�̪.�P.�[��ʯ�!M<��n�{[��'�
z�O���h��0�I5�H%l`�Y����Gk�):9��Ē�}TS�P�S9�y����R���c��j���Vg�� l������j]�ީ���$�Xo^���V�=ſ�V�������k��(h��9ϖ���FLH��"ج��=�w�7ܸx��>�W�p=y�^$o�k�U�����E~�cl$��1��ć��s|�@�FB�&W@u!3wj�ǰZ�7�����@vp#M�1}[���6�N�[p�{&��_YnE�U�@ѫ
I�%M ����0��V{�nOcŉ�"��P2��|"y��ێ�=�D#�F�?����-�D� ��ר���IwY���v}O�6U\�uנ��j�r����>��ɋM%r��[���a����Q�[�=���e��0��v��Z�y��<�W�S��!V�Mg/j%B���/k֝�R���f�-W�'-���s��Y4Z�+��Cy�u�/p��W�
N��&�AgU�Px�_�8��q[�n%�Bǿ$���"K��f�m�T��^A5͙WH"��,${Q.�7�%��֮Ŋ�-��;�=T� 0p�L�31A������ߟ�p����d 3w{շ�b\��T���<VMB���4�O�'��js�sf�<��@�;:��%�.\�[�D�5"�ih����vWѩ�f;��۲AB��m}r���>�	g��F�y#��]n[%Y����Tb�C˛�܁��U~�;L��	�W2||�w ���!���j�o�]P���ZꕨS!ge�,�h�h���S,T�Zɥ(�;vH_�H�F2��_4�!��б$&���-���0����γW����zs�偂�r9wVk^����Ĥ��d�B����JV�U��č�ͪ+��óY��3�)P8�S^3^���5��i4��ٓ���SC�P��^�u�@i��v�[b�f�Z>[� �g�-��[cz�����ޙ���O\�����:�8.�d,��=%�$����C<�p��Q��,�=��>�Zx��1��ٮ?��E���2J��T�`C'�Y�c�� K��E�#���j�
z��"�:�'��5z�z*�iE���)�R?�{-�뼜���G�Ub��d�#�UQ@<���¼��"e)ˊ�cuD�%ܥ�<-.�J/e�G�>�H�F��Fp�ef��ְ�V�2�?}�݉4�L���S��з+�gy��8̃�#��yOyC7�&_�/4A:�/���QW_��ȋ�v_�iKH�=���q5�}UI-t�M�:�ɋ�e�Ƶ@g<�25|Y��X�]MnL��#��O_1N�o�[��y���Z���d)!�<����ig�����k���T;�tz*�n9�χ���1�~��Olϥ��6�������s�g(+Ԕqí�tQ�~��l�$�/<V|��M���˜�E<���,�TB%��}��gv2��|�Td4��V*~,,o7n���s옉��j�d�����	ʥ� D��'�NZJ����_�a]*1J֏w@�W���0���ٶ4��:r��$mD�$z
��U��j��Yt �����.M�-O�����X�p��X`Z�?gR�m�ٷ^e'@����푼�/N�5�0?�G\�ü��L�u�Q�T��%^�$�f�����;�PI��Şjf���0�8�����L�H��~\ԝ��H�8+�k��%-�_3�JC��#��E�/N���Q�n��˸Al�e�v�VE���p��i?GB\Z�p.4���eć��p�P���ځ}�l7?1�OƘ�Aλ8��������dG���B$�
�L6Ӌ�Z�9N
���l@���BG��*��N�K�n�H��sj-E^aؼ��o�xK >@r��cL��P����'�nԿ��N(��M?��r��!��Pm:}�Y��%JP��}��&^�X/�t��[�1w��xQANF�D�E��i����QӜK�G ��@�Y�ϗ�ݽ2�x���8��_�We��
ٰ�NN$���AO�}�p�kHD��2as��-Xq1��WCD5�fG��j��,���!�0���j�����?*�P��L6nL��\��->2�0���{�r�Eg<�����`�˹��%� �Ǹ�����g�Bw�����9�_�Q�D"���.�e*�E�2�-�^\.���Ҝ��"��� ����nWʧ,��πW�q�R4���$�i�@`'9��c��^�P���å��re=��k*!RDa�-1���]#im֪�>���eU�Z�M|Y���&^GF.:c�ːè��6t8w^J�g�
A�n����w\�j��q�m��i&uM���ল}��B4�f>�L��Iyn�9 򩦧��1��20_'�~ƍ�z!Kr��oҗ��Oq�.|���U�hϰ��$4Jl,�m�i�Gÿ⳶�ˊ���=�M3��@��c�%����Ùd.NMq�9��L}:y�\<�2�R�z;ˍiuG�j�O7��Q�%�S	�T-�y�3�{��䶪ga0(i�k�O0(�0k��T9�%$ ]�AX5� �U�<�|����+�}E�=M 6ي��<��^�w��Ήǌ�eAg�&�95�@�ǆ|�A{�S�޼�؜5����������,3��V�ly�R}Эa(�P`�ѻ�0�����~E�T��UU>j�:[��'��in]�ɔB���������[k;���Y�x\��o%�;��ͅ���]���,�قD��5����ʠ�F�p�k�!���ϝK廉zZÆq]�E�P��ۄؖ�ſ��B0�x�|�"�X��fح�Ǩv�Z��V(�(3������6�d�K��d���֤*te��)�i7`O$`��kX��p(HZ�x�Ѷ9�5ţ�
��c n��n�� d�4��P�f���\�}ko�@s���T�㡲�TX����B�BZ2�7Vi 4�{>q��b�e�eM��� 1�z���i0gU��+�4;S'�"1
�ʐ�ri��Aҕ�C!�����"����QO���E(l6����$^ Z���2�߻�/啹�	P��(r�+3�#��dX��a�6ᩭXp�o���4֑UTĬ�����_��B#�u���v`	v���`cT��J��w��:b]��B�'܇h#��aF�&��.(aq6���Y֫�X셫_!�[r]�K1�H�Hy�Tz�%�У��(J����I�2�jŗ>�Q\�"t=Rl�_��7؞㲊�3�znA�ű�5������e��S�7��.�����Q4���]A�/��ܜW|����%_#�	���}��g��QAA��^u�q�D���%�8��&��H7X{��I�
��"or�"���VШ���e���61��5��%�)��_H�ާr*p�h��LE����}=��wq���Aa�H�y���A��C��w��^��+P�l��H�pjD��$H��+�-�Kv��r��[�V�#Y[y��O&�NFX?P.S���^���Z��Ew�ڂq:��֌`��#�[5ڿU��.�RJ��XX@���HT�����J��ue",�@a���!��ߍ�镞��_.�&�f��.W���7�����s�jx��
�9�����q�R�|C�:�=��T�B-맣$�w<�RQA�t�Zit���7%vo
�ԐS�e�.
d��_E��xW.N��������u���"+����GV��u�eΫ3{㼊2;�(E�ִ�R���XU��F���U Bnc:��N�fx�)��uI^P-�����N�lL[�_S؍�/ڧ^�z�T�cб�%4���-w����Cb��!��rfך�1��+c~�H���뇊;�/���3:�{���� ˤI�[m�{��ZdK�7Kk5~��ɍ%R��M����D<�G ��g��f|������I!�y��̕���/u��d*�6\%��$r9%��R��FBr���:vO��=��i9
8��|�k	;���2�"�yR�=M��g��u�ۿ_�Z_ �;듕��-��Q�UM���Pn� ޙs��]�^N�&%aWF��nG��c2�5�r��1g��1)X=�bq|��r�1�$��?��2��8�����a�yDh>���<��Ќ�A}k�$j`�D�;�Axֺpg�Mh�O��n��Ţa�*��.dA/���c�߆w�{𛍥���m�iů�!�ûy��k�VZ�f@��##����A�"�|��g��!�)5�K4Mc���S�LOR�4C\��~��b���D �h��g��M����vU7����94�
"($����9�є��h	�kPRrZ�3��n�
ۉz�����0p���� ��I�[T�+�/�ډ���S��~Tz;�#W�E	E�9�� R��:�P�v�nX���B^�����Mb$j5ɭ�}-�o�Ɯǭ�d��1fn��8�',�W���3P����(�J��V��˓��-�W�cfZ�kI�� �~7����a4���Oݞ�0���1�K��/�,+�h�������ݬ���Ūq���� �Lf�ղ���/W��6��������nx�h�`��#����ɅfL���fq�黨A	� �}0>���B�O�D�V� о�܌�BP2c��U�$�Fo���w�}�Q�ۃ�����[o�&_������\�q�N{�Q	f������u� �&T�����N�s�7;/
��,���P=d�$��3y&�D��t�˘ժ�Hu1��쩕��O�*j����\�1�z)_6��$�HoU�m2�f}|<DE��>�����1��B���������=M�t�>C���Ñh&�X�4��~y)՚�tZk]A�͋R8TUu�/&�+��A҂9+ 	�y8i='��͡�<�'xA����2m�����ą�W��A�Q{��[I��8�"UM�p���Om�J�2S$B�q`�#�#@��8	-��Ɣ��G/="��������Y��M%�� �bP�n��k9�e'R#M��G��Je��.�M��td�m�X��{�Cw o�t$~�ڡC�CH��C�Mo�XZX���w��qS�^;���+e�4+i �xjX���{:�($mV��l���l��>���U,��[�/3���"]c}.4��s�dM[�\�Fr\}�lUmdyXc�rq���g����zi�a"�L�b��wq�e%�}���;A��$m���2�l�i�-�
	X�9��VI�_��\d��)��j{���郞T_6ܻz�
���l5l@Ji������W� ͉(��y�k���ѕ(��~�-�d�v�_,�����x�[^�����Q�*�^�ܿs#��������h>��&�%�dϣ������!𾦒�`X\�s71(�cc^��.�Ŭ	ђ�M��n�&�@��Ȉ���4�>�2�bژ=�#1�=)bOH�9��LL/y�̅�b(��?��`:�m���Ư�&7ƴ�J��HeY�x�.��Z�͏R,�~�Y�����8*dT���vO�1���e��kм�F�=ߦ��Rٟ/����v�~�S��>�YF��b���I�Ak���0�@��AɮZ���ڳ��T��f=L�*9Q�@h���煨�[A�����ζ�ל�h~����Uvqm�c8��8v�a�u���,��x"@%m�����8�Q�C�Ľ헕e��?FHl���&��!�PE ���x3gN��'�_�U�-��#EaT��Vt|LPh��Z�Q����vX皘�`�
�u�����Ԑ�W��y�n/L؃�r�Y�7?�lJ�CT�m����ӏ�:/�֘mp�R��Jx�C�������Ԇ�H/a<ԍ�
��Uk�C���"-�W���i쒭F�v^�yv��E��]�s����ۇ�}�"}p1Љ�Rm��[���Ѡڻ�Uˇ�t<�o��و>�ivLk�X�%Y�p�t�0z�HrI,w��ZQ0�,�+=]��Tk
�Z�:��=@Va@ځ(�+ςU����S�)$���u^�J`�}����c\�5կ/�8
�����fN3�\s�Gs2��l�T���_Qp�er7��SK�V=;@��q��+=1l������"��=�q��8Z×X
V�ǥH����'t!8)�~SyU��F�+�?*ĩh 軃����?���G�����/s��xdZW���T�6>��>�5��Sj6�Z��D��.���O;�В�#�.-��0��:�L���Փ�W��F��JbrV��gZF����$�%#���Iԡá�����D����9nF�D�em�i�'Jf�'���:2���I���m��jq�}0�E��fd&i�ɖf>;��}@��½,k���֪�如���v�-�Vt��	�$ڷ�����"c������+����|M�D2j�|�t�v��8�Ky '}B����	Rò,� }�bӚ-�ÆK�dzۿ_ [�#>��3�����X2�93�g�(���4ck鳋`���r��a��ǙA��t)`��]���[>�I�܄qnT�_3sUE��~�ZE���l*ڂ�?T���V~��pxi���\�Lt���}!��3|	>iOV�QBJj-�M��pA�x&�;�����$�&@�1uw�v�4yB6dT�q�]�� �l~��d
+(�u�l�X�a������� ��p:�
����,U��Y�Dk�����*�d��.����3�{Z<W��{E��\�������?`��:0-MfX�R�r+D�v>L����*/��2��l��_\�ZJ��JvҀԆg�s�9=��r�6����[3�@�/���9��V��gtevp���̗�]�P���	mp!iK)�B�����8����85��S���ps�n(((v�����.Xd5#�޾���=���H��h��W���:W^m��v����j��;l%*}�a�!�hH�L��	)ܵG��@5Iȣ��nZ�����W���Q�ˡ鮲W�H-�Ŋ��sޚ@���`ͫӇ�>ܒq��H��iEY�_*�o>İ�X2l����1�O��P��2�tɽ��֏�|������_#?��A�U��)��}��M���Xg���1�5�|v��e3v<$ <�E�9�u�����Ü!�;��<L<��!qE�Z�t�ka��V���BM�@X��ӍĴ�,2"��-"��@��:�}�}�C*���{����4X`;���׫���T2"��j5Wp1�T��Ԩ�/Ӟ�k�҄qJX���g�4H�t���_�1��)W�D�.תl��I�#/��D�07�:x�嵻��e��v�Lb�[���r/3@E����r�6�}�/o�6?&򲸫X���,��p�a��-�J�w�U,򀾅��Eۓ3wO�Y<W��X�>�6��A~�3c8P�Xړ��F}](�k�"ئ�[�\���u���8�re�M��E۟м��QfM/����'��i=R�|���v�l�.���YP��2]�Pu�
��\bH	�Hk�,/���LL���+X3
��o�c��]˅$�n�X0/I����'����A��\roaZH�/u��`����&��?߹$�\���S�3�gB�[x��#�[5`AV?����
qTadl��[�[PG�;:��f�z����C���$TR��קp"�H3��F��?�q����%������ߍ���B�N�K�C���$����Ӓ��������&[��0+�ܕ<����pM���WsG�"��/80OG�1W�w{t��#�;�ùu�Tg�������e�FK"ƣ7㕶��Nx�&��J�
�I3�g�U��h{m�I�olPו"�MO�I�����6��J���d@�za,+=,r�=�W� ᝒº����0-4p��q,����@�A2T:��|=�	k�̸��=Z.�,R�;�����1*}X�(�ۿd���~_�vA�l�*�$��	̵g�0��Zp`�r.,�O�Vm����*���/_4G++�έy2T$�sYE�c6���� ����8�B��rOB�%��K���^�l�'�e�o�cx#�|-�i��g����Bl@�<ԫ�~wG���_�
	Ƿ�gؔV�6�.,�N�_�?J���f�_OlR>$������F�X�b��m[��%#̬� >�B��?=k1)�~�oFqO�O�>@oZ>n�Pbz�j��<�}tX��!��S��vKR;����Y��I1u7h_4"7+n�'%�rr���z�R�*�]j�c7x��|����q��le�!x���k<
&`��,��� �4IM^���Jg$!C}Шwb����'s�&�vX��GB�N5�דl��CtP9},_l��a ��#9q46�$n�@ ݤ�i.+Q�D�=ǣ�"�++�.���k�����O�o �5^W?��ߟ��X�W��wB�K#��[÷�b���c��UHq�Yq���W���j<"���r�>�����&�ɇ����y�U������t���B��xip�f��uӸ?�׬P���ώ6��c��������SRu?,�Z��������&�<�L�+��4�S�:�0�����o~6����3������:����"�%}�y!�K�8���|�Xu�xɃC���R��
�]���J�O(���~���|_�3Dph�-��y�#+�}5��D��r�f����"�9������G��yI�Syc�f[���u0�>q z���m�_���`�S�Y8�e`949�^X����ut�])�JOA�l	�UyLBw��mȲHC�� ����l�.�����G�����ǝ�k����`�+ʤ�2��ϳr�]��0v��_�c/@�f��������;$?Hl��o�/� ~��#�B&�n!�o*����QQd�.�*>�p�r��<A~���Q��*�!�@��j�;��@uP;	�ǜ�Nn)Y-�\F�U9�#W�h�H�k������9�q�ռ���]���)'�gA�g�s�VF��`���`Hjc���)$=�B�w5&�!��k�+�(����j�����jW�\:�����J-��/;dm�`��NE�lYk�LV�R����,q؏JR�)i�v�K@x�]��	��-�k����+kSuɾ�*B`�`�o�C�Ӄ/lr�S]!�f�O��1Y�BL�"���O�re\��z�5�\����1��Џ����fy�a|��%��{��6cܮ�q�����i�',����F���lq�4������7P��-�	+�x�J��vir��/�m^Q�.�v�	�|PŰ�l@�%��w��P�$wH���AN�CcS���!���eAlG7cu����-u���C��1���e����������.iV���1]�>�$&`�Sd��g���`k��A�E��x����rzE�y4>ޚ��Ѐ��c������	�#.��Q��q�J#,n�p�h^����O_	6n��&�U$���o�$!M繞ԏo�T�*�A�eu�6j,����h��u��!��[�<��d6����~9�z�>;���
~p�B5� �KOe_ܚ1h܈��o�'�#�x�~��b��'2	wv
��L"�+k��?��v@� �y��kI�[A����/P�7ӮzwSe*,��c��[��9�"���ߢ+IX�򌼤��Og��p�w<��4����F�0����3�ڿܚP��/mhQl��B}���[@�|�	қ�~�[L���9��F�2Á&u
�.�Ss�+7�2�039qL_h�T��=�V��5����Ȑ���5Jz#�0�ĸ��2R��2�ܴ���?�O��h7!-+j;�)~�b9�i�k��G�/q��9�9%����R4��G�$�K��n�3-g�ϺVt�̩"�)@x	�Tĵ1$�G���ڈS:]{t�G�L
S�tDa����$���*^��^K����Ol�C�n܊��g.�h�w.�|���������E�Ì���_ΪB^�װ����3<\b��ە�]$D�����_OO�?8�?n���i����|���O2kJ��=�}�Fp;�<y��.���� b�+M��� Es�@2�m���"�ҧx+!qE ��5|I�?8�-·_^��b���|1�����M�?��H3W6��J	f�Gm�jJ;:ύ�[h�b6�7B��x�_}jV�;��h�S��=��	���'S@��Ud�3>0� �����V/w,� g��ÂOo}��B�D�N'Hb�'����r��{_����bzt�]A��cߔ��W�O���G���D���iF5K���x�t�.mfmG&�_�3j{wK�¯5���6c��9ޟ�wN����
���qn8�5��Hp`u}�I�p��z-{g��+�'�N~��*_���Sw]L)�������;$�ſ�{��oǩ���/�j8��E�*\8�.��W`��^�^�G���k��Z�w22k��a��_��S��<Ա9���G;K��J����gN)G� ����NA�!Jλg�i=�r�d�$�����[4B7I���Uz��M}��Ԃ�j�o Z
z�ɜ^��Ni�U	���Щ9�'t���2�,\m���	$H��
�
566�/�V�[��(mj������ʬۨ\����U�I<��
ݿ�̑�۹���y��uH`kS���%qr�zg$�rY�'������paރXk�y9�l�8��K$,���]Z�]�,�iwʸ��&��ϙ��5,��ˋ��p�&[I$ٻ__m�s��� ���`Ӱ��N�o������6��TU����G�Y"�rJ�Vk01&]��}�	xb>"�|��Ě	��ܑ�.��1���Y�� 1�uR�2�P�T��{F�H�b4�]�ơ[�Q/Jʓ�D�ɨ��̭���+9��e���8�:CF9��� X�&�(:���;6��R4�S����Z��"ɓ�9�
�)��]�����y� �lJ`^}C�LRH�}
�Ę���l.��{��������������.���ᨡ� �`�&۔�ke�	��UD��g]�=/��Z���!��|��n>I�@~J�K��`?`���vj������\��c�o��n���Zٳig�t�qR��Xdy@�`��@s:6Ar8i�dbC����YmO~��Ҡ���T=݆�Ak�1����nY9WŴ��".,5�:?��v���H׈�L_7_+������jd-�uoN��9z�"����C�� ����DDh��5���Sּ����i�D��W�菘aw��{ ~M�%��9J���2j?f�1TJ6B?B?z�0�=�|�ri���V����ݔӶ� ��W��[�>9��G�F
G�o9;t���'����oG'���m׾���띣��� ǻ68�g �!�D��P��^�̶J�E����H.]�4(�,^�7M�.](m	%�Xp�1����^�"EЌT�[炩��Vj;�p�G���,&��Z8���ۿ�%<��ւZ4<��G�7���BDe���9u�l�L'��ˊ�rUQR]��?yG ��-�׉gn�HR��	��(��5�ϑ�������hJ�R3+�q8b���ρ����
}��=��-�)A��_�vh\�e�r�����'���͚_;d7�q*Hl��5��u5��2S��8,��F^��(��EM�#h�q� F�u�#d���M$D�q���m7��,�X��rZ�Do�2k���X�X��xA��6�2�D>�6�׼��[l��y�i�u�]Y'����f^����z�_�O���e���<V��.4D���~w�͛H��������?]���E.gH�8���	~��Q�A՜����j5=�e�A��F���Ct.a��#U��"f͗&����ѷ�ٚ#K�
n��ą��Ő2�4X*I���oO��Ҩ?ʟ3�dS3�������	�?B�>Oڇ%Q�����)*�4���q^NE=խ́Qں%k,��=	�7:��� �����,�� uM��ɺ3��V����E�*2�.������+�k�w,�k��&�zB�⧹��c��-&��cp���c���(Țg��j�-�8��Q�D�e�>1��pϽvub����a<��zC	������q���u��k[�����y�&����6�iB�߲\�����?�r%X9'UoϞ6��Wn ���e͐K�Hq&i��	�z�8���=����;�����@��^Y��@N��^��{q��~��"��كY�\EE�V�d%�p:ӊ�X��}�t��'#|Ob�3Ssi&3?#k��4�(%<������=&��It�:����X>O�v��9X$�~}5��}/������g�qq��0�3��mgFV���%��O{{{�ۄ�Mp�ܑUm^���&#pG�(�K�Rkf��@y�O�3���!.#r1;���1W����EM��\\s0�z�$���PΫ��k��봀rXc^3��G���FS�F�Y͟����@���V<��EMH�H�1��+�����Mג�J��k�%��a�'ey���b�&ܲFUS�)Wͫ�d����4Y�a����[c#~p�S��mlG>U1�����C�f�5G�7a�RuǼ�rU6���8�:����q���M�9��ݹDa�]���Pb�����L3_K:si�����O���v�����.������X�p��8��V�j���n�2k�8'��\}@}f�5^��4�5����qo�#�������/_	��Uؗ��B�WU(YC��2����?[�t�Rz	��9�p�(�D��;��5�(^��
<���лo,h
�*�V����R��ɹL�PPK��U/)�L|��� b�bG��1l|���HlX�a8��»-� �:^�<����P��g�8��ea����]$�ſG�4�ư\��N���=�[�0ٶ_�� �U�( �!����|�t���p�vk�P�XU�X~<8�FyHE�H�33����f~.r�	��-��&�g�oQ^܋��9դ�Xj��Z�w(K�����p	�M�m���$��W���;���4f�	@�u�Գ�aq�]e�j�'��;�G�!҅`/=]!���QdJ��̍�����.jY�{�7�;�^��A�/r��x��s�TN_bX�	9���h�#XaM��nL��4���[_�n�����qƠ)��1Hv�&����B�;H�/s������%�J����N1j�� �&	xB@�A��7�r�y�w�>��9a�^m~Ȃ��P3����8#�X�� &���;�N�;�Փ�g�J������A���z�k� �*�ʢ|d19~�y!��n��[˶��Mw��0�Jf�N��R����ɏ�ٌQ��Vi(���Tb�n�D�1GHh�M���ζ��d|�9RG�^Q�!n��� $��R,��G礬N�Q��T�7Y�gf�6e�b�㕣8g5$�|��C~��2�������\8������MȞ���'�ncqm, ��X�"n'{�%P���@�r~��?��j�������j�p*�}��@�6��d� �ۚ�>`����}"����+/1��ՙ�}�u%Ԃ̕�֖֥���
TV���;����I;.�����Y��lz��y��H�sn�ϓ͋'g.���JV�]�)fX)�5j_<��n;��'�-��g�(��s��b_�z�|/�r�O�UĘ���$�w�`FW��b��oSH� �]gZ����.�(��3�damʿ�?��s:���Lo_��n�OFji6�9x��[�0��{�B4m���ځfR\�<�]��I[�^C�'$�6_r!i�L~i���:�)F�
��P�!M`ԥa�a��V�D�Q7@C�pb�d�M+�� {L勣��>LAm1�zͬTOa�"�~Xi�6$�;�}�r+؟�|x�{�*�/Z��X������Xx�6���,lQ�kI{�+/UE�F`@�t,�8� �SLO����G�;!I��В$��ę0��9?w� -v(�2~���a�� �Oj�[��;��&������j�RL����W���0��$MBH�Q}h�v���FO��Ț�~5I3��*�8}�S�m����)#U̯��@�(i�+�5 ���
;7��ny��~@ܧ�(�(���Ћ�w�-�ȾW#} �@�����0z�=�2�
�3���d���7��J�������c۰������Q�Q���@S��SIJ�� oq>�u�rJ�)���v�@�%D�Ҕw�H��j��F��_���}�z����E8"�}��+e��D���GnQ��V5v������+�ΙϽ|����h���-��@�I�+�}��H��iv���m������x��8s�NF��z��4(��|0��>#�{�Ka���ҏ�,�=�D�}s�>R^T����_B�ra�þ�������a(T�9�!�y� J&���E<A�7�,S��켶)\Y���P��mV�q{��4-="��:���4vN�u���↙n�W3�O�e(��H �$?�������� A�F)�"
$��\��gvYZ?��N�;���l򠓉�㇏	TD�ë�K�2�	.d[W���zRl� i3���e�`ޤ	�F튃�)?G#T2_�|Ǥ���#eE�C�/g��=�vr��O�� �=y�R�0f=�®�1H���j]��ZC�pT��J q���m���{��c�*m��S��12�����ݖ|�|�4��R��@#ۭv�LI-	k��G���
�0b�3ȶFme[���Y�?Y>��$����S��:�2���hb���V]��
�.YJ9�a(�#Z'����z^V���70�ҿ�OP,Thb۪> �9O�̾x_aִ�SMA��*C8���GRH��^��X�GAC��O3����oBp�Է ��q��]X���d�}R��
�Ie��M��k��K��x���.~��S��-3�K�b:�!�[`�d�5�SE��5�+��k���y������ߨ���ʯ��Z+Q����\���������?�aa��;�W[�����-��	`2��s��gd2w�Q�ኅL[�ޙ N. �]e��?�Q�e�0�����U��iDSf�c^r��1#�me�ئ��E-L���+Oݧ��uXyS� �@%[�V^�`#b���/r�UDd�dq4���٤��ތכ�Y�w�'?�St(��%���)/��c&������sI��*񬳇����<�,A��96n��*��f�mz�I��廜������䗫f�Ђ]ƫ�l{FRi�G��]�r���_Eɨ�@��4ջ8�|�;,ڒLL���P�#�WJX�-Oe���P�|��e^u�޿�i�yR����dx�� ���I�[�IZ2V"u���M⮹uɆw�^����g���J�]Z] l�)z��e����9���Us��dOf��3 Չ�ʵ����s�����"�-7�_�u��ac��|�+��a���M�dbw_��{��wɁ;� ����hY��HPe6����D��ǞBJH����������c��z�?!BTȻ3�\)��L�h�F��98��h��)�ݛC��Ub=�O�eit���Hv���ANIi�=0�4�S�n�b׬x�	FQ����6�ж9�^��n��hH�A�#�Z4վ2���6����@Qn������Ep~�� =7�������94�Ew/��T�x�%��8�zY�-T�x:���2�]���X%zRt	F� ��U �̯�f"��<u
8�ɋ���Ʀkՠ�㵥|��i!��F���C�,�֠��v򢻭�m�T�C����]�T�g@2�×&0�[7�m��z�c��"���8��AYa�1Mx�Ec��Ǝ�QOs�$�U���ᱞ�R��5��L��3x5$�IW:�h� ���Ej&������:#�UǁETh�7Y�Q
�l��ƛ���G�Q6��f�����=�ɦ��D�����x�A	�Q_�~�i/���&�8�tK��Y��K>�����4�r6Ze����0ad`�wV���i�*���:�@]�GkV�+�i�%΋ �lT�c�f��������A��ǝ>	��P��]$�i҂��ڝUgч�J��WÃ2�9>�Bn�����*�$D�b�	ͫ�4���D�c�QL�)�4���[2O��vtL��;a������p�i���V�9Х�Y�������w=xG�p2���a^C��8��R�:g	6�6�O%�@��FT�Gls�>�u��b��\
�غ0@.G���jX��B�H�3t�u����=�zoV���V��T��9p7rt�k�u�Y#�}�*+W���;|'�.�Qਤ�P�El��!�+\��?�P�d(k��
��j�DaO��	Z���V��\+�����l�Ւ[��=㠪��*o���6Q�59��j�3JA9���U"�|��0t3�;TF���&o��~*����u�:Z\��y�~�w�=��+�'��ÿ�R��f����m�B�i�cW�m�?3�R�%=�n���
�2�|%$�j�=R�f����pё%���^S51�"�DF'J�%3���F#�m	A�?��c��T'^T^ݢ��8'�[�i����;�n�!��q�����lC�%�=k��MXm���o]ܩ{����@�'�21��;WO���B�tE
>��4�!����������F�\_�ǫ�'<������.ng)��w����������q���J���9�B�!A��E����D�[8#���7���R4c@w�fSM
_�I����&.K�z�ƶ�r� xU]5���z]g���c{��t�'X/S�c8�'Y/�n9�M�mqF�,r����۝��3���v8�UW�׻�TE>X�h2��s��x�x�� ٓc��X_g�i3��a}X�5�a�@���r.�u�*A0�̕J��:z�vO����T��i{�JD%����(�:�U(Q��ԑC�'������/�?�D��
�*��=a�m|.���f:���1\��N�.�L*c���{p��]���냼v�T|���NL�u:9�3�=H�hN��w`�j_���zR�i ����rH[w	� U�	��\����V���?L��������*��@s�Ŋ@GRW�qɝ0����V�n��6.|�c\�4�X�u�"%�JJ�(�� c�n��x�۝T��7�]|�>��#��e�c0WO���
T��۔�����?jK3O2#˫��F�{E�^���~�=���H$:� qג��>��b(�a�2��7���f�'(a#�hg�_{�麾v�A!@��:bAP��/��݁�����_������E"M+<b]f�X���8*�pc��0�䮯���L�\�	NS���K���ǆ^�Y�}�/� �~��@�b��K� n�i��9�-��|��V%���#t���;�?df�5�H�B�L+az��qj��t���������;8�]�<X`��#	^a�:/E��jgJ�9��<ƊK�I�r��;_���d�����@(�Ł�T/���c���l��HI�[�M��z����WfV�� ����
̙�E���?��E��I��v��$�����&�����Q�Ր0�������0yz'����zْ��Ζ@�� ��i@V�EN��3(t����G,�x���!]	�?��ۧ��%�Š�U9�t��p��#��C�N�U�QG5��(��&���!V �c�Y(8j�j�ZῨ�����)�^¡-��"���\l�����J�o'���d�zѴ��H.�6�+^�r�W�A�&�]W��b�ۿ:/���Q� �ʜ
�34� M ����������|��r���O�	�(�&��c�1���}q6�s�E��ͅ]��|�G [��<��-j�zI9�qǿ�����0r ���_�l�𷬥�'t̡���m�*���d|�{�.K��%��ꀶ��&=�͋'�!x��G1d�7l�3ķ�W���!��H��98��|{��eMw�!#Ǆ�Z`���-�2��W��SH��D����1���L��Ըz�}�L,V2�O�KCjM������5I` ��1%|;�S���􁳋�y!i��:A�tn ��������v^�^�x�<s���o��{�/��lbȷ-]/�6f떴��ǭ�R����c.�cl��L},�wKJ�ԗj͹5,�G"R�������4�ԕ�1����:V����sc�#�� >4�ɺA$��X9lOL���������2iT�]�\`�5\�Z�S����^�������+"W�m�JN�ͫLu*��DX��b 94��hΛ�Af�h�p�h�8�>ǧ4B�P���u��l�0���g�w���|����Z��)����0s]0t������!���q��W�Cj]7���U;��9R�������
�ኙܮ�������9��|���J[Bm����a1nS1�b>ֳ1b�f�!@0)�V��ܖ0�·�=u	�4����W39��?
�\mk&J+L�@��1�b��f/�(:!��R9#���ф 4���кb>�����o�L�7S�2u(�׬�&�{����ܤT�M{u��n(�6����q�[��F}$.����@�����t*���?�ą�N��YY�������1b��>���u�ｺ��M�ωN>N\
X�~��kE;BbS�n,���o~���mt��bI'o���w�C�+釸�R�x�����ڗ��zS6��+E�t��;g[J��g8� ۠S-��'�4���ԝC���{�~��Ұ8�QLⳒ�B{>ToC-Q��	�!L9�|\���<�%�b�0Fѵ�=IM����Z�-/��,��������?X0�������� j��gZq���vE��8����5�1�WL�4�����~�����˭�Q�k�y�C���@t4��
�Y�3�d�R�ubj[�{$v�BZ��z�	ޙ�RȆP��?A���w�A�P>��ݵ�����4Z�][�c-��c� �2F�C��_v�❗��d���!N+� ��Dc��T	�5\-�<W8j'q�v��(��4�
�	6�^�[�#�Oi�@?�1<��R�T��6��-�x(�L��<6�I�D���1��6�� �}��K��k��L�~xQ�p�O���)C�mSd%��WY�9JQ���
�0��R\r#�x����M�g������L#��]�-�l�X�E�}X� �ٺ��'�X�.KE����DԋP�E蔺���*�7�� ��gl���c֎�����IWfsh��<�N�k�8�[���g����%����>Q�Ɨ:���ݸ�=�h�-�?58�X.#����ں89#�U�Ќ>*ܑ|ϭmW['Xc�ih4^~�	�S�G��I���XJ�!~���8�uI���S����z�8�JM-a	8q�8qwu<��f��zy��#�ȴ�
S�i?*�c$�3�|A�=�I��s<�vid���0��%HKs|��0�����s�A�n��P-A2}��w�\L���Iv�)��mr}��H�{;�?;�e+0�z+&�3���-?� �k|q}��,��ω�=haN%t�AW������s`��A:9�j��nj��4�������[n39���#��I����������@�<�o�TE&a�q
��>t����༻�r�j}�4{,ZalQ��C�b���L�~��8Fwg*&}g���ȏ@&��h"�=��iτ^�6:����&��@j���+�=���\>�z�,��U�����_�$\�V���t��.�
�i�-4�֖A��=�xJi�SB&�INpt��:`���]�ހF�R����4DZ�cڷ�����,T���=�������ᩐ%T!J�5b�mPCf]57���7����29-�}��ؗ/�$�f�/��0��IRX��L4W�|PfV�3w�\v�Eˡ�*h �Po�>a	�l(r���Փ5�1���$�59
��}���	^���s��$��V�g��sp�ע�8w"}��'�Y��W[X�yEm.�!E�\��j�$�A�. �z����)ͫ�g&bԉ��[
e�9~b�������c��'T��F��J���~WQ䭱H?&�j-�z�DX��nah�NJOh�e����h1k�[�'u7��A�1���!������9j[]�5��B� ��@m���~�zdy�J�vއ�W��Xtư��&_	�nx������h�/d�B
G��7��*Z~���4 X��҆���2V�Q>
�@�n�7�lԠb~XZK�*cBH/=M*:�9ʼZ���UM t	�.GU�LN�9N�|��?B�_ܩ𣌔\�z�,��)�c�@}Adj+�q�6�O�4�-�Il�[3�� ��&�	D^aSi|ܮ�q���Z�x���-�W�����	��5�'�iR�~��%��ˬG�����>��Ð��O���L:n��&)jcʁ���m�����(:x��}>SU�����D�i�M����/�R{�[J�S�>�|���=;�?�cO���t%b^
L� �ߕ����Kj]Z�Kxj3���{��/�4��]��ը@VWE����M��O\����˓���`��;�S㶗z&pc��zF��l�#�EX���Ck����V��JB��B��3D	#i���Oj��{.W����!�(���B�&��v�Ϝ�ԣ���c����x�М;W�������v��qy9�o^��%�~�f`�C�`�����3�<��8��f"k����
M`D߫�I�7|�D��7��O`Q�
0��H�Ӧ�o�D�^��*�����m�ކXv�ӣɋ�1C+1��(�Q<��H^ڳۦ�V�d���}�=cś�˅i)�d��a��&�o�A�(g��%/��X��gg�Q �}	�����~f�غ��z0��T����q`��P+��+��x>����T�h�|���g-&���8w"qB��N[�?[����*��2��/`?���s��4��Jɬ�m�3������3<��M��8������!��p����<�x�o����!u�['P]!���-?#ǁGr%�
-.�L��c�����@Ebс��	��9���;Z�涣��(��_���z���+�����`���W��Ӈ��ǤP9<��BT"���>~!�$Jj#����Sϲ��@���hK#ʢ���?��>��e�Q��8_��lև�ظPcz�{
Zh�/��ۄl&#N��	��s�O5�5m�֫�Y��!���mUX��2��!��p�L��L�c���.N�u1��3� .n��"��v�!������'�Z�V�F�������K;]�����7ӗz���?�7ܛO?��4���#];�Q��Oؒ�k�ɨ0aAe��q:7���!�ɳv���6��Z�m���=[}��6AK�i�(��]Mc�%��VC}'�<���?���\�YD�o���S�KH��z��dQ�"���4F:?�k_'��L�:3��&|:X�AWi�N��}@Y>��|�({�@oK�I-i�t˽�>�m=HF9Mة�\�k��6iJ���{�Ҁz?�F��9��24�MW�_E.���X��U��t=	p�`�f�v�yii@�)�����l_��@�t���̓�����,B+�F� (YO/4{JԱ:��ϕ��41�
6P���!�Ml�ED�r&"]P��)W����坕n�1)��~��<:8���U9�]�3��EwWq-L=�qcc֐���[w���6Fl��~j��#n2�NG+8�E�ɶ���b\�iM������e���bv\ij;>ȫo���)>m�y��Ϸ�x>��ҙL���O����M!�<Ԙ܈�n��	�z_�	�J�-ub ������d��{`�)1�\yu�L�d��f��%H��}�K����o�tp��]
 G����z]��!C�r�d-��`vc����o\z)�6�^�?�=���0�� Լ���̹�LDϸBݥr��WD��Œ�BLW?�2�>���� ���l+H���V�q��	qT%{��������)d$�Ҕw���o
��[��4�%��*�Y�[�X��~�(̭��!>A,MC=2ST �7�/H�p��Kz���K_�a75=�%��߅��һ?�Q"�����h+�Y�*���s|.K�nkv��y��S��V��9�I�pZ>�B�.��,|�sQ_;�5�ᠵ��L�m��vy�R��I�j�_��ח��='�P
�OУr��2�<��k�^o�۹a�v��;��<G���B�(�H�')j�ጥ�.꫰"�3��Y�(�p
%�[����r���.	ĕ�	(�<�ւ��Q�J�}L�I)�� rL�ɯ����d��+Yћ�I~Q��~�	פ������Ɩ(�ש��/�a�"�������oc�����*����o���J�m�}E��M����!�
�����_�� �Mi&ms)��H6L<��H����j�bj\�	f*P�/Mȏ���>O����۲95𒢔O~dO�d�L ��H�`����[��E�ʂR�� �x�"1�(��:�2��D�Y�eX2��1&�G)���"��P�2��e���!k*�XU��.|�;>� �o�M�f�Xr"wn:hdetԊ)r�\�q�dOf���r+%+�kLr�+D�po3��պ�T cpJ��?�3 �8�ocb��ѳ��M�'d�>��%��gӓ�&'�pj��r�$���L~)�Ke�Y�.��J8TYm���hc����69^��w�9��1�N�ކY��j#�U�rѴAAD=��#��u!�7Q[I3��Q��ꖕ\�2�jd%�E#Y��9����a�2j̡M��P��0�U�������oS�/^������J�p�Dܡ�$�%mA�ǉ�y$ԸZ�-���IG��(
����i��C庤��s{]��b�y؎�]�O��ш�-��*�[�5�r�Qb�C/'0m�6+Z���4�h
dV��zA&�������ZA�Y��4��/�E��*>�]Y���^��% o��)T���-���[���\�23���v5��V�r!"�ݳ��t�&����<�{ ��u��f¥�V�r���(��3���)s�ST�����~*��7�A�n^��.l��[��NdBL,{9&U�?C1ISO�tybC��Πl��!j�8b}ȕ��K�ao�E礭�O~=l_~A��C�+��!>����w���ws�7>��YK �kTv��N>�o�����
ɍ!��1�'0��(��h��7+��Ȭ�;�S`s�R��L`%f��	Q���>�&�U�6n+�&��i��5�(r��6�:y��:摩"�c��9�3�� �!q��A7�1Ht��s�����8;�qS$��A9�-�G
��^�<N[;�R�3lv�.F�@xFs�e�}/45x��r���BZ�Β�mL(Q���O�J�P.��W��Cf�Ϭ��������=�/A�\�
������$��ܰ��5I.w:���Ȭ+��uk��q����|����w�9�N�h��cp~k�Ιg
1�e^I�.�pD�^P���Ӎ�� �m�~��'���P4��c��\��|d�^���etHf/�td�+�xP�{�K�2[��&�OVW&^��!�	���b,-\���(����/�L�w���zT�.���(Sd��<F�,��;�rfa1/���w )��1l��#�Z[L���;8<EN��w��r��!�l��1��$t�{�}�}�q���U�?M�x�~w��՝ڧl����9X��Md��%���c^��K���)��bzDީʝ����gB�D��ê��C��n�q��|��X �\�2���nPJ�"c�!˅ъ��B��V'�9��.΅�߮S���-n��=����;�}�+�I�@�1Oց��P�@P�%��#h�'O^��'^c����m�>��e|�V!��^��my?�!R��5����:��쀹Mu�1���8�A�򉈄�T��,�I$�̤9�sO�.`
�{�o[�]"��Z��+5����I�Dz����Z\"���F��_�˂�<���^a�*�Nփ,Dm �k��kY<Z�B��:xەQz��a�`U���2�U*���c ���ey�}�K���fM��+b������d�;F(�B�ZK�H�oͿ�Z�:�f��-*5��*�ݩk�qW�Z;0D�$dR$pM^�����y$�+`wyB���	�D������F�:�)�e��|�ǻ�����:������bIm�y�׼\u�0Uj�!����<r��Lp����w�$�|�$w�a~I��/X$;
C����r���9J�/ܛJ1��v��@�� 'b��L�L}�uhI�I`���P	��i� 7�aK`�Ο_f�������+`����k���V���US\��B��pwd�[<���8��G�6�9^(~S���ف��ǂ鷚;,�{������ǔ_�����d�\Yj@r~����dt��i��xa3�[���5C䳟�o��)�T����=���WL60�7ZM,/֗�/Ձ:Eϕ]>����N*�(ǡ^4��g��~vp�1��!d��y������D��l�����n���ѥ^r�W|0�+衧� j+�P�QJ��J�"ΐ��(,��q��l]7�����C�%���p�F�B�0�?�&���3�����k6c�����N�^�r{i<��W��Ds���lE��ӌN���E'�N���~ւ(ﺨ{w`!�S�"Ȯ\�M�t�pi��>7Ɔ)�C\��s!��K��z�P-���j�藊�Js�Xe�έn��̉�4�!�0'P�y�#!䘻l^�}�+�/C%)�(_���\r_K?.����3Z3C} �\��d���%�A�@UE<4�؇���ҿ�ԜeX�|��Vd���.����uh��O��`��ޛA>UW�j<��
¨}b�!M�]a䢆��b�CS<{�!�ܣ>�,ħms�=����Gv�h<���<�� [��Əd傘�'�\<���B�q�6�|��s;�HC�>���9(��[�F�/d�a�.��A��.d��� *�����W��<�ӻ��+���Op�"m�C�4�(7��S�ԪU��� ڰ�ddA��H�43v;Cb��l���1��̰<�/<���F�����Η"��3�%��d�W�Ԙ`	H�Zר�J՞���z� Q���f�S�(��<Up��x�DF��c$w;#H+��%NJu��F���4)5�A(0($����?��)���!�+K3�0��x� =�f�H6 6�H>>��o���i�FuU��<?�������9��qxZ�QJ/p�N"�K�В��d�<O0J�Ƌ�猏U��lc��r^M�C`J`�b�r���ʏr^0��R��\}�u��R���,�as������3$s�;?M4A���^m��UDNy
��~�u-���x�\+J������v�K9ߣ���i3��C.664��նd���(���Bk�Γ7)��g�线7�0c�F :���P�8 �'�����M�)mzNr�@�bL^g��<�(��Z�Oh:��ޖ`H(�2��Lb'߉{2�FQc ��G+M��-���14#+����%"�͗�����L#S�����ցaSHэT�UK��s#rF ����d;�0��6�8��u(k$k�"21^�MG`�.��f�xnNF���?��Dr�I"-�!��F���}�j?;Z�0�9�^�"�յ�`=�����Fԯ�_Ӵ��a����&������V�gw_��� ��[��X��Pi��;m�L~	nF-�/�K� �_���֜|��C)��5$W�)S�s�O�1����`�k�=�}=ev=|	�~sxPA�\��;�<�"�n_@ �k��ŏUORM�����,� ���'"���~�o��-=��[����6cU��C�����[�f<x���Ѽ��¥sC�ԗu)cY`��g�Erc��8�h��f9mħ2H�USYi��.9��&Dseh��9���ӎ�\����e���,z0�h�%��o�TT��,���:x�~�����i��"g���CG�B]5���*j`�y��|�|������'��	7:�hz �	)YFcԪxN.Y;p�����}��Hx�-�7��-�HĨ��N�P�Z�y)[�: 6�h7�~���H1�.>�^�WcY�����+���������֩T��%��A ����IŎ�z�h%y�>b�lrFڑ��iW'��-f��d)�.�;���Gb� Nh�'c����:��e�'����D��{����J�i]i��@ԓ��9��̽3��b���H�RŠ5���R:jQ�	�<kZJ����J9���|�e,�_\�Vw	k�YQ��<J �>�hԣ��Y��-�ͻ��e?��2?�+��#)�����x��x]F�"�ݗ�N���O�:|u�?�	�40Q�Hr�v�kM��{��{��9��A����=��si..�P��@�]{��$�)�.����6z��#�z�h��%�F�< \��D���zq����mg 2Ґ�d��Ѷf�f^+��7#���%X�--q}�p#[�U�~=�P�EӇ;�u\W ��SO�E1�����"���A.�xl�oR���{�\�I��k#�z\#��ta\���(����3��x�o���Cd\�o~ ���k`�� "��G�!�����w�S:L&�H���r��PX�~ry$��PΪ��>,�B��ݑ������RI�;o�
|��S�?���X�Q���	"�,"�+b�����3`�>P��H!�lA�4A����Z�/�;��4&���Da7���Qt��[�8�y���������!�*Q(�R�ɘ��}
��2ԫ�.��П�p�o���Y�	I� ð01���X�{�s� \��y�EG�G�����8$�*_���=G���q�3S�Q&`��|��]��<�cq^н�&X:\�to	�2=��/wM�l�k?�|@مT�3�ާ��9���,�p�S��s� P�,ֿKR���3����4��@��c8[�欯n!|a�uK����	����0"?�@��ss�Z��0v�!g�%Ԝ���*R/��ƄB�A׉٩:��	_��/b�Jr�~8�v#�|\��/��%�͛t��L~��`S7X$�>v�;��r�w-D�\f��S����i��z<��O��lY]]����&��FG%��n6?-�.�G*��$���±��+�#�C ��)z4mV%�nwַQ����q��I��&{�jR�r�6�ى�
��y�����8L����v��O�.�$-������ב#3Oxl.oQ8�˫�>P
haD���)8�Ye���0JH��t'T_p�{~�F�W�\��N����2/��f�Lo�k��ʻ�OJc�7(i��w���#��q̋�`��qt�:|��j��`9Yz�=����Nbz�cLB�*�(z��9.d;�&o��3� ����U��ԃ>��E;ت|g��2ߝUԁ�~��	Y_ ]���uE1P���FE� A��|�3�d��ğ~&X��d~������d���喐�~nۖ���jނ�|�z^V��n�����KRݮP�L��8�� �9w��nD�P�	l+W�PI�A�*[��D^�xnr�LpkW��%����-���� �i7����}z�����x�]%&O0�G�<*P�� Fo�a`�®e�D��J⚳�8�]^��r*��dV�M���S�8Jf���z������l!�d@�:��Q��{l��u�21
I;��*9��j�E�wg��ކ�c�X�&�ӛ�����ڗ�jK��-פ�C�n��(J���cZμ���Xץ�bJ|2u��uKVڧ���~�.��c"���R��3�Y�wBD�W֯�n襼��]�?����EE��3�3L�+o�!���K�z�7�~�����p�9 �RZ3��{��N����ʩB��~v��\��fC�Q�N�(,�5 S�X����<�w��r�R�Ot��\QF���D�x���{��������u�l�"����O��Όi��+��\���N��Ri5^���n/�2y�]��e{�E��
�r�|O������"9��a�Ɗ�]�kNR��#�7�}l1yc�r�N����a��Y��D����?1��yM�HRT�SOӌ�Ħ�j�p��W$X\vnC�7/����O�Έ�餾���(�sV0��S�P�59�+�9M�H�W8���>����U3	a�H�B�X6e$MlP�%�!��yJSL����QOW�z$m����G3�6�e�AȓDJLV����@xԮ [� �������e���CV#��-��4nbG�D�C(:��2y'hV�o.U�QS���#<�w���q״\	#E�88���)
�g�FRy��̂�eo��Tݟv�G�$'�Ձ&��iת�?.��G6�2�Z��õxO�X��D�����9ccr4���Y���s�/z��P��@�c��_�
��_Q,�}�8�Ks)��2�����K�[��E�����ÙZK65�X���-h(�BY���R����MC��ت�?2\^\�S��3�'�5f�ۆ�r|�c|��;�*���v�V�?AI��˭�r������ɳ	|�=�8a2��3w�a���E6s���ui�yO�	x�p�U���>-Wx�Q���6�v�gWZ��p��8H������8�:s0�����ė��i5�e�2lT�m�2IK�-�q��/�1�N�ۀ�m��H�;�X_������]f�!�nd�{/Q���R ��V�!	z��]Ah~���$Wv��Տ�kS#�d�\�G�|!�VH�������j���3Ȑ��-��QW�T?!&9�6��(��Y]�Ͼ�g�>Պ�q��{�~���]�Ĥ>YI�"��т���g�؃���^�������ɓ/^�฽ɰ3Fn9�l�<�n����F���6a9	.�%�tC��7T�A0��9x��C��3l�E���	|����5-��ɥW;>3��ʟ�Ii4su�cV~��X�T�H0�'��#��s �g�s�S��$�� ���;�B혨a}�\���LE� S4��,����V�a�����p)y�}:KK��5�)��Mj�|��߆�Gb��i\|�տ���'�}N�: �S�Bt��1�6 ~L�,�;K�X�VZ*��6���뽻>����a����>��;[m�0uoX��E|�	�oH >���	X �1I�קIl�1ƈf7�GH�����)h���|q@F4X�[�7*FJ�d�5*�c��.�/)�zN`��q�ɾ��o�f!�ף��tN~�$q�	��Tl�އ%bL�V}#ģ�V��ׯ��Dy<7Z��vL���Gz��!�YhO���5�fȔ׬��+�;,vk��
��-�Q�Pt�Ш����Q拭=(���Jj2�
��U?��[RG&tݘ�෶�ߙǑG�0<SW�;�A�sb��l��=�kX*��#ٔ1� �؇L���mǒU���r*���]r����.k���+��w;�*Փ��3O�ˑ��|ϩ��j�m���d�� �"�[G�m Z/�
SI8�Q$�sP/�%V'�2u�#t�/��/��������"�.6I�(���Ј1]oc�6aCص2�t��/7��x�fj��	����N��<-��o!Am�y���Ɗ�/І���V�r�ݫ?�~�5ϥ��:�'�x���_@����
�������ѫm��9�Ju2�E#�>]�^c'o����2W:���[�������<�6����zl��9N��K@}*X���";�������/��	+ygT����[C���CO2f5���ぬ�|��$�J�(g��y�B�b�.M��^�~��w�4�ɳFQ���/�e�-V��Č�?`��ʫҕ��%�h�%�0Vͽ2EU �0��Ր�k�xœcé��b5��_�&`C��.�k=�Z��S+fscI��=��X�J�u��A%AW)B��T��c�.X�0�z2��p�N��;�A�~^�v�#ոV���04���'�+$��\����n��d���T"m�u���T�h��#l�K�H������S�4o�F�%��� ��#q�>��҉���@Ʌ�&ܔ�ϒ��-n;�5)ώG�ӈ��8�E.�hTEUѻ�c"3��j�H��*·�y��>i��r\����^��8�U�_���{�ue��'��3ʗ^�P�����k=Lui�⎢��x�6n���~ҏ��y��>�V��`k:�0�D�J&�7�j�R �@�I;^��'>�� �d�M�Tq�/��3� 0���*�!�P�]Ml5|2c�+�P�ɜ�Y#��%����{|x��f���8�? f��B��0����ZM�c{j3XZ�!�����I�ݯ�a-7;[H䇛j"�1��:n��7I�/X�&�{շ�h �hT��!nT+aIJp)�(nӫ�g@qVP(dz�G�O��a7y2�����p�g�Tx�ո$8��g�ʗ�EZ�O�W�����w� d���sQˋH���&_u�c!�K䐷@M�j�=i�ǚ2��U�d]�0�\l��M��K�T���X����Ie�lw��?�V<�t�^�:�>�:Mޥ!!�����3����C'9����wD��v�r��l���fϮ-�̓�n!�YĘ���A�M�����F�¬�˛�_� ȉ��0�	(N�x���Z��N�ͥ�flH���vcC0��h�7����$^	�)9$�8U��z���H�ĶAx�Z��}bƅBeI�Z�h�J�����0�b��eҡ�+a���[	���E3'���ɺ���G�#)[�t�#E��x֕b+��$1�~�Up^Zv:0�p�ڸwN����I~���!���^��:�A�6�z\Bhq���x�#����ؘ
!G��}ZvRPׇxN�e&�YFIќ$���G2�O=D{N�O�i5K$F>���ܽW�%�Py4��~d6����C����K�q��f4��Oe~�K��Iu��qb!�֢89�X9d-��vJ-�S�z�*����b[��0<�r+�y���+U!G\�MGs#�ם7`��{'��h�|�Ux�:���<,OE=%��kz��� {��|��t�����M��k���GB>�Ԕ�>��/L�>[�c�`�V�(iD.2�u`���ض\x��a�mP���뵤������
b��S�YTs՝���[pq!����z�7��g����R<
@��!��������U��J��0Yl�6��b�*Xj�5��"���tC�p�o���]������]	=�x��B�/U��V 	���û�*F��L���q�*�W��PP�A��q���$�kP���I;Z��z=K�e4~�����)���ۼ����v����[��wu���/��r�.���g2j=�cU*p* �
?.LD�$6��c�K%׻+���)�����Q����"'7:e�C:4Hs�H:�H�@���m�w��m0�E���.t��8��V?-� ��s;;�
T;�����JGY��p�_(�r<,�pa��C��M{3��^{��d��?6e�y.*-PX��ֈ������������}�K�(��}>�A�_B])~���>�hq���:�E��Y����@�V 
�q��,��0=�V#|o�i�Y�ܪ�|���������>{KL�,h�Q$��2+N�r��D��qk=S�Chr�P���̻�J�f�a�k��t��K��ſW�@����t�J4߰xyqS��Rk�]�b��<j 'nT26.�Qt��e6��Jk�ɨ��<������������`�tEV�ٲ��Y^='%J��F	# �A�q���4\�cxn �Ќ ��۽���Mv��,Z=E�$��W�Z�wLz(�d~����S嚭�;��|95>��Q���u�n"uf^����f�;W��r~�ݦ-�Ԣ[ �
��x�WS���b�0��ԗY���-_�V��|	L}�d�����Lo��N1�J���nq'�V�O���b�1��0?5����B�~(�>nǧ�Ȟ��x�/�|'�iW�����d�g�5�Z+6�5w�|��[b�0�b�+MFI��A������W_��
gD?��w�m�^̠���E�qɚ����|���1��s�����>��[2D��*
\�� +G	-�S�x�2tN��w�t��|ݙ'�q� �v���>���0��W�1/E$�C����U�)lr|���I{XET���)oO+3��\5�<�[D(p
�պF�I���� [sό��¤)	e�v��&���q}Kb�&�CU�y��Ʌ��q�%$�]�h*9�{WၨN��(��s�/�d��i���P&�7����P���1hD�Z�֌�$�1H'�A�~�tbX=X��
p�II@f觇ӆ��fޥ��/�s0�������}����o4�6�EsgVm�VG%��<��1����4b�-�πX]҂Ц0<Â�[�g-Ku�Nk�I����yM���%t�/-��=�+"|�H�k�V��D�3�`�KI�m7�ɷ���>իL��Z�jixRIc��D�[#�ߎw�U*�qW֖\�>"�F�6�ٳ|���l(�H�����i�|*t�Ř<4#;	I4��*F�N�ϩ���ڸ�	��k&O(,����TO���#q���N[DA���v�%&�N.P'��>~IF���I4��]~N�%LyP*��J���%ͬ�eL�x�RF3��:�᫭��:&�v���~���͞���q��.�o� �+�53��v�v>N�j��>M��2�=�&h� ��N���[��a�ʦ.�82�P?}8���^����l&=� �7v�I���6�EK���4@j�tl�����NQ;��+�zLmU�����gI��h��|f�mɎ�+E50!���,FD�H7S���� ����c3D0UҤB�D`G��U�_�����#[�����܆��,yG�1׹��dP�W��Z�|� u�A��"�T�ˆ-� c�Rk�W�w{Kh��>�I��s"[Yg��m��;�f3Y�d�s�q�/�LY��lC���h��ʛ�~����s#"�5��n�c~����>\����D��F��5pQ��_�-[�q
�2)���{�V���v��R�b�i���O1dQA���Ҏ�@�z,ͼ\Y�X��=��Q#�³��[�ى���ب��a���4����Xw�{#�L)f|)��Al(���փ?�?�)j�}�⋣_�(F�2���x�,&ٍO�7�z�!�"b����y�w�3.:�ӎ�HĥB��8C�kI,7��M���;l�"�1j��2�X�Ý��+��pR{
��e
iP�N��Y���a�|z���k���+���Q`8�Ap�q
�U#�x(v������vϿ�9t�T�.%���	�Xu��D#̹D�a�bke4�K_R�cP�G�{�''�N?u��顤k>9hr�ꞷN�������ڍݑ�������"��x��*��߀^���*H��I9f��"��XD_I$6���O�O�n�A8����]������Xk�>o��A�t24% ��
9�TQvZ�8葏7��m��#*���H�&s�,B���sY}t�I�k9�j$�~�ճ߄�¯,=�6�Ap��8���>���ځG�Ax1UG�Gdr�IBp�y������"�9}r�|�Y��S�uJ`���DWRz^���]fy>��Õ���׊0��<�n��0���-	;Y��/��F�p"B�Z�s)�8Pⅆ�oę�I �OҌ�`[����m$I��D�
��E���OukI����u`ڐ*�(���}�;����[d�]�w�C�.o")�6�aNc'h����bLƜ�����g^�}�>��j�V?q"O=V�fD��;��m���ÌV[�E]�?_����>H�Y�m�ؕȿ%	"�v��mq�.�p��|)������vjJ���l�<q^;�|��P�N���G���/n#�M%#6�g�N�� �趓ť��ıi��R�&�Q� r�uН�9�$��Z��Ś�8誄�G��%�D�Ž|��wo<$H��
�T�������]���k��C�<�ŋ4��e�h�$��������_'�`�J
\n�{z=;���_����}q֞h�;�Ol?.�p�j.NL�jl)���95J!;�	G�?d�{����%_$��DY���'��:��D��Gl`�gU������$L�����v�xb���,ł�"#Di�Y
���#����L-Zd�4d�S!�&ϺV�s"H�#�J:����=s�:���X_b�n|!��w[v@}�6SвvC��ph�&N8�,��8���)M�x�#*+��'��^�`��1��2q��8l�u}�D��F؉���r����䵲�L��z����ɂp����k�����5l���R��A�\�#����	:-���ǘ���Q�ٛk)Av��%Dl?B�[ȹS+C�����S�:|l�i��D�?n
Ee�f����|��S�y:�ls@��('��aN��Z;��_�/w��!��K� G�I��]t�2�m�zE5R�^�<
Tq���:�ݏ�&e��gb[�iϒ�h�p9��-�2ü$����`nO&<�+�ɇ�� [N�l�ں�"�����8�@C�Tǣ����h&� ɪ�Y�������S��n�%��!Y*k}����r��'.��D�4ɨ���I)j�ϴ���s�B&*�j���I�1���/�9��-v��]�[���Gܫr"�W��gt��޸Wpɒ�#"@�hN�*%?:��Ib=��pC������tO{y�-��5{�U��#>8(F6>���V-C=�L3tSX i̸�ol�q�pm[EҜJ&��8'�j���6��уL���S� ��V͉�SG�5����z�
ȶ��v���,�1��_�3o�w�C7�jыl��N'�#��-����O�K����\�8��p@WE;"�򴆠���9k���>�]���L�vo\�a���t`���'��I�t�F�Ҧguq#--aƛG�xe�Y��{k.��(<j5�7`b/��)�����v�u���o�1Np	�Xf8�Oȵ91�QH)Vy����y��c�c��R�;��V�[�;�=r���K.ܵG�G��a�N�O�<4דs��@|^0�)��C�f��J��Es������cb�fӠb���%���X�J�ą���q��@����Մ5wc�P�v:n�����s���
a�����i۴k�m0��B�Y���t̫��ضߧAE.s�y���Q5�_&A��8zU����n�@���[6��G���4��E���7nU�J�� � ���)��Zhac-�]�8�?S��Z#t>p���)��[�Z88M�8%>TH�ysrVරb����)����c,��,��F�ݔ���GmwC3.���K�����ʗ|��d���~8���Y%߯�AM��N]	��7ݨiɱ����͕������LZ���IЌ�W��?��n&P���f�D���nQM� �6�[��#�!N�m'�(GI�S�O���"=�Ό\J�/��ZK?�?*������y�fy��& ��ᙼR-�D�Ơ8��XHڗ�k�0���#C ���t�T�kiq�#�������f�K����h>Ke+�[Ek͉C�h�9#���CVٿ�ǖB��N�H�f"��,�[{���Bh�S���(A�Q#i[��P�V}i_F���"9��%���ǿ�&����'�0������REY!&]��L�?�!�S9$,+��,��;����hѽ� ����-�w�"ۓ��"��8����,N�W炇ѐ�a,"�������/�B聆n���� &��1���?pH�`�z�G�̕�w�w��<�̰#�z�������k�F�Foj��͜�ey����sB;��=��Sm��������� �*ԔW�_�lyX��3P��:c����a8Yˬ�}�<aV	x�8�
�jZ.u�������ڑuCV�41��Q��+�W�f���)[�	��1L,܎�����k��iV��v��q��!(��)���N�{o�ی_Z��f�(�げ����8^����af�K�g�;�	��R2R;�!��J�Y�?`΋��-0����d�5�������}z���.�i���'�����&�S4V�S4M�kY*�ʒ
�
�a?����s =.Y��^�����>eST�	��Idmۺ��ݟ����r+�_T�Z|mR��Fz!*�$M���%�x�&�M�*�o��66�}+J<��-譴�A�0��X����)E�`[���[�� ��_�k�7��E�xo��m�JaWXjgF��y9���ь��:e,�a;Œ©7�[�����K!�?m�0�ȑ��?⟅?X�ΥJ�۟iʴc�Q��ac!�LJ�� �r؝]jC^[������&��E���<�c���{Ys�����Kǯ�Źj�gf�J�����^�5�F�1&W m
r��Axyxgv@W�yQ��^�|�WVU/:k�IUG�	�ӌ>��[�4����Z�e3��eq��;2��iH�7*b����;���u�_�c��Ʊx~�[k��"�oE��`,O�`�� �� ���F�aá���f��> ���Y�B�x�"�в��@MrEae���_��ؼ�����\� �N�Қ
A�qZ����M�7������%�Շioep�"n���r.�֗�g	�M�2U���c��g`c�=��G��߭*�Io�P�_��c�����M���K����a�z���84�o���(=�,����m�T�ғ%�[T�1LpNVWk�7��=���y|ۡ3�X�7�j�`n'�0$.3
Up�ؠ׷ EI�Y���� =�H�[ >X��i K�y)7�sc�4jB���\��?}�M3Эo�j�^������T�0�[�3�Y2���9B3����&�ukʅ��wG,'��z�G�T�V�;���ģ� �(ۜ�; 4��Sr�r����=��D�~ڍ�ۛ�8����WV���┧�?,��9���^pH�p&����
sjFx/REo�U��>��I�o5��='�	΂d_ϝ��j�!Y�!0�C��`f�	�~��,���,�	��������z�,�	%=�`�U����.X~H�.ܘ����<���r8䑟�=�O	ۣ_��w3K?P��%�z�+�ѱ���Wo�ΎO��d�6"?xv���,HdC��>vca�{ y�5_����E+�!�s�Ĩ����u�W�41/�rbV�`�U�_,�M�"fn�$˄���3}���HZ�O�e(L���HC��5I8�����k��F�Q���x. ������i��゗@=��/��>}l�`��[˄�`�0���^�`��'<@���e�N���xӘyw������(�>�u�a�X0�ʱ�#YQ�|e�^�?�ќ��
]
����)6v� 6�V
1q��z����Ėކ�T�d���+��k���W8	��I�52Qv�͟d�7��`<�w	G� �)�,]z��@��tJ\���B{��P�|�l�{OѦn�l&z;�^O��]�+��"е-�U����)8y��	�ק[R���D�!�S�->��@?D�ڰ�b����Oe([��8�$��7��3��r�_�m�FAi��E��0r0C�W�
X�݂�3h� '��؋�}��4F��%�]��Ɓ1+�a��s��&?�圊�t3�5��K�I���T~(���3I?a�\g�<b�ix�����pj�,�|_1��J7$j}�4��>��D�����[G6R����MN��.{�+; 0g`Քa�|�3R�Z�p���C݋W�jg�t:zbі_��eЎKT�^&��	4��b;��	��C��5�}�]z�_x� :^��[�*�=���9�J^�*(u@�@�f2%}�A�Z|���B��;G�j��YdV˰q��9G ���m����U����B"Q�V_R�e��A��=^�ނ��\��Z���]�˛�꣪$v���^jŘ$O��4�GxDiF�n�2���*���v�U� ZP��/����g�kKuX����V��x����x3.� �(Q����ob:Ĉ��޾���뒋{��&���q+�<�u��ם�b�s�K���hh|�$~���&��NA�B��h%�g�����'_�s�%�)�����(L�7�=���?X��'��o�Y��i/�i�h/<��AP����G[����R��?@��E�2~x�'NTк�'G�c��z'��2���˩�]k���?QgI����w���S�
�nb� �� �. %⍢�s�u!��_#ɗIml:ս���A3�<7�»4�?����"���B-����8<������e>�}��p���x~j.���KS�c^�� C��E�:N8�dj��R+�F�*�tԖ����?I:&�W'�6�IyZӰ.D�PC~��p�-�˦������s��ԕ#Ir�9\����'XR�O����i��� q�&4�>63p�h����Q�,�f����A�
��g3�d�K��fD]�n����m0:���s����_%�ݡ2Q!��E`���.r)`n����=:P�)��y���R���6�e�0��a�H��ļ�{�CE�M�`F���� ʋj%@���Lx�=�0[P��u��{����ogLIԟѫt�@OK��40�>���is*oo��lV��*�»���]���]�'P�Z$�:C�Jao�����b�1Ŵ"���x:k_HDM�P��YB��<�-������f&%�0��X��� �����P�4��te�9$PP�L��"mUH+�������p���B}��>\ܻ�lm��tևL�l���F�����-6��<�+��n�iX.E'�f�ݾ���ܓ��-%�yS��	�lH	,l���w���w�X�+���Œ����O��))�3K]����J2���5��N��1h��m$�{�?�)��2��eC�3��Y�QV�gɑU�R���9��3�ZM��E�����mN�c�+�9�2�ZMu�Tyk��䣋+yІ���o�؉�2��c�tKQ�S��_Ku,�����+R˦J~ʩ^̌<��3g��(�*�%-ϰ��,m����P3y��������1����x����ʮ9�@����9A�,1�'�l�;)C���ٲ��h����O-��$�����e��T��hp ���a�Ф�4e���5��TQ�H?n���T���-8!�W�%,�����&�c�6��DdA\�%��9'p(7��A�8�����6��ͥ�7($�]t=M�6�6�1��~;�C'IX�$D?�#��y1�x�V�)ͭ�5K����a�?���P6<�p�x�PD���5 �S;zk��j�
K�7���J������9}�5wC���?,x�u�1�a���9���c����Hd��W{8�$\�������_�,�X=�ػ���ӿܖ/�m	8W���Ubh�s�vnNnm�� ���f	o�� �}����+�
D����U8UF��*޷�Q9�ϓ����U��Pj���S�)�}*C���j*ט�V�M�ʝ�|���S@�)fG
�]��AȨ,B��&J���x^���}�1��ؒ# =< �E� �-�P������	Þ6u�]���:�a)��!���������/:}�~�^���X.��ϗ���nk
�׻�GX1A�����*-W��x�HS_w[JӀ!�gb����0�/����C����_��c���'�+��w}�Гi����l�*�8b��N�b+VX��^����L?c�gS��E�XP��=>I/>�8��r��}�KVL��^����?�j4<v���]�9 �xHzܠ8{����
ΐ�8�&��B.N�j�a��aJ������I�r���@� E��*>����3oZ��Ddb�Hj��Ɏ��7<�����-V��r�4��@� 	�� ������7�d�����[�S~˔�x`��;�0�����:�HQ��1tdc|�����ݴA2���ӛl:)eK�)��ND�T��t�سvY0�N��=��l��M�XA�̆�jm^4����\�ʞ7H�'�(7u�R^A���	��^����B����'uȰѝ�2NŚ&���`��a��qH��ԎD��wÉ�p�UكNQ5�RF;֍�BZ��#`ml[�Y~7(�V�Zf��ں���~�نF���Iߎ���)gLx��K�|B�k_��GhM���_O��P�o��#��Rc��q��:�L2�'|4$�����E������'�|Y���u���1}�\��H���	�Y�����+%Wcs���*]���!��3ˢ��eeZ�q�ݐ������2j���lp�n,���+��V�E3+.������HW�ôA�-��� �D2�x�,�7�|�;�]_�|��Ģ�2�2�h0_FUo~�j�t�I�Ͽ~���9C�Қ�2��u�C��y�*[Ϳ*�_5���<&�h�9&M�@�͘���CF`yn����<if&�D�yBO�y�<��`-b�mL\�?�S$"�β��K�h�F;0ТC�1�%U��1�d�%�|�C"����J�jM�%�Z0h��6r�/B����\"�����ߊ�z�E�Մ���� �)�p+k9$��P��ȑ�X��i`iB�Ĥ��R�n#�+?����@e7;�:�DuFs�#AtF��	5X���0mĭ4��L��)}Ȅ��$8��an�Q�¢Af���Q^�.$q+@�\�'~;�o�!���P_�R��;en"�.|�o���<?K���@,ݑ�1ra�ҩ�x�WPt�},)L���9��I;Wm{�V�����P�@���"�kN��/H)|~�XF\��hj�z��g ����'�g�ĒnR�Ç����]O|����P7��x��	�J�O�e?�����5�#~�9�G����A�NS;���٦�i���j�(y6�v	�αޝQ�M
a��-�,AT�'1tS܋����_3-�jÖ
R$N�����]�"n� �~������.�bpR�a��2��e�y��v�#����̿�Nj,S�>��i����K�ns��pcV<�74۽�����Ǡ!�KTb@���G}�F�W�ӮC�PG����*p��[�&a?l��#�(�=y϶	� ��xɷ�_��VN��8m�v%�$��1�=��E���ړ3�E������WZC5[�k�����*vʕ}�QԬ�yz�P>���6~�䐏�E%�Ú���`�V����),/��&���t%�閔Ѧ��Kϲ"�R����=:q�N'.S&���j�i�y���pJd��h:�O�Q�ϧwg�XG�4$eD�@�<�!0B�������N<��l9,s�z�x�2
$�����ɧ����cS�Ǖ�KW���>Y?�NeWi1�~������v'R��n�R��bϔt'"��0�~"~�yK�tCw��{�%��g{�ւ�۲wԸ��_4i1�l��潪�7�`�2��'%�F#��!�����F�~;�hu�����C��L���m�Q7J�E'\�꨻�1éx����IL�&\�K���)ON�|?� �����%%�+��_����k'D������)kc2�8WԶ�l�ᔊ
Ji|��Y�	�-�?7����n[��6g%0^ּ[��P���-SmEc��������8��/����Tȕ�f����hZ�������Б`+l}W�A�`��}���^����Am�"Q��K�?�&tHp����PN!�	��+�)3/�n�<+t'T}��ib6�Չʣ��*SsN������ɤ�!��}���m�������:�3��d,�� S�_5
pj4�F6�c�a˖��rZ!	��I��-_�o��g���'�Y�2������]&�ʛk1f���zbKxv�T	p�2C�B�㯑yS�d��:�4`�j�Y(��Zt��V�b����n�?|����(�1Je��l�9[��m\/�\�5*^�iNr�/6� �
I]�9 4�P@/�ͬ���-���-8u�$V�o纊� �l7+��
��3زĸH
������l������k���S`֨;()L�[��^��8�HY�UT�IqF�`_�b��>�|�w_��0�CŻ�dJ�4�oP�ry!L��{+����%��p	�L��!	���AB��I�G_�Đĥ�kX}Z��<��,������M��s�,��m���.\��AK� S����G���e��B"$:+W�$:����T8�.�[й�ji�$A��.��|�Յ1�O�� z����4��5A3ϝ �p��}��h%ܓ�)R�M�fmS��M]DǇM1N����D_r�Ó����}XVg�ꍼ招��#7W{�6�e�f�5�IjX�֑W��� ;�S<�I0����o�Λ��I�8��gًw�B+�;��l�1PnY`�&o��L(kA��v�q���\�e��W���,��dț�c���Y�ie�ǚg�K� #x֢c�Ԥ�|֍�T�����ޢ������Ϝ�wɵ��8`Xu��D'P)�n�^��tt�&ʹV	�������c�ҥ"喍��_ T��X���Z��3ir荱yB�3�hld퓌Ug�R��_yl�5z�(`��/6���r����c��T�g"��SՕ�+���n�n�&���~��#���պ)܃�Мu6���;t&��iB�_٣��#|�_
K3'���kb�Zi�*��7GE����%i��/c��6�����e�,������6�+�i��~,��n�u�7��AP��Pn�g�*ugx���C-�JA�U���D�k�#R����/nKDۯ�S�)�%PW�;���݄�> � (!~,��X-��1,�i@+�di�VCĹ��g����UՓ�u���a��|ږ��S���i5,�i��H�X	O;n�J������C!�j�.[�;��m� �r��2�E���-"8�Մ��]�����ޒ����o
��E(�;�ߊ7v��M<}�k&�7�$�V�u���Y5��Wq5o��o�nnv�b�wK��.#��S#�{9#In��0��~��c_��X� �hYm�W��+|e��B��fsMc����N�Mf5l�g�t�W��)32��z9��[�*�<L����b.?3�pWk�y�)kk��|=4?�&eQ�=>�� ��7TD\X� �1+9����b��O�Ř*xCx��#%-9�ox�Bi����������3�����`c�>�<?���Ƈ�("��P,�;�zp���CF:�*�Ň�fD�����r
�}{^a��ۆ>�pO�fY�jme��x�_f[>�����w)��*��m`r���	&�^���p�C6<^p"��]�P�#a	|�D?�]�vd���9r����7��}R#4g�k����=�!wd���X!D��{5�SQ�%Io�w������)�.Ӧ�o)_\�3��R8I������U;��a�p=mL5�%j��Q�p������eg����1�����Gc��-$U�:��VZsb���sU�q��H�h]|Ts�Y�M�����o� `�Ȇt��>���]���E-�ށ�l�f����SS��R���(��%�$[����<_��U ��k����"_�����a%M���A�Z���ȕ��`�/tiN��6Kg"�q帺2u�!Uػ�Ֆ1�$��cv�\-&5[�t��Zx�!���ڼ7k"�.�=5���|��� �I�͚��T�U����v/������ |2�\W���j7�'|�
�ܘQ.�dY&jVDP3�k$���`���j�A�lf��($��~�g��u�mЖܲ�mq,��$?���+���q���7��@�ͻ��0:�'Ng�$���v�Q�v<��^d;�W��9 G'�:@����r�Ren�N��F@\W��i�K���� 70���~�0��ֹ`SB�|�g���'�VA���2l ��H��E_��6�Q�|�k%�����l�D����t�;e��P�����������E:�aJ^M��%]�m�Eן�ãx���ܨ��>5�"1'ŐMG���qG���L���m�e�C^ʀ��tk�Z�A��(�+��j���T��H��摖��!Rt���(�D^�'��8}��r�4Q9ǻ%�CU���<%<�3�.G`���_�:`��f��V��i������Xߝ�������GSm�i���]״>pL���}_٘m�#����(�<+D�홏G���r��CY�B���� Rg�3,U$Nm&;	���콚N��q/�Iٙ�Ʒa�4wp��{���^μ# �)f��j٫ޙ�3�T�[P@ŧ[ݻ ~�Z�J(S�9�0D��YK`_��pl}rI��x4-͛%� ��%�&j�ي��;e.A��yKna6�i������I�7�U�(�Pݒ�#{{H�LcO)K6fG��E@{E�i�w|��n���`|aIQMbͩ�|0��!P����Jc�k������� ��[��2
��W�CpD�	�o^��N��N��W��.Ǭ�)�[�� xpG(n��L��/$�
Кu�ё,��e�D#r�����G��o1vP��J.�%t"yn�ܽ˴n�8��r��9�AL��}er�ܓ���O�S�u.�
,.�<:��`�\��t���,�1Fv�u����I��,�- y:0�Ne�@e�m:�}������s�Ѵ��z ���rT�R�+g�-�-�z�d�
A�]n:�t'sVj*��������ܦ���F�S�^���.�5�l���z�g��/�3�N�]8��Jp?��"��q�����+��Y&~�m�g]�7,�ҩ���Ȥ�/&�dyar&�O��G���1w"�����r栗����kf�ʟ�-fV�B��T$��ߓ�7���P���	��	 |���$��@�/�uӳ}��<�_+���j��פ��������Ռ�Ʉ틘�墷�n��y$_�_���#����I����y.�N&#�2��Vt"
3�������Se����(�<�{>�����\!v�~Je�����TD,�..��[@�׹I;
��:��v8-����_�%�e�ŲmA��+g��a�"�F�e�Y|}�񸳿o���R~E��!i�j�\�hc�A�`�[҂bQ�i�-��Z�!)��j��)��<�u��`��5%F�g���rk�V���ӟ�硐7��^KU�P��{D_S�6�'^/��%D(4�0e@��%������Tu\�b� �j'�wu:nV^� v�q�������
��=(�M�{@DB����vM��r	:��Fw���^=�V 
`@���q�4�((N�G-2C��u4V_a����W�Y .dC�cA&<6���
*mC%8?q܁�LJ�Y;E�%��W*�y7��!W�Y��i�Oh��� ���<�%�I��# �oI՟l�"� ��R6��?��批"XD��!�,[��B���Ub���x�������ʮ��Zw4�)ɀ��C�!��g�k����X�R6���&b�?n`�fW6��#������������e5��C�?�fD��e�tM��Y�X�?�kōl� ěJ�^ϟ� U��UV�O�M|�d9���D���	�d9��IE������UYgQf��l�%�����dq�f}�����%K�Dsn�SZv���y�K
rw�~fM���!}K�z;���Y϶L�ޱ�y�+�잵p��	�~���j$5�vIo?/Kq��2�D?�w!�6��m��x�1\.T���<��G4��$���a��S6��#�9[�L1�c_�:��p��V�-��F�ORݎ�کN:k�Ck~�������ͩb8�^ ��Ǻ�yP`�՞a[d�n���l��۟��1U�~��̖aga�|Ã�n�Li<�B�T�C~�6e���	�M\`��=rr��W
�&�V2A})����bQ&�C���\��qE�8�cj2�``� yqޓ#�����T���үp��~�O�Ÿ6��n�T�n�0�^Q��̐&t �s�'���x�Q�".>,��jMH����
ޱ�X�:�@��>��ӛP���	��/��b6�h�΂^�j�7��t����f��#Pf� =�V��tc�����-1[���0��2�j��y��g��VMe`.E4�t'�b�h8D����Xq46h�1� ��c$#��jsП���qW� �Z�NKZ��$�U����꾇w��L�u��] DtZk�VI�7R�P%��}�?ٙ�T�Q�������7��i�+�#ZM�(A+��Y��1��}�&VX=�6d�ur�)~�O�+h� w^��M8����j�7��R�:��uJa���j�6U��bP�k��$�>�Ȩb;;��ʼ׾ƾ�V����7b)`/�AQ�0kC��H�6F��@ƥ�O�,�&�ʪ!��(�\�bB�h��)8\�<�%e�᫝ܿ�f�IƖu�	th�m#�Ǖ�֖�s٠��	��1�qԜ������4�B�t�K7��7�U"l�c�Ҙ��<#�ޜ�݇��<CL�A��J��U\��ࠣkaɶ����Q6{�1l���]l*bmE$������G�0-�-��Y�N{i��N�CO|6NXQ��CoXr<@��V��B��x2�+'r�g���޷5p�G����6��͘ϯNRr��nu���.o�B���k��0+V8���-ԓ+�֡G,��a�x[4�L'��_ﾥb��e%��)j����7�4�y� o��������u�BK�؉���Z���aj����R������k�u�Q�.�������ҥ�m��{=�~��[�w\��ٮ�%6����N8��l��Ъ"5���X$hQb,��~4�ڀ:m�j��N��c���BH��m%ȐU7�=��&�FdC_�Z�o�X|�C��A[ń�{�?�"(����Eq�6��n�x��?��AJ���u�ڤj��~�T�[%=:�t
-
�����o
����uW�H��ꎠxK�����[��s��O��Ǜ���.AJk��g'�d�Ƭ�U)��u�lb(�)���W�n�a�F��ʡ`�Kͥ9~v����]��k�Y[��V��O����?�V������&�{�5��g�::�fja+�0
^�nD�=�h����g����g�����͹«��jE�\tB� z�`��;D3�ʨw_Z����5e#�:8�����(��E;�hq,]�+'9�S�� ٰ+��*|�D%�U���f'!���x_"w~�AB�mwdb�)_(6�H�0�-��%#8��e���4���S��d�4�M������9(_h���&=G=	dm�%��|�)�t*$_��8�="M����h��2ʉ��:ə���$����\(Y�����y�55����
�������`\`l:�u�2Ry�BMq��n���!�'�׶��\�ZKwl#� ������ ��4���.ė�{1�d�lb�d-��Rd�n��YۄoE+@�S~ˉ��R��n�*-�O�*}z>�����K��4mF�IF�H�G.P:�5���K�S���@�0Jޔ+e�ZP{�VT�"��!�cS'�P�xF��~�YG�^
�ߒ4�F�X;[B[���]b���x����s�aC%������<�ҭ���v�y��|��J��i�;w��}��G�'�7�y�L���5Mا�|š7��L�>�-��3_�����)[��D�8	�i)�&�v�� k��z����'Mt�oǡ��߰��#UJ{��{4�˨��N�\Z�ݖhw�%8���2��^�E幂�#ڮ�z��Fu�
h؛��-��9;t��˶m�������%�^�L�#�9�>�K�*�����h�����<h&�d��~��\W�8�+D���K��{H���'�E2������� Q1�Bb���Ҷ�$r���+�[[Z?m�T����	�b?d8����N^�^A�%Ӑ�}!��r1U���q'C���
C�E�ϲKEv���3��|����	�܃�2˴� A��1�	e2��)] ���W��/�5%��_Q��7�
�t����ωi��%I�W��8~6�I1�]�b�<:����>y`�ہ�#g%�T�����h��7�g,��ӚR��F��#F�5U쉞����I����B�.:T,(N�!)�������� ��2��*�����p��`��ɿ|�m�L��TJ�+�G�DG��?�Ղ�hR8���Ȑ�h3��̜�/W\p.�w7H"��f�t�v�Q����͆pul��O�?��l�]�N��iE�4��/0�`CWj��:*T����&��=��U������ ���bUgGT�ؿ1�,9#�编�@|QN���*X-:��@��әp�"���i�4|��*pͨ?�'� K�I�����!��J_�����Z�\؋P]vg��k�q���\�J)��k��oCܞ�3l���t�t�rI&����6�\�KX-R����2����:������%D�}�j|����5t��6S���^�*%���1�%����\
"z���q6|��CP�}���/9�NO��e���������TL�J%�T�t����):���<��S���'b�g'�h1(9�� �e�M?Fo�'0�
��PA�e��r:�L^":���l��*�;2������ş�s�K��`�e�����J�OJZO���,P�Q��.e� ��C��.��ʬ<eg|���=�`��A>�+;ႣA]�餓���� u�3�%�9�>�xl��6��V�.$��3 ��!\�^�o�-�1�U�#�l�UL�D�	H%��'�3$B_)U�� ��iv�kbU�9Y�!��D�o��e���d���� w�e�����ˤ�?��@��2��A"L��s�h_��N�q�$X��,� g-�6�d�v��f�����2Z��Nʄ
��o.��@y}N��F�Ȱ�ze��f]ٛ��M}�Oj[k�5�U*��7�	�Z�ߠ���,�Q#d���'��� %��@D�M�����j78Y7*�Mb���n#����n�	���G��^�r��vC͖�o7B���������kSl��(��np�%J������67��	�[S)/�9�˨~�D���5���A:��; �~ o��{�c�oQ�U�&�ǋp������(b�`*���`���|��YH~��򄵇S�L�t�uK�GM�h����0�B	O��Y�}M�Y���rM�JiG`�؀ �"JZ�j�346�V�%�R��i����9z���\�ƾ�%�b_�$B%?|�qT�!��M�{M{K��av�+�#�\
�߆YBi��CDM�������|}��:���sk���W�!Um�w-
�Z�o��t>$b_�`2"uKc4�U!��1�t���LJ�0�o����WԷ�6��x��6evK��f����j�u\����D�MD����H?���0�����7ܙ�LM��9!��_�޴8�2q�� �=����U�G墂�$�{U��%��Y��Гg}�O������|�l��X&{��G�}�� �J�k��om�s��w���0�'�B�)l�wI/���E�j�׏RH�ޫ�"�?�������S��䎭�ӓ�uW�#:��T~X��b.������+b���N�)�Y�	B����i��3�*��t���6�1�q��w���A#��{��	�]C.P$�2FWLr�u�����.�����ں�s�<��h������֢g�yqĕ׏U �RF����Bp�R�-%����*�>���MaG�؅.���HY}�kd�[�������ٰ��]�!ﱳ��m�a�H�r��Ϲ�B�nMZ7X��;I^H=��)^���>�BKҹ%�.�ݏ��q�?ϪK5t�9���$'�0:�<C!��
��80�����'P�<i|��ެ�~�w^�f�A�E%B
�!�Y��IV��$�r�	��g�������)�Zw_�]L�ˍ£0t����jJ�n�����P��_Yɦ�W�Z��d �.���=i.�?��ܐ�D�'�� �-cnXνI�AH2S[V�vo��1f��wӱ1�5 �y�������p�6G�l�F�&B�@h	�R���C��ț��������YO�N�����5{�:�#��9��B ����9Y�m���a$iJ�UY?�u�o�'���[�hш�4��j�P� ����=�[����3����c9�@vٞ7�w ���u�;n���s�e����:<�/��j#V��O�(�����ל6���[���|CL�����m|�4���!�V�(��rݷ2 ͟_(ͥk$�Ŗj�9�񩪒ҔR{m`V��7�0]����	l>~�:�u��w��+Fɴ��a��jM���V�ۈ�<�h&�X�I�(~̍)+�q�/.y�\)�:�?��Պ��mhQ��YY7�� ��&*p��%  ����Īƚk1g��� ��+��X���e�wGY�)�b�!*�����э{|QԲ:+j�]I,nP����vP�*���ߖ8PA����)������K��q�J���d���%�z]�����������e5��n3~	ށ�ܭ@�X�X$��z<؆0��o��I��7jҐQ��&<�������z�"!�E��Y�LϡO"��9M����_�	B�i��ɡ�+o����u_�x�/S�WF0�
��W&+�H�ȮvIh />��c~�-(��	��G3�"r����.�)�����-�"[����ݏ��^/�s�݈wsR�ؿ�G`3��8�S�~?��ȃ7�Z"�t)3X��~F���o/%���]KK?'��ޙсA)Y*;��I��1���v��,�1}Ȃ��?WԄ����������|��!;���N�y�I\cGc;�<U�1@����~1�}w�����	�o�<.�Z�j�����Y� Q(NƜ]2�g�!q����>�A^3����2AM�D�a\���s�R\�?0vJ��l.k���t]6'�C$Q�|�sA��r��Te��X��V��4���ή�*g��L��ÿ#$��S쀒V�?��g�;�m�f�2vYY��,� w�_��PA>l@�7�SȆm�Y�8y��:7�%�-�"8>!��DU M�MQ!!^���D�^��W���0�O��ω�J�"\֌�)vS��s<�yG5�<]�qL����Q���a�e����ӟ�n
2[kI��8OL4�^?a����
�6���_�ȼ�]/��v1D�]H�@�yv���G�s7O&s��A*��S@BPT������͋��cུ��N||$�e2>[�nZ���z��H/Fr���3�̧:߻y��1V6���bHB���Ǵ���4�Z4@�{�F�ܗ��DeM����6=/�h{(+�xW�vj�m�h�R��/�������Og��L��B-�zc���r�t��M�M���Ƕ�k��/�6���L��-8����g`Sm��[<1,�=AN�S��u�l�.yVL��6�j��a�JgŹ��v�|"�ً���C`Qps1p����,��Ȫ�L)*�����>�٤0���+<.��M{����G����s��6�Nf����@�`�m�=#��C,'�O��R\�_s�̟��j�}����Wz�|�H����,l�?Ǥ�X���if���0·�7�=�0�������|'��S���o�=v�*+~Q�,�E�u��VL2y������hN�Nj��Y|�@,Jn�%c��E5a9�p:o��M8d׾GQCi,ub�!J�/��'F�w^Le����|��M�a��f`�X�����#M[r��O�N,Ay��K(��$�L�7b��($� u���� ��~��X��ǽÅD
mƼӀ:�������1��
�zcݓ/(�4��ZpQ�\��X�E��Cr�B#���p��?���Y�u5	��` >�{(����)s]����R����V)�&�_�D��9�M^�g�����	@�Lo�)DE�'>Q��D�h�fzX��P`��A�9K�%Zӑ_�C%��o�S�07.8�K�.�����J��g���.Ѽ��[[�����aD>���hR1���NK�R�ӏ�]ȚU�h��8\���/�z�b���,�~Ӕ�3�bx���<�lA�@�B�	Y^�e��6O�Q�%�|r��K+q���)$C���"z�?�U'}B'�ZG����CԹs|1���_����[��	��y?�����v��?Z����ͼhx.�R6&&ū4Bgɖ���?%��5r�[�=��qd݋~99��T�.��q�2D����Xt�dF�Y+��@&��җ��M߸u�Ub��+��̞O=���`n�s��Z?=b�pF6:�Jz��N�ښ'd*B�4T@/&�z����Z�Gh�=�zP+т��� G-X�o(D���CKj��e�65���=�eg�#��7�XxiS19��,,W�7d�:	�^�z�	��^�aT��8���W�q���z�X<fa��B�=Um��&	+�Y���\nL<�+	�@3E�&�S��`B������㟒�C]:����� 2�=YN���ul�`YJ�FQ�y���c�H���'����r?�MS��<NM�Z[���Z��|k�����Z:0��g[2Fj7�,�҉����0��]�<t����{�@��KpܸX���:���7�0���qA|hs�	���K\Il����̟7ѥ�5�+�m���ؠ��8Nj'�J��@t\���@�#�=�TQ�w�w�.�<<�x �'g~�������VR�x�~��2��s�K���6�����'��0���.ji��)cH�t�5�>�89�-��u�.9�����p���L��F�C��1�0{]���Y��u�ͱ�y��V�ծ��lĲH^\b��tf��Ũje#�"K7�~�6�p���$�������@U>�Ϊݚ�� iC�qO��q����x�>�2@�P��#��l�8�@�em @���|������$γ�d�6e�ѣ���c��4�H���r��-GC��)���ɉ�ʫs��(?g�Bb�ph��F��(��=5H��6m��.j�րOs>2��*���k��++�VR^�!�깒���/vs�
�Z7-+Hjyᠬtp�2:ZK��p-œ5���>���پ�2��Թy�I���)v�N��^��(��t̟��fT���1��9��#ߗ��	L�«crD���N^��7��;@�t]����N��_�Z�v�)�ۄ)`�8�� UwB�>��j��x�~s���KU��5nO�-t*��]*]�w��>�5y�Yi�)�I�T����l��H��E
0MPҭ�;I:��9:�%tc��$�wRp(n���c��_L��I&���X��v�k�T� v�!�+�\�=����-O�5�^���=���v��>�={ihe,��JI�դ]��jC��;�-Xn���\�����ۿ��,{;-�i1��V�Ye�>��0d��h���j}�Y��Z��d�/;Ý����읍���C�O��U�9��C�X,Ym?��8H�ƕsR�"���ӵ�R8Y�y�6�w��!�	�#b��X$Ⱥ^��hc��~����H�!�_|�=�D�D��lL;M�%#U��XB�h�լ�t��7�� vHK�ݽ���%��4tձ_�� L"]�]�h���N����4��uS�f��F��h���1,����!�P�#��`%�@�G������ ��������ݶ�}ټ�@��F\F��C�X�� �9�v*YQ�?�w�c50�g�RtiEH_Y߄����a�*sK!��ՙ$dWV`ɭ���H}��}1�Uo�51lJ�H|df)��%�tr �WY:]�L����������1߹kH[o�A�x!t��I�C8w�w7��B�j*�{n�I� ���J�@�t�-�kD�S��<��B{�r�`�s�.H�Ec���ؽ��m�@����'10w7Z���u5
������q���wH�ڴ�2�lm�؏��\`�XnQ�4<O�֨�?�;���#[n�({��C�+vI�q�J��Ea��i݁��	g�N��!eW��2�,E��1u�P{�ߐ��Gx��J2��ݑ�}��T�L�A�fg�Q�}
��M�(��g0T��jt�Nųkr��)S%�b�l �J�!@�a�I,B������nu�o?s1�*�Cw���8v�U�����q[#��Aa���-ǿSAypJq�_��lDp�P�
�}4�gь&�y^c3y�?sxۊyb{��I�H�N"�%��e�����=�����k�6��<&VMz�,d��5p��@�+go���R1=��<�p�a��$����XR�ߍ��fA��Ӿ�n�#/�p�AG���F��o�zT*۽ޥ���W��B&Da��G���.=��A���|�=�3�p7y�L�J��vi���N��5��:'�Ju߾ˎZ���kD|�y�P��N����l0+�-_3�d��nN��"�ot�
��-� ���c
��W�_Q˽|��/�N�RdF��$3���~:򲭛����^�R�
Ǫ�\����7}xO��goZ�{o�$�?Ȑ�8���d
$�
;�D�s"T\���9��,9�e��_�t�]:�"��ͷ�nY��<�����@��QVc�{�G�z�T5�!��"8	��S�8ݭ������Ũ�+ݘu��ɓY�9W�b��*���xF��F�[
�����q+�1��цp�e���#7L��ޛ�|�F��XqI$�'�1#j����1�ްL,�A���|`��Ąt������'��h��X���I�q�[ �"-�v�������Mt�QE���,b�smf/��&P��9 ֐WxP�Ĉ��G �VD_-�]^
��n�rm����ƉӬ�'�,�V��↸�&�K��fTݘ>2^��KYL��x��Z������𡕕k:��_�k`���H�2�7����A&���:1���uVd;��9)6_�XFwt����}��4#�!HH��im#�B��+� �R�}W�;�J/�������,.��>n�P��8Xh8�F��GK�
.\yQrU��<���OD�Ҡ�V��0�o�(]�$r|2�Q5�f�T�b�b������g�xLڗo�f����2�Ǘ���z|�ux�V"��gV#�XDtS��̹��q�R����9��*�%D��ȕp+���w������ �(���g�#eE�@�O�m_'����R�t��N\=,CP� ���3�U�$�{�H18�o?WD�ط��w�/���SZ3�� �HT�&�!m@��z�;m+� ��F�E�^����\�}f9���5Th֙�ݎį�?BX�vP�Q��GP��Z|�=K����L��D$�J���tP���h��N)q�C_Rp�r�@p\{| �kn���eГ�0�sq'R{�x�S#�r���@��r��|1��KkYa��m:���r�e�g @S}|GFI�76E,�'����Wu/*RW+��G�|����b���c�L� q�0%I�2��VB^�3�&�9O?Q1|��.Ž�'�at�	�A�&��w$�E��h�Ml�������z4��#�L9�솵̶�z@(��m���sބ���W�4��j��%S���ˉ�T����t�u�vK�1�R��sX�V49�]��� 5F���h�..b"����X�`���zaW<���7$C���eEy��-�#.�ʄ�o;�u�M9o�]p���=���F��'�i��a�"~�������Fy0�7�κ |d��?�|��*G��Nt��a��{ �+r����Lr9��r���VM��p���2������}����k�; ��F��mNK�.5G�#�i2�^��ffo7I�N$M�+|�e�f�{�'E��. ~*S{���^\��ͷ��C��f9CL��RHv)7|�_���1c�&���vv�~����n�g�o�r�w�<��KW1� ��B!�9n���2/I��]Ӫ(%:Tڐ��w.��_>x��M��0�z���G��y�U�J6��ᅙ�L�h�l<�t�Qh�}��������Bu��w*0��H��|ϟ�v�D��7�䝩��c�,~v5��.�w�t���U��F�;M�(tUxI^d��|���$2��D��,l|��[�38�mm�1��]s�`�>f��&�l�����nF2Xe���5C:������g�sa�a#���z�|^����=��3~��P2���i�[��i.ash�3�fΦ�1�E����Q;�	�t��7"��0&.���p����*6s��;����J/��;���-e�=�}�⮷���	/��ѭ��8�E)�1�$�W���4��Y0�Yv��z�,@>���u�����-c{����:��}'����8�^P�������r�VW�^���5u.9���V19/iO}�jv
5]pj�"�n	 4�R(8]~���Y\��/f�������IW����z�Ԏ�Е{7�p7�fC��m��
��}3�&9V'�U�.bE��Ų؈�x�?�nh��/V���LӐ�/$�'�t����BU�^�����x��S��rbFK���r��������fA��A`�ceb��М�=FK���G���86��s�JA���eC� ^a�>R��7,E��������u��2h�eYt��VQ��#��f� �;�b�N\�h?daV�Ne˶&���ca5�`�~)� ˝.P��qB�'���ֿ��J�{��Ռ2$0x��s��~��Tl������E%V8��Hߤ������?�4{�-���K��ɰ����'��T�|�	��T�<��v�j�J������+l�b7D{��~�
'|4v8$o$?]3�Up�^,��c�vG���B�(">�Ź(&SW�i'�B�K�I���T�S��ܐ�	��|=ٱD�UN�S�g��N���0�G�K�B�qX����A��٪5�z�it��gC1��s
���n���:�%�xX;��>AH� �4Ü�*Q�m�y�TK��uT�0{it+�
�:51`����n��Ҙ��l �lt�T�h]�ex�X�p,�?�}Q5����f��Jڇz��/�=�YU���Y�A���:?� ���`��0���Ĝ�ϑǯ��ó-���9؋פ��K�f� �R���� �^`ʸ\��I��:~�A�h��	��>ܜl���EF��Ǯ�T*����&�ӏ�j0�鯲��(]V��E~jB�Bz������S;��0.�	Y!/� >Co�E"��]�!�E-.T%^^�m�Gv���E����q�����@�>ي����/�� �$��n,� ���ԝk^Ѽ��AϘ)��Ha6ݷ̻�N�{V��9�o/Ȉ��kpkͽ��+�~�֎�\SOEνi��B}���Øn�S�+�z�(����kdda��J��GOG�󰓯��z�����K�VASą^�P�g2ͫ���]�Z'�#A�[�'���.� � ߔ�pI�YmTL6_8w:Ө��G�3^:tǸ	B61 }��hT�}����xjI8O�A���)WGP`�����9�����~��0}+xLN3O���:�5i5�Ao<˵�9�nAʹ� �ǌ����}�zc�"�J�C���CcA�ð���+|�� ��-��FD��'C�l���M�Ҩ!ay>��Sʉ��/�&uEw!���ʤ.h��W����'TΉw�`�t���ރ%��N�{�nJ�⌔������t����JX6"��
�7�qD*�M6{�B��V%��c^���;)����Ţ<旨<���r i# [{��/���5��6�n�>#��<%��R!@�쳟OI�$��aNw�,��"��Z����Ӗ�'�?Ƈ"��pA�A�Or��b#l�2?,h�v';Th��_��?")��(�`
��6T�ȫ�[N����:�js�m����V'=I�*��> �vq!>`^2��'^f�8r�ۛ�#qf8Xʹ�_��PWXa3O�*�l�fD���@s�)�Ч+c�JD@�]��Ț��F	����Y�IFp91�:��(�>�h���A�[a�3s�O$�"̵?!�Jlp$\��i>a�]�L���)'����S��m�7�s*imY�Y�Z���[�Ai���y,����H�Z��_;���7AiؘRy69��r�����32�3�Σ�1� � ��M�Sw�A�T���C�Xâ@cOISqI����vI���w
��f�*�^���y�NL
���<m�4�|��J����SW6��Blc�cF���tf����pZcz�{�-�%!�@ ��=�w�ȉDϰ�i��_��?@js�'�@�qB�����+yː:y@X1�����3��|�ɍ�6L��I���b��L޼�@�у����X	<R��RF�}���MA�Ս��'�{D0-��ǎK����9�hɡo��#�P��.���ޙ��e;ZY����{p��+�K��i�q#^)�����l�J��̳��nvZ����v�ج�@��G�μ����9��G�H������+�j�����z88Q7�N�"��ow���%x-��@��X�*F:�zG�YB辣��^�G*t����kb�]�Z�55!�`y�)�at�x�]Hf6�T�_�u0�\�p&�*���&	䍃A��XOOu��w_W�m� J�&�[W@
�Z��]�C��J��s���0Vo�Z��GT�� ^��(�'����br�x��jЈYQ�^z䖸 x-����-Iqy�����ƨlH�GI޵�?��[>~]Y0�P{�M?�!?Fr������g;^&>ZBE� =�a��e��x��V �A����	B�Y����D@Q.�z
���ݦ��.�_������<����!���c�0����B?�`d�9uK�V����r��`��ɬ�ڼ�mQ��t˸t�c��m�yF�v87ć�-���K_��D��?<����7eo+�(�\�631�6���w��:'�t������O;��؇Ã�A�!\VQ�O�主h�Y���Gǂ�k�����Q�[XFD$�e@_���'b9���|�*�L^��h��o��3zo˖zǠ��^�e�|@N��J m��е$��L�o'��n�\�T՚���/��3V`����t�E�������'���W�\+s��1%�!��&<u%�y��^$����򥦎[��P��y0:쫸?���+q��w�$
��-%���쩺Gȍ(��v`�H�ԙԷ~����E]e5��d)�aۄ7;����iq��N���H=�S{C�f��rĬ��X/C�&.6=��=��U�Y&LI�I9�:ۆ[S�πˋ}�	y[�8�{k�8�u��̡R�HC�W�bw�!Xft3�;�GJ �m��6P?C��y�m���-ˬ�,b������dpP�%���W�9�4��k���*���Ʊ�`��u�EH�aE����#��P�����/���RW�6�wب��ۥ>�r�K�$�L�}5c����R��;�]��,��2s0���A�YG���jj�#�3��{����*�̻y%�0Bw��UF�DI<��n�zo��U�j�X>M5�^�TwG�r���h.��O^j�ԓ��h�`���&U���[Z!��V�H#�"/Q�����;�^���l�؈.|8�C��R �쵔�oD��?�/e�>*���v�.�fԛA�:�bker�$���g���s�V��oߙ�cx�R���ڃ7Y���i���Rʽ��V�)6Ih��ݢr���r���.�M��?F�z.��3ZTf�4�G�ِiu�q�O�ԎO��y�����#��i�.�#������Ыµ��T?�;�N�O��f;�|W-å@��:��s�s�}V{i|K]���A����p��;�:��[%�л�};g�b��n����j��?�),I��+up�D��˾��x62���E�oߩ+��B�2ҹђ���7sy9��
���D����vu��w#���Q�[S'�(\㯬����I�|jKB��^��a|�Ug�n�6��m�&�7"m�{�[���N�]�w���˃y�z�^YΊ�j��c��c�}�A�W���24`���x�`�bSԈ�"\�n��
&��\���j��e4e��K�Xmv����/�[
y�����h��#���G�w����
=4�w�%����Α_)�CB��0�YO�ꪕ�"�O*�+��ݘ����8�t~Ǡ�C�d���XpI2nCa�����N��(6���Ɲϒ(D� ��Bx�)d{� �؍���Ib��b!�ODvI�.���g�[�Eq�ad�N,\�Ȧ�JS7[�2��u�c��,c���Ѕ�C�y=-�����Gc�ko�6y��dH�k�ߓQ~i_!r�[��:�%��Z���_�
�

t`<3\�s㨓��c��b�KR�u=?�I�(��>�c6D�k��'��6I������Mo���{=��kv�G�cU/L�q�-YE�z%G���)Ǟd8d����m+�	1Bh1�:G�����<�*@=�JJ���Ps����dA	e�mKS�3:S�E�(�]1���^���׷�����!�>sp���:�:5��ERH��W���R_u�ze!�k�e�J�H���c'+�����G����r�;Ci��-�C΢����g<��TX;l���,j�Z�2$a*�)����%sl��񪅨%�ɬH��Q���q�0���Ÿ#�^Fէd��IB��߀J��Ka{z$���]�����F���AP.�q��l&6��?S���v4�n�{~�n�c���s˃@���J��K��'�hOA.�x�1p�f��PS�ʢ��}+��o�b�ML2��J�$K:5�m��:�K]`�l�����Y%�����_���b�+�T��Lc�=��f�G���1&lK8׸���t�>�o>�����L?�P :��zm!�FC��(X�!�f"��^�~U)���,��h�HQIԷB�?���V�i�X�eh�-	�b�̄⨞v�E&=ٸW�o���(���!C:똠!}[�Ow6���e#~u���0'KŒyA�i�#�"6�^�7����8x����_<�\��Q�G9s���((�\�9y���ޮ���D	�A�m�!� e0��a{�?���ޝfO[��br`T�PB��S�:���/���N6R�？��ݔ�:�|�qO��L�p��3b�4�/y�Ȉ�b����0�o�}�͟��IP�.���;4�+xۀ:����7���
e���G�S=GO��AZ����{ᒷ(�*#�N���-	9���%ǀjվ?R}�uY�i�7�������Ax����pFQ%��Ki�:Ć�`�<"GHG�G�<.P�;��|�[�����2�W�,'�N���J߷}���^� l=
]���/�F�=�ϡ�j��ztR'%����R:�&}μM��eO�~�A����ۜ�cA5sH��D ��wo���m[�Π�	�<߲ @f�Z�6x��i�!�}�%Ӽ����4x�_�*A[:y��Y�|�I�ܡ���q����g���)�?c��űd-���K��z|��Q�~덫H4����xO!_=����jT��mq4|���v��IABr��i�^�6�xb(��-49��PR���`�f=�x"���"�W�eU��r�A v�����&�?�aa��v��z�0���Z�����k�����S� F�
q4���YS�j��oi�{��؛��$O{������h\��:���]�)s,s{Ahܑ������x�O�����nD���-S*a1�:S-Z�%����^;�8�@>�� ?br��_VB��&ϣ��f�xL�RL���3":��*'�R��~Ue�������:bOjO��C{���N��3�\W�����*�t��ЊR�l��?�\"9�C}'�� �~�_���F�ꙩ�ʏC��5�)�1u���i[;����~�1t*
8	��BN��Pv��eFx�$xA������a�o+5�+�z��֢.;á9��ڙ�n�@ �#qR0��+rE䄫3��,�����{�[x~�DE䧨�3��1|�֟Mk���^���zO�\~D�x�
P��4���&S��$����`Y�Ϗ��Y����&tuu������ �-P^�W9��y5��G�n~o�����)�v⇈	�I��aX�Xl� Ǡ6����}�ܰ�6_��y��l.�Y����x5"�1� ���b,���������J��qZ�2�x�(a%fe:Մ3R��*HYpUY4�;�o�m�k.k_�����x�����t��f����R�+�~�ˑ��-e�MT3����H0��<�,=�|�1?t�LPȌ�Ub�6�H/�W�v@�i�&�O*,L�'{HNv�9b�+ę�#�KA�� [�艟�|�F�!�u䓊�6��ˠ���Sd��@s���[�J�ED}ʗ�vF�e�j�o�ӣ�B�����Q���dta�O��͖ʯ��m���^Z��mŪ�0�K����D����J>&������ʔ��.6P,�d��i`G����-�kpV+�/`QA�O+��lۜO�׮����h�w@�_�ND��(x���[�Q:�O���	Go.�@�c�x͑i�����~:�S�@r�D�^��ό�*�h��c!�#]=yV��b!q��#�Ozf%�=ΨG��!�f�΀�r�5�,�j<��ڨ�c<0��G0�Q��|�t�
9oY�!�97�k�d�Qnf����Ѡ�W�Vs�ũEw�K,�|/��p9�2�6rP͇L���׫�=�,��˭��[�6����!�!�Qwk��J	��Jɤ�������K�5��G�
�okI�)�L�;�eۘ�P��%5��L���!.,�w2����ːSI�%E��]�0��OLv��X%i�}4�����Hf�R�����6Y�cl@�f͕RJ�$}��.���\c9i�]�����L�(�
N�lw������1<=�7�]��3�Um��K͊me�{�q��YJ�:�!?�����8��)�k�1V�S�jl|K4䯳��2�/ׂ�!U�oIZ�2BZ��S�#�Yy;�P���pK޵�"��;bx�Q>}/$��|M"&nW)A�#�u�NX���_m_W
U����!v>�f�]�K<8n� f��r��Q�z��-cJ�$�t{�>��̫q��M?�����~�����6ͷ����e������ϰgwM���-�"4A@��ߞ��Cx��opѯ[4��������a� +�����(ٜN���~C�����Į����S�>�p�-�?�mcˑ7e�l>"XDr�`�!�g�׆!�/6����:fʳ�����M?��=yk��	g0>%�)^>Y7*y67�V@گ���a*�
���E�ZgG^��udsP~J�!�ASHƥ��ܲ���}��nPD��b�,^C�^�ajBG��V�g�'%/����t�.�P�J� ��p<L�!l���R9�c2<�v;i%��꜐f�q�l|V�za���_���������|�����(M�Xg5m����'�z��lCd�
����8�������Y�uQT8��7H��ȋ��K&J��/ #���0��F[��h�*�Q���.ʝRG�)�2�R����8lq+�>��sݢ��!�|sv�m�̫�6�cO��Z�w��&iz����B@~u$Y>����Z8c�3�p7Z�9�R�I���:Q݈d�i&�ǌ?+��}�T�sғȳ)$�S���?�Y��,�J�t���7g���mW�2AH<�B^g@��*la$)�ċh�_d��{?���s��6�+�
!*m�8l^��~�yz�$�G���u�����z���o�����¯���H��`ګ~|O�Vh� �&�co�zTu�.�������V�����'�^��w����Q9[��X�l�]+�o�b	H�BO���a{��v<�`�|���5޿�i��U"�7_��u:ԺnGoe]����+�-u����R��0�}e�pf�H�y;,�852�Ғ����Ef���k� ѷ�gG�m����UD��>�L�_h\Z4Q��Nw�{U�G�RE!O�|>�U���!:ԗ�ۀ2��,+B�z�Y�W�u?,�5�h1�xWHF��ɦ�Ν��D	�$�k�SVaL3'^Z �;j���"�9���I��S�+��N�t�c�|���T(�����T����"���b�����',}���}q����5��-��ϣ�
H"��*��޹��t㑺T�tA���['&�((.!���%j��7��r�&���j(ԧ��������/-���K�\C��˫�f�2���j�0lJ������a��� 6e�򿔌��/��ù�F'��н$Y.�$X�־��o�}���J�Ô��c��
T����2���d��Hv����1�Dt�\�Ǿ����⳷�T������:�;l��6-�̕��.K��33�aO�ɞ�̓�$ϐךB�2��Ϣ��X���M�#m7R��x}���]|�1H�\ҷ;��[�@�`δ|k�/��0!�8S�	9��V�k���y�a@�o�G�����{-T��(!(�>r��}e#ѽ�Pn��R?;)\�4���A�^���j֍�� ���w�*3a���o(_t�8 �B��+�/Yk�y�.���(�י��y�F2�X�\�TR~�J���j�bA	O+̹ʸi������.�q^��B�YgY���c�Z�=��k����o7N���+���pۋaBd_E�\,PR���3ч������i	�u_�����iޜH<R�Ȃֺ��۶W<,�7#(Zu�Ǜ�2���\)���
x��ŧf�E&k�l��xv���f�V	���i�S�<��^���n�\�s����������Ȏ�O1�I��a�t�6�����R����I�Y��7��_��g?$�L%o�HV$�Ĩ|��`�[�-]N�+��ϤW[��Ean��=�i[� �i�dP]~kV����,��\Q���/�q9 9s��go�v
t�D%Z�+�Iu���P�Ӫ��0���cg/|Q��%섄���Ț�%�N����q�Y
0�p�Y�s�5��䁀Ҷ���~v��r�e�c��@�ȶ�צ9�'�Ȕ�Xd�@7�d=���M4�Z��퐛b�Sc>��k�����U��d���N+�e��hO �t@����uN�c�f	�aCܳ��^P�uH�u��g�L��=I�=��B%TވH�B=N�"��)���6�
"e�����M;s���#C������_�Ɩ���x���Az�vK�R*�~�����r8��9g� iN��{�D?��[��x4�H��HZ{y�����,(�}dq�&�����['�L�@��7���귧��
عlM�p��O"������7�<0��}mǵ���Bi�b���0VV�%4k��!�{��Aa���}�%�W���;Oۡ�JJXq6uO���31���g^v���'9Wr�qS�.�7}�0*/��e�Pέ#����j)��Q�ɚ�צv��u �Sc4�u�J^$�̂����V�ʦ�V��y��܁\+���`��N\��#[���щu)��A���౓�������f�O��g\�oG��?(ņE��/l���#.�����/p�C[Ydwۍ���)x%��,���b�ꔎ^�e�lZCvޒ��E���s�VLѳ8ե�g�)bG!Sm"O�{e�Z�W�n@������^CE��,Uݔ��p����e4%Wi�_g��ݜ[d#�d���j��#�sZ	A�#BxC�Ч@�pZѐ?S�֐�ڟ���`0*��#x��~��hE�+ȑi��Iy�ڷ��s:�����դ�44�Q�h>�B�yKӝq���)�9"����v�ғɜ���N��;qআ��x~g<Si#ӓ�S7cG���,�E	�:��1*loR�z��S�{�'\6�[�ی�m������܊����V4�hv��2��\�7ؤ,�X�b��ׅ��?��yD�2��&L��"S
6]i��X�h4�9�����\�����]˘��Z�m0:>�fV�jȷ��+��j"U�-Zh)Ս^�e�uJ�W�k>5a��;f����i$\�6ۍۗ�{-k@~��pX�m7prj�c��Z|W�}qV`���m�n��� ��һ��%���©����Z�=2f��s�
a�AyvϚ6V�9� TZ��� ��0��Qr_�#���2�,�"������P�ƍ+��N��9���"ѰGp��_UK���4b���ڨI^��Q�獿6-�Hx�4��"��-3��	cu��� ���4�*G~1�0��/��]�q�����ʵ�!e����8F��#�߉��a2':E�(�����II�+}�5^osr���&���r�c��G�Q���Y|W�\6*	\g��/(�Eo���f��$�F��cY�00P:�{�Vy��>�������\��oD�[��Qc�7r^c�>/���o�����o���	��Q$B?U{c��$㟎����7��՚@��&*]>�5۷cr� 	�c|�*�����Q���e�g�Uz��m��	S�ϋ���(��;�#�I�7�ʀ;p�M\x�D�()K�B�B��NC�4(����%���,�;V���x07%����v���kD��I&Y�o�Lu�;W���n��2�ci'����l�ͼ�K���~Fc�B��%�|A 6Ñ���ƳΉ���`����RD�]�~�π��WJv�8��/�w��Ѹ� ��T���i�u�.z6��ζ%�6��2E����MQpj�
�z��8O���[>
�eW$ˊ�=��"����w���٤�+Q��j^:��'׶�yW|U`����Pd)��=j�ro�|����O�O�]eT2�A�?b��X8X��l�_�e����?�n_S����g樓��7��Y�����#��=4������q�H�QZ���?��7��u8L�,d`ROh��,H1�'z��!�M��{[[�{U;I���ǆʵc�m���Rj�+$�Z}�0���e�����4Y��� �����=�4n��Cŀ����h?kA�.y����d�v����#�#~W����/u�=�<��؀~m���#�|2��*�4gj�@�/[C�`'`�y���iE�g"��� l�����k���r��d=p�w��w� ����h)�%-e�e�n������J�:Ԭ����@_N��sf<����\���;U-�����?;�o(�)7�=vnj��^�[	�X��*\r��r�������L��2�Ғ����Lr?B3G'\�I�ec�&��%��?��,�,�.���項��>G;���y�/�S+�%��4���F+J%��4�.z`�][��G����p�)�t�w�4�ɕ�������1:GQ�^�ye���Rq��h���ڪ%�h*�۪�ǅĎ�o��'�b��g?��A����^՚2S
7{�մ��]�s+�K�(��'c��I���̋�W�}�F#x��f��<�fvk��Ր�l��b�7@���N�T�@��X��ϭ*K�Ԩ�7���᯹^і`H\�ҩ�-����*7\�6���:U9��P�&9��bP=��P��H2�N>HH�=�M5ǔ�X����@p��� I�l�$��#��)i���r�B�cw7?X]7�sՙ}��n��{\v��ӿO�v�Tow�K4`I�+%X���{��S�fQ"��{đ�R�@�?�KQ2F%�o��ᑵ������j:5A<�_��6GN�}�Xl͇ޱ4���o���Y5bc��kq����;�l,I�u1��w�.�.�"iN��?�QK~g=![�?�/�6��f��\:Z �����Vٛ��%�ԝ��c�C��1��k���Z�y�2���sS��0Af	=�o�_���c��~%�����*,=l��	����"m_8�ɒw�@J$&��[w�L0h �qœ��7�n�U��������y� ����Y����NI	qe�~����sq"^: ��N�y4݉l2 ��c��ʄ<�};/2-����hn��zдWv�յ�Vֱޥ]��f�<�~I�ul(�;dAY�"�b���.�O-$�ڀ0;=�a(G��C��6����!�`�u����4#�����(��v2x�~�JX�K��͆��-/�҇	�Ӏ�R�R'���n��N�P䈧-ȟ����~�@s��=�g�;�L8�6um򸓫٧�ƣ�/�O[N�yN.ks��Ə�z������j��{����Q �u.�>|Y���L���Bn�GT~�k/��%�"�=����i�9^�L��6^xa8�e��J�k܄PU8����g>|�>�è�(h�A�P��u5�{�z)�:0LIOj'��!{˰��Ӧw��	��m���~����c�s�t6� QL�Sn>6��@���)N���GZX��A�kw����=>ɋm<���t*�:�:O=K��+��&��L� �j� g	�7��C����`$����p'A^�8�'�T����3��6䍡Q*P����3�/x�7T_d�m+%�����o7���\��ݳ��%L+����� m�
o�mj����L�P���]�����v.��/H�J]�I�}� Kq�����ф(J�\^��:�ĳDՠ(�9�bE[ �n��nc1�T3�|&',Cr=�`�K`�鏳Y.bHN�:v��������s�%ȷ�(�gr�^�`�%'_I4E�zwb����G��A���2��K�ٌM����@�M�i��@��-�2-.�@�hv���b�\�������u��gcZf�t!��AW��1�VS�{��3�4�p=����� �3���wb�����zB�$�>#7�!�	J�6|t���`�qE�Ɵ��]��U��.���C@�;W�ר��M3�������K&=�Шpe��(��^c��f̤]x(�c�7|u�3���oZKt�%L��a����E{gf�s��<p�Q���A;�@7��u�U*�;�>�?u҇hY�����e�-��R
�P:kCl�C�M�f�A01ܮ
&���"�"�3�H#!�b} �-�i�B����J��8i�(Uʤ��G����H���tn�DIZu�ĳy�ar�4���my*���EU9ؾ�ڊ$��īփ���6@�Q�<s���|�pk_y�fP.��O��;��`�E�?"P�-�#��,��0^etR�W "!"�������B�̓f�tO4YO-9v�k+b"�r�-���H
������E����9iP��ݺ�1.&��Fn��BG-mȘ� �Jm���p���B�!��V�^��+*`�KY���#�����`f?`r=��BB>���"�ɴ+y��Nek���Tsh?2PSX�/��o_�D1�J��y�������h*۴q�VF5
�5R����KT�'C�^GD�Q�3��6G�����:ˤ�`���Y�J�x���8�~�L�hʂ���{��e�0y��f��Z6tOj/�ԉt����ҍ�h��\#aS����2����0C�:�-��6�n�FL2%��� �����"����}yj[�%V^)��R�'��7�:Z��#���U(���@]=��/(�$��T��>��8��+�6L8M9�Ry|��bZX��ܓa�b��x'��A#Y�G7^<Ƶ��:ڥ��Pd���O��;�9�����xz��j��)���:x����~�Xy�ߵ�z�ng��1k|�ˇl��ȳ�}��[IɼT�N�b��%?F�B~���N ���9�l�r�Ok�$�3w�+)c�Z@J�����3#$=��V`���5�&�U�!��F^S��A�^����|�q#���*(�u)�Ep�1���8��|���?E_(�a'�D���KD�>=0t�~(�U����r�%��L)�>�Ѐ���<�8��4��I��I��Q�=��PWw�k�<�����x~q$)�-��ou��#��2���6 ���O�@ڨ���U���������@��Ԓ}PeBT�-��yW��b��Ml����Ԇ���nz�'� p��C��o�9Bq���S�b^)(?������*h^��D�n��,V������b� ә���!z(�c/��	�Ѯ�1�ϣdz�����v���c�2�gc2�W�oS ��I~�ז֒ ���U&i����GS`��J��j�^O/	�"����E�J������5�0�+T�d�t���� ��M6�@��V�iw\g�va
e{����M*��b��� ��L<&��U�,�:kG��fo,�o>CbS�l;8��د�8��9~�6�~>65yD��(޿�����AI�.��y֏�rVU��y?q�ʮ!O���l�l0B��4mf��p��4!t�<\��֜�(B����A�O'ry��Ӆ���Q����A��S���ӎ.�&��VTxF"�"6�������$2<\(�7ֳ%s�q��(o�����d�D�*6�����
���T?Kx��|p��sD5I�jM�����P]���M�Z��L���*�o�^ �a��*�o�ڜ����8���������i9�6����^����� �7�w�H٦O'2N <,�J�xBɋV�T��=gx���d5���*���F��xx�1�c�q8i�}��0�T!�:�Y��d��o䬋'�VQ����~A����2��کM�[�`ç���!��α�V?�_�72ML����G��w!������ʖ�7b΁PB΃s"=���.�#����V#����+ޕ�ۅ���b"��d?�>reur������o"%��1\��>s��(y�p�
��G@ڭ!�j���|<BE���ݠ���&����-jǔ��y�V��Q(Q�MU�Ul�j�w�~��Uze��>�����u��P�8��A���c���.�7�A��}a��آ�kY�/��&��
�J�p�q�H���t�ݔ"]uY�|��C�� u�Kv]p��|�l\�U��~��׷�iLp�ގ"p�A�L:d�f����u&��Q�?�Ö��۝M��gl1yVx-r���F����ۡ%����S�8>w���t	BԐ��t�bq	����F�@�R�Wr� ���h�@S�/��X�G �����Z�z4�s6ؙ>�G���S�i��1���x`�����v�'�RK�����+ri1
��oI�x���Y��� j�}�-LE�u���=��q�{S��w�'M���L�+�B�*�R>a��Ԓ+b�zUk e��6��*�y#����-'p�n����A�F���f�}�r~�*)�e�;�u?��h�E�b�>-ӣ|:����
<�э�R����'�S�p8Vr�Z5��<�]k�[Vs�E��!�%�a�2��'ǿ��/�N�z�b.�g�J���t���.���m����9-���ە4�V�f-��ſ4ST����Di�ܱm�Y�1v	klxk��2�o��#��T�x�i���EAO���ȃ��[�\{!�nO	"d����t�[�ք��G�V$���m���~e�۳�@h�`�wٲP^��AAr�+oiO%�S�1��R��w�ơ��� G�9����ǜƼ���{�3_�}Tv�K�`g�gl.��߄	3�aI�N`=���E��:��K[�UY��)�	���(`���I�7#��|r_<2I�;\W�r�d�qB�8P���qH�ឪrt�y�,��IEfƝK������px-�c��%%���["(QZ�(a�&ylVc$ ӛ��>����Vu��T�b�ܠ}:�<��&����k ��s_?�k�%ϱPV���\��\1�z��i�j�@�� ��E�/��č@����~�KR�<He�J'���x"d�C�Xo�Hm����e���-25����Uxf��Cæ��_��.,)�=
CzL��^؜5��H��+�0T&Q� ��.�d*;�]sC`��	$�lnޫ�4ǁЩ�j�=��v\.�����a��v�+��.��r�`*�ϥi���sڜR�yE����x����3;~�k6�fj���F���V����j�᭧��U�q�(J7ť떢�;����8�R?�<E�ER#P�I�;9��b��y��Q�� �G'���h��2�ߏ6&���8����.0-��;<��J�d)��b��ZI�,��O�5�|^�\196�4�Z��lR��N�tz�| 2���S&M�a�	!Ջb�{IM��t�|�Fh�W{���}��iy::��Nќ�����@�$̭8.�K'1�n�o�Qo������h"���ϒW}c zLu���0зY�j'Dd0%mV���17H���X �T����h�A���~7e`�B(U/@�Lj��؂7ѝ��gw�S7 7� ����l�u߬��v��]E-�8ޓ���x�ЃZe��ܮ��)c���u~�p1WZ�,@t���/�ɑ@C疸��<�l;�-Q���;��~��Y��<�G�u[�ׇÊ:���k�gQS�3Wv9�ݥ&�
�7�S�L���#(�P�q�����m�����y:�\�Eµ6ug^��,�7�2uI��$U�m�oy��̿>!8Ʃ�j;�o<'" �%�~Rq���k_�Q@X{���0�݆�w�	��Y��3���;1��ȣ9��賸8���=�
�iS��~����^fPҨ�_!r��ԤoO���'�P[\,�9�S
����>���_�e�Z7T:@)�%�l��"hlN����o �1�7m�8e}s�!�U6G��]��=;"/�d�$[��j��"�S)�,��0�Enp���хPB+�ɹ��͍�F� �c �X0K�+�Ug1�%I�=UЅ1?_х��T��k�է�g��B�!W)z9rk�������P���EUX�������^��'Fs�y4����$�fDW���\t�+��љG�Q
�$�u�<����G������6�8@�Zާ�A�.�շhK���J�0SXJ���ĥ]ŗ�� b��BGX�����^_�^�W�b��}[�����ie�|�
l�fgUCrL=C��7XJ�mt␳�&$<XW)�e�;qأ(���`㸃�[�|8>>j,��^��f�a������]��n8�-�U.�Cͤ!@xc����f��y"��ƙ��o����e+�X6���l`W�
��|_�)[֚5��G:�� ֚jt�����S�=t ���3Լ&,��k�ퟦ<%�h����^��̤|G{�Q&pL�7WZ��,��×'k�X4oHrA4��;��ϢA"3��MVi�.'�'i��hTW�yڪ������a��k\��G�0�b;��J�\�P>c�[�@R���
TWۻ�F�[�q��Q�xo�ȇ��&n9F������u�bz�S��unӺ��d��gL���d���(欳^�B�G��M���K��U����wط.��p�=����b��+����%W1bo�ƌ�p�?���yƄ�ŀ3���[^�c��u�o�_�� �����X�����},�C�'���WU� >��^�d�]��J�3��X�d��E��h9,�kAVՙ-����kP������x����
�E�m-C�7Nu��Z�}�Ԕ�VMfc�(�����:���o3	� (��)�P��	�༔��s-���.�U���Y���7~;�Y�Erǩo�t���N�}��O�
��]�c��0?�6�c��rd�"Q���4 ��w�u���y��b@�?Gk4�+W}���D��眫c�Pw�7�
�%cM���Yu�m��Q7Q�����ʑ�U(M��ݐ��LH�oJS��<�y ���/�,�x���ݩ�Հ3��CPJF6�%ǧ	�^�7��R���7�%f��R��0[L.�Ǡ?�|�%>��}B���B� �Q�x�`��{���I�HC�M�����2:U�md7Ń��w��d�T6��J�k�2��K@�|��5�rbS��/��/Y�t.[\p�F@�dY&,FT;�𺇰R����x�%C�3X�䏀� VɩO�T���R ��٬B'[��R�oTi�P�j}��5�� �t�w:|�<�7\y�[��Os��+����!�+dV�J˦H�|K������a
i �b������H���Iv�z�yM�����Ȋ䯦�8:�j9����x&A�y�ʋ5��H��%l�X�_�k�s��	9p�-�{��r�L�S-e�)���qp%xcy�]�t�/�F]u���<#F^?��X�U5���9�2Y���0_�>%�3y}�(�^c0і �pp��J�k�G�(��5�+���&�~X4r%Ό�I�6&8N4�*k,��7��j;����J���u���b�T98��D+��I��2AD#U�����A��֯�`bK1����9*�=�p
�����ʏ�5 ?h�| p�}B����oW!ܾU>I� ,Z�݆{��7]��0Ʃ�JiZ�R��\3��I�2Iy��_�ge�ϯ��!�����<�qN1^u����3)R��\fg�M����e�	c�iL9xtxB!R�A�:4p@p��,�$�b�s�0羷��?@k��9��x�u[J�6�|�׉����@yr��<���"K�t�5���x%J4|!}Εgr����z-�s��t>��u�r���r0�qV�^Ȭl�_2�����X��պ�:.�$V���\~����O �T��H�����ԝ�s�Z'dPy��Oqh]L����G����e	���&�I�ϭ���Ɵ�|m�XW����y8��d�d��_
�����֥�f}���x�Ă0k��Ipl�_c�H ��pp�m���'q1=�d�뗭랉���$xzo��D�Ώ[[�8D�
��ɀ�Sﾛ=�K�Ğx��t��%u����9{��+FD�;ߖ�O�� �a�5�dC���=3��nP#_-u�Јّ�pP�t���e>]*�z!]���r�ܪ�,��R&y�5���P���L�p�7lb��<m����ƥ�bwG0�@��Hա�{��-��p #:�����pβE�R�`�c�<�,�L+�Q�$�W�_����=�oH���:A��Y��;�	�@���r�hD"pE����͙�(��Ƽ�e���l�QB+��;L�o݉���z;-�i�(����.����̃��"�����C$��<���������/�C��l���_/�%�󮻗�q֠χѐ���gB�&X� Qp��`�VE�RDK��<��y�],9�}��%˳���_���b�И'dU����w���F��t�i�#<67~��a��I+� ������z�'�e�'�Y�}��'0�s4����$��?��o,!��mzs6&�|5
�>7�'󩏘�^|�]�^��������|E,��.[�6�V�kK�����ٜ�\U�������'\�O��j��_6B�[�����mI�^�Օ��d�ȋv�-~�ن0\N0�4)Nj��n�k�n��n2��4B�96�6�e�o�.�L��.3���J�Z��
�Z�Us��w��٭�۩��1X,cl-�dlK���>���m�O�k��J$�у�JJ���1�J��'9'����[�$~oRd�Յ
'���=č�t��a����OLO�s:���t��!�\�}�"��~�7u��>�:b��VR�QJ��⛨�%ڥ�ؕ��YF?�oa�7v����.*�R��K
����|'�z�Wi���0��O��u.���N����co��7tZN�%k��!�J'+��S�!�]*��4�T��m��4k,�<W�#,b��٥S���"IQ��t��
�W[����"���
�8/Z��<�Ҫ�$�����w�o~�'bѡ0���9�N�@���n��w�����[5��l?ֿ�]���?���&��rb���]�{�>�OG�$��o���7������P�	P4E@�T`5��_yv-S+�L��i���ao�N�`��&������ϴ���$,lܾ����R�߅��e�S�P�M����dh�e��]�%|�ڛ@��	;�C:iUg����o�!vn�4%n����~��¸��
C���ef
���Ǯ8Ǿj��k0����78��귖jLgƼ$2On�I�Ӏ0Ius����VJ���W�V�a�-@� 4S��j�h��y�K�>yk�\�;T��4�5�h�&tP���ב�C���P����n�H:�Tkw�#,��5_NNW���Ob}�7�X��4���ȧ����<�6��]\rc�!���Hn�����c��y�k��(��gwi�z�/��b���biI�ހ��%}h���4�����N�?&��1���2S�S1^�{���6�(��Sc�F�DR�i�	j����
�}�؍�������?���]�/L	�&��/�R����F�w����aL���9��k�Y�~7���㵈 ���2�ƘZ�W�Ra�{��Aڕ��Y*�ǧ^3�=�}�A�45�!���.y��#�#G:�ٲ��JHC�!`�XT�ۦ�=�
^fK~1�a�({�A�@�k��uWr����֣֞����əغ�������sڋr���ws��L�*.%�%�6�g�x�z0`��cʚ�>�^a���%=����q��0.^SJ���:�/JJx?6o:�i�D��j��zzv�p4��<]͞�h8 &G�
���ۿٸ�������|�"��,�#-@�el�h���gT�`��~���SvK�=�p(�̴�����2I�Pа��I�j����
eG�����T
!9_*�Tz�^��3�L^&�)�?�6F��q�dV���Vw2%8��"��̷F�u|��yߛ��D�Qyw��cA	;f~�7�����?ؘL���t�L�/��9��k�Ot����������x�	.�D/�8ʺ�Q��S�6C��)_��0�j���E� �4��H8Η||����q�ꖨ�~N���{�Y�J���7	� xP00���]&�B��f�'*�&	�+K՞"#y��40%�rR��%����Ј��Xa�#���Aԃ��Nh|��z�{w0���i�!(7;@ް�
�_D�s�����ȑ�5��R��d��0#��2f��ȅ�M�Z�&��u�&��j4���|+#.C�ɷ�U���HB�������s%���cf�ˢ�Z*���pe�Z�I���&3V����$��A�p�m����O�Jv~�����������Dj�]�<ˇԙ%��_������2��ޱ����%�e�M��u��3�NL�q�I`S��6Eg�����|��G|��zh[��:=�ѿ��y���(n�(%�0�=�� 6�<�����`�y���������q�G��$qe�:�}�U�7rY	�^㳻���3]*�cQ|�"���W�;�Y�vf�:������TG$�?��=��VL7TqH��a��r"���Jfs���@��͵V�3���.��Q�Z�̤�0�R,�	��)�Z]�O֮�L9-���w2.Uj]q�6��t^5�y������R6�,���0b�{�=�f����hxqP2�� i��'�((��7K��hx�ʀ����o	po0�7��c �0�/���wi���h8����C�,��8��=���A�㫮z�p9��d�]�Ș@IT�<A7����$�j1LVE.b��������龳&C��e�!�d31��)�v��2%ou�z�­M�Z�J�l�}��?�0���BY��P�N���O�u�7�B;ɥV�߇*��p�#��Kf���"�If~�L0�)Ԟ;�8����>â�7O�bLN�Yc|yvgٞQ�OQ�@ܖ;
��T*Za9�����F�l?��X����t����(mus��暳)�	PI�L9!ŖZ�$/���(I�ZWM蔫�ȷRv�Q,�I�a�[�7X��ru���ܹ-j6���HP����R���N*t�*s$I������Y5m2/�,nrk&#s�C��O��<sRJ��0&jAb9�ӹ|Z\ϒ7��Ӧ�0B���mi�Deq7��I�c]�/�	:�t�x~����i���(���K4��6��|�P-�1����w��v9#�-�Fo��������ų�s�˧ض/�9t�#Yز����n���ق���L�z�����7{����Gy?�q�নu�pc���Z}��['���3���ϓQ~�Q�1��I�*�KЮ�1���\����Ĳh��֚_A/�y�XR�)��n:i�2���a�K4�\�/�M»H0x|��|8ژ����r���+��(/�k��o�ާ�+�����|��?�%-� W�0S�v��i����Δe�0�kC޺H�ai����#	X��c<rIֻF{����_9�r4)� ��D���h��o%{(#��()ɦ��"zHR:1=?(Ƌ���{9C�E��E��T�F
��#��d�x�K�MoཱུDͷ�6-Aq�|�������o����	-Ccx�.+�b�^cL<"EX��"ڙ.��:��>x�v��!CTQ��f����9��\Ӫ�4GN�<��������Uo8tn�}�Ve3�V݉�/�L)�S\<�Δ.�o^� Q��z�N7��\��Q����Q��G�Q=�v��MRf
/[�&Kk"��@D�4�z,�K���Ҙ����e�:�
�j�J?�����Ƥ�������9�eG�f�1t�����w貿$��]��jy�R�f�:�S�5p�&N��d�dn�_�p�}������ =�=;1%�f��3�u;���	�5��9�%��l���L(���G�US�zDo��uM�7a.&���Ϭ�]�h~�p9�V���-�Y�#�:�Q��;�ȷ
1�s��1ųXR>mQk~��I�0�m��2�=	%gm!��Uƍ|MDr(�ƥjg��Mz�s=����~��DS� 8��ʑ��ގ��w֖h�l;��a�6{�Z�Ԑq��B��@&���x��腒�@za)�S$p�)C��D����w���܌��-��_(�&���Jo��M��_L;Amt����DtS|Ƨ0�=tk�5Y�6��<��KR���骐[gE2��v|��		���F�]�\�'02�Q�S�IzZ�"�YU��/O�H����h\�䬽� �U!.�k�;��A���oe�1�kD�p�v*Uz쮞B�?�j!<���m�%m3�Kz��ʓ6���[ ��#��Xh���Z��V�
��<��E��@����=�&�*f�ۅ�{ӇS��@<�n+��:{��A�P�?]���t��NEߋ���Yk^瘲]�W�ǜ����o��{~����Wg�7dV7gX�����~g75լe!�2(��}�^��#���2�>�"Ȟ1Yro׌f�Vފ��x��]_���Z�$Aщ�C/CQ��9&1���"�贸8�ص̨9�X����ʏa��;'��._��&ЃZ��:/��\����D>��.��BJ�P%#�x83:�'�%�x'�	|����3�c��Z�Z���!?I[���� �eO#�������#����Y��g�cY�;D�{q�ҕ�vs�/�`���]�A%ys>�ꗈ-O�p}�Ev��o}@��Tٍ���D�W0��s��ض1���|����'LgMU[kJ���9�^��������i
>�2#�<@�q�R��V�˾��;s
���s~��8��KQ��օ̌�i��2v��|���Q�Q�jK�cA���#9:�-�T��}�{Ɣl��\�G�]��t	�[�gI�؎5��Q>����1Y�矃����TS�(v#���(8/>)����Dݙt%�ÏKČ9 ���S�����cY�	#��0R�綸�I��ԯ�����.�C�sr/��#���ʯ۸���_?mnNw%��1k`�P�|5'��rg���G�=f��
o�,t�d-���bZ�G�9�^� �cA;V��rם1Y!�
6)R��hc��dTW�+����}���vXP;ۤ��,�d���%�W�~��������1�u��̓��}�
~yq�u��41q՜"p�r���O`��}�i�u1�]U��)4F����Z��ɌL��5��iM�fFD=7�M�֛��Fd&�'�BC�7������2�nt y�E�k���j|�|lǷ�өB!���+	Lqo��^V��Z�ж�oʝ��)�(�����)�lv s����^����Ⱥ����y�O{���H{!-��\��E2���1�ԯ�ea�q͚�-�q������^��!�Ms��f���E�����oƬ
o��iw��/�IT��Ҿ��Ʃ<ћ($�r���'6��ܭ�]�h����K�������~��L��j���B��	�Ÿ�Ҥ�aY�F�;y��b܁���>g�"�ۻ1@ ��T7�kA}3��5��<B����#���u6�*��Ͽ���Wr�IL[G��������3Fhdm[*F!�۔����-g�m3c�r��	����2X?ޙ���{ܨ���Tq�޾��р�c��%<<��7�V􀬮V��9(⡄�ٰ�B���h^��4n��DI���au�f_��q���.�,(��'GC�TveN�O�����5����峿6^'8C�rk��~#~8kF.F�������rˮ� ����y�}����i�G�b����)*�G˴�ь�3&��W.� -����Ԭ���鱮����[�������i�h��,�A2�_��:˝�)5�|�Ȟ���𧯇'����z*;(�k3��hS�ݜ�h_�V&��B5�mL�0���
��vx���Z#�,Y;�0�x�@l����P�t�����lP�䏵]����9����H�����~$�/Xe;�tYd[�J(�Z f�&�S��t����X��S��atX�Q}�ޚ�v��z�B�nsޫ�.���'��M~��\�6�tJe�N7zc��릮O�E�8� �i)K噇OJV��B���~�~;"�ȉ:	�s]1N�;����r��C<��XP���j���]\]O�.���9�"����dK%����F>�(_��-��6Ԫ!�&x��'����z&�ůl]U�/�:-u��ă0qg��d�L�C=��`�	���t2�D!�{��K�Ϧ��8]q���c*�T�Ѝ@����#U�A,P.�UU��	/��%S�̱�%�#�8<)����L� ��oº����Fw�]�]�U�o%+d �!Tt�K�BL��L��)�h����ͭ��-L�X�)���,P���=G�@�u�`�C�<�;s0|�O�Y�;��G�hXa(��{�'��9]�[�v6?�	�~J��3���Ō�?�U �kt������&9yk%�/�m�z�@�s�@�qW6eG=�@�Z��_
gTx���P&o�
{]
��n�ʧO��R?���t���
a����8�s��/Gp�2ܘ����Ǘ�H�4� E|��[)�y�h}?�t&��M�0���D:�\_��T=;+�sڽ�T8��Dd�D
�a����Ǎ��S�c�0�\�p�?7G�Cnk����c�eYż!������vr��!��C���W&)�ʵ���0������� wˎ�)�B�Od~���
e+�3�-�'aI_�k�rȒ>��X8j�����
���^�9�i���v�H�ǭN��6��3���0:�g�H8���C��L(H��(H����V�e������F��N:/�2��2v]F��A0$����Uo��<�
<���|=��[��[{}ƚ�}I�*��c��m,�f��E�(�,����?��t�L��Kp�CL5j!�9��6e�����p�j����ij	���Ҥ�ڜ;�(�p��2sc�hc�� ���Wq0�0��5^G9WV��O{�9���{||d&�7߁�2Ry�ɥؙ�oasT��%~h�ϛ*Ϗ
�.�h�	7b��� ��W���a��|S5�7����A��livf��u[�{�8���a�͵P�$�)�����wpFs~
]��FK9��#��N��v.`Փ���ߍHHJ�q˚l5çF�%�A�'���B��x���J"F��>I��L.ua������b�z��<�
�D�}q��lis<J��� �17F�u��
U��,����[4�(*��v��ppRUjB�k}��^�L�9̯(iA@��?���!��.�9���5wvQ����~*t%D#�,4��[��񇀒��v9���
�� ��}���)]���!�e��p���X���}#$���N
0�u��kl�{� ęQ�J�TcjN�3��w+��f Oe���H���f�}���2qZ1���񯸏a9�\�cr�RI�V�h5��˫a�>w������j�ST���|��0�4�|� �O��7�.dc_�PR��2+,���dľ~q�F��4��"�V��e�����j@_�'���R�Y<�����GL���1�f�L���p�"c�| �8�ˡ���1q��*���͏}u�[ʿ�Y}��-�2kKq�k�$�5}4R�đ��.�C��Vɹ@��L�uJ�[�����
�`����p�28[�nͩ2M8&.�����f�B�9_�I���,�7^H'I�pC�^�i��eg�z?�5U�k"��gLn}H����P���1�O�kFB����:z��i�����H��&�= ?��^^b�um�OK*��S4���(K#���j}������ ����Tm���� ��c_%@���e����ʦ@������q�����@�a�B��aE��ɽ7���>�u&�N\>�I:"׆0B
x|��l\�s�*�MsS����4=�)w��"�<��˓� 
�Ss&��\�ﻥlD�G�H'lρ��3�r�ŦAo��tI���%K����͛.Õ�#[&p��������4(_��B|�-�M(<�sp���v���N��d�׷V����<�Wᰵ��{��
��;���{Jxካ6o�䊖���zRP�j��uڬ	|���=�W�t�s��`ƌ�g�ϗ��Ug�E�v�Q�+�9ڎk�-B����l��A�U>����W�ӛ4���q��^��_Mt�X�#��<K��elo�ՀcR��6N
���#k��"�㵆;�9�O�z�&yׯR�����F�3�`��>��u	;�q�L ��[�ԗK4iw�3X蘒�"_�og�C�-��*�U<��V8NE]4O;=�چ_����%t�[Yn�������e ����O[�ߊiks^`	L߹�W�pۣ;��g�JY��I�f2h�$�n �h�¹�|�+�����^ؙ��8)h:�$<p�"���_��"XW&me�Uz� �S*6$�ǠF����3*9F`�2����OtږjC��n�,������VW�H}b��t��䳑��A9�v�zć?aYR��{__��ZߡT!�_����c;^U��G�YB�F��S_�k-�rŀW�.�oۺi}�Jī�8�ݒ�Ȩ�n
�i@=�����.!B��ӆ��3���dΤ5vJ�r7	��dD�$^�1|O�����W>�P�l�XWl�$�AA�,h4l��]dm�u�K�C�3h�*����LN�;������<��Z��Jz���ώ�Xq�GMp(L�9
pUhP��ﲫ��w,6��:��Nm��ؽ?��Ŝy�bl��0܇Hv)�O��8w��Z�G$�$~=�(�jīg8�;ō�>�P�!���	f"�2F�������q�;�e��wFQy��N��͋�$m��P��F��m���&Œ�����w(���ڔPxX�(�	�keh`s�D,pƛ1ȂK�q��9N{k,�4��0���x���L�\�x!\�R�`���ťH�����,{Nq�6�%�ң��pL��Mr����e�-w��a%�|А*�^qH^�I��&Oݔǹ��ܿ��f���S� V���t�8ƾ�ч�|��z5�K �6vG���
�|zA���7#�0ѩ��=�v�ϊKW76�c�Q8���f�%���2��Z�ɐa�"$�Hk.�7u�
/sTr�(J�`�N|$ 2׎��Cl�!��~ݜ�
��t7�J{G8��f�?*��40��Yx-��<\�tK���CN�0�]��j2��Έݤ�2���� ��Ē�3U\�EJb��Xښ���?f/���P>	G��c��0�S����c��EB `�,�eI":[����������<���"�Ӹh���¤-��x7�Y�d�ٖ�]B�@{G���/�	}[�)`
�܅�E_MO�	�g�P�m�t"��X��~�p|�#8��x
�+ȋu�ăc���}�~� {��%y�J�C�D<�6��.�b�O:>��6X�W�~�/�J�/�X�i�o����ڄ'����晐[_���ǉ5:�8�xF~آ�V+Sa�k�� �F���:z���O^��c�A�Y_ _�qv@sɜ�ԕ�gS���b��1(˦t�vM�QJ��0���=�[x��fv�tufG2[A�=��x��	z�cZj������i~�A��V�j�F���e����jc�/LT]�/E5��H)(c���17Tk*�\����Y��:A�u��K�1��"xj)��|��~z
hn��e�Tt(����q���5�?�g��R���YRʯ��-z	���ẏ�E�N��QE�K)���n��b4�{uO*.&��*B΅`狵�
nd�®��rM'Hc�A�p��b�vZ�0K�\I#_��	�M�{<b�E���ت����h�08e�߸a�E"�����3��}�>�!���_{R�������X��^$K�8-��]X9���l/8��h@bY�R!pZ4�*�Z����+�Z�HOBS����>����4�����g�!e��r�!"Y�����j'�!�Cѹ�͵��-.#�f�����'$����wq�Ps[c�՘��5bhb�(g%��H��孨G1%75���.�y����.�s�r����7ZeBQ�*+i��3��;�t���F#�WR��6� Z+#��O<�c��cW���W�T�m����M��z�u��W�����!אVom:<��J(��Aۆll�
����u��݋/2du>3wb��vd(�&���_"@1�&/`�����.u��3«e�W���<��EA�����F�%F�J�J�
��lĒF��ߧ-1�A�/ô 4�{4�|�ca�y��s�1�?Ӥ�V�ġGr�����'
���m�W���Pq/�S :گtA�g�|��WS�:�;�~��_[�'�>��׹�+���r^�!�����D�mm.���������`�x�;LF"6�*�Gԉ�s�������1+ǔ*j�&��?���6Ҋ`}���3O��T~A�5�����=/d7�ØϦ�.�A$P���k�l��Մ��Q��`ڗ���t|^nW]�$�n�����
�X�d֫/&pe�;�>�� �Jif�-R_}��ɴ�3��"�"�Z<~�x��������Q��D�2@�x��5
���K�	�z�����'髜mM�%m�%6{h݄��}�'�)�\\y�V��y.�{f*O�d�RP%�z��C�9��\g8�ʬ�n�׏�g���%Tr.��@�z]S��
F�����b+�s�5�S4#���4��S��3�YҜ��'�(�N��ѳ�=�G���!*��%gׇ��O`���y!W^ER៲"4�D�٦"�ݤ�k4���ou�mo�Y.^��f��ǥx�ӦЗ�6���𲌍�?�y��M縠�j��]0�m����9��BN�x��s<���p�a�� �~��?A����(�u�0)���F�9.6�Sj(��}S�E��r��.��4{�0NK�`��Hw�Wa��7�`[�X�f�#;G��Ɖ: �Y�C�X�M���	?j�k��ۻ��]�[VJ�P&��5�NW�n�ܴ�݅��X%��wZY2a�y�«��DԌA���e+���� 6bL8���o�����kSgn�u��
�`J�竘� ��/<��&�KS��Q��*3A3������U�w�Fd��/;��
iiT�A�<��X5�>dJ��zw��$��J��@F	��.���A��~��}#Ex�Kˠ�gr��7}�~�Bnw���@b�|MI�1�X	���!�6�)��ob�J#�[��ʩ�R`�OP�yL�5���Uv�m{�}ю5r��f�ơ4�6�|�҃;�U��rpx@ �84�n�J3M���}��(6 �q)%5���y��>dthͼe	�W�������Vֻ����SxL;���%{��3t��	�v���°����ݰ���Mku��+�p���,d�2^��`l���ȻTPch8o;5k��N:b���ʯ{�]�I��0����DY@���k�"&�����u�,���Q<�ސ���E��S#��P.�
4�g�k����}�P�_2�:V���НVN��d����'O3PP堆H�}��5�9���H�o�6����N	ə����S!�A���J!��$OfWO�2)p����q�9�*y���~��Im(����A<m}}wkrMش��_��9�������y����	Kp(�+� � w�j�g��x����1r���O�-;u����*:P.����oҧ�� �e42�h���%:�{�'�F���@n��]5����}ժsZ�P|�lXs����X�+�=u�3d��6���$	랪�.�n���⠅ި*���Ǜo��s�q{4�wH���T�={�؂E߱�a#���ۈ�g����3&���$�S,pf��'(�k���S�t�å_��b�t$�6�
�])������%�9P��0��
$[�X=�؋:�m������{�h�À��+uiT��߲�x���D��A�oeGO��l=G63w�$hH��;�3��aoR]yw�I3�}Lx��ǔ^�-b=�/��.veF=����8�Q�y3�(�7��g}�m
��` �.Pa���78QD g܏�i���7�&���E�]���1��"q�J�Xr>6����>h�rm��Uѭ(�폕�͌�@�V�J�Wh��W��c������2���vOAoL -R5����y�CwS����ZB�E��if�*�ĕ
`}�%.��vI���ݷi��J�8vܯ�莲�
_�O9Ɍ!�WI\&���V>!�v+^I����6�1P4F�j�~���Vb�g
sr8/�Ѐ��k@��M�i�:��=�!ژh������b�:���e��Ջjx�A�$�K�����M�{�|���p��@�f�?�>��*X�L�����{Q@�$]�jMc�>s��U�2��bdH3)Y��Jz����R��"q��-0��ΰ����~ )�f7i�y&d�<ɾ�߳�4�o��#�A���h}K>V��96�,:�&}��k��K��=tv
fu�{�������ⳕH#
��o���>��ĝ��N[F.`&�m�zd'��
#p�����;d��N���_�~W�6�O�8i|t����.��gW�I��wl��"�3i�si�wG�Zn�}�!'��C���_����xO0O�Ѩv�UL�uB�A��߀	�{����_IG#�� �����-V[����\1 ~1�"�<W>��'a�`R�6����Q23�N<4ٹ%@�S�7c��j	B,!�]!=�=��^1 �������۞&��{�cA��3:\��2|�-�S�~��b��hJ&0 0<�:x%�>j8  צ	��$�tX�R��a�ՎK��x�t��"n0���K�}A�jɁK��;)qJt��V���d�N��g��MYz�Ul��7�O!�Zh��
r��<^�?Zku�)e��t��vv�y~Y�q�EHs
q��)���	��&X�PD������;�VL�y�`x�Jܽ�#x����"Z�����>[E�/�r��i��j�D�o��a���NvlS�$F!0/���x��yB��"���څ��H��&�\�w�k�_�!`�PB)��������Z������ɥ���o���U�c�uW��ݙ>�q��z��;��Rym_;6�P��asխ; ��cNJy��胠����=�M�6%�7F�]Z6ߩЂ�ҝMC�R�-A\�gW���<�8l��ϤY}����Ci���������oWz ^r�0l�ұ��	9�&�L��hB��\[p��`e�Y��D�}�Dw��HMO|#�����"�1�O��k�m��V���(|e"�R�P��9���ь�Ӫ7B��sŻ��!�_H��l�������s1%v_��
Ŕ����J�La��ul�=� �`W.������s,M_{����К�h�H2eZ��u�Yw NN��f�-���*r��=%,�S ����`d虻A�,���5Gb2��T��N4A��K��|�uљ9sw�V-៦9V�/2/�>=k�e(�_����m�F��fl�h�o���n���Gʢ���_ �.$�X0z�-yߚP��
1��a��7��!�!���Y͖�%ƨd�\mjdz�$���37he��Wz����5�	���,8�R
���x��:e'�P͙�@O���U�'T��0�w�z�yb����yV�y��S��F�-C4�����E$�!Z{�Ka�M�"���ey��|ܴ��0�}xT�Н��B2oNj6�\�V�rkr��3ߓ$>g�S�h�`ї=k��ost�mpȔ� 4�B\oԼ�1c>�~�<la�|���%�Z�r[3�ǥ�.	����2�9�o�AЛ��t`�����#&�-�����E`)��l*_E7������.$�,td��˯_>�H5�g�7��.2B��a<�׍����p*w�s3d�R}�&^07�N�����!ubTĈ��e��������*�5oC<����Y	юYi�G����]Uq�V��Qy	z��k9HM ��OS�U�/T6��v �-�.�MA�Ʃ`ygV��r�F�P��QR�)7��cC%E���^9��)p/'��*�Q �/�ۖ�efU�Qf�>w>�, ��2)5b�.�ޮ3m�?�%��������t�X�E�؍��a�n8y^��Z))�G��mm8��|1�fS�3"��,nQ���SM��P���y�����!L���*��b�v��20Ŋu"�S�AK���x�a3�r�WٙѬ((	)�� $���AY%E,��> _���s˶�Tg1��~Z�r��BT�c�˝
X1�m���#�a��KAf�� ��"9��7�uHf�/���a*W.����U1h�`�(�x?�Ղx�0q��N�C�@��y�B��l�[��~I�*�ܚ�J�A�Z�ND�3��d�N=ܫ�{W�����m�-�Ų񂂽i�_�tX�-+�DLR��cYn���	���R�~�����/\�-
��w��J�ſ���N��º���P p��^�{��P��n��Ȓ�Nͨ·��R�]W2�p��8�R��|[P"W�W�3Q��1��c&"wAx�l]�L1�`�e�.RL���N���C֔#L�:8҄1�r�����Hn�B+��u�³c!��+I���MZ2�:"�S�3z�x��p%�����n�������ի�`��������2�b�͋Br:!��s�ﮪe��*�+7bx�*���{���$�� ���$H��Wܑie_H�-���QK�Ǘu�#�߄�0�^����n�g�X�g� �\��AR*��Q\��n�����Ze=p5/��l*����/�����T�uXl����y{�À�:ą��ڂ��݌�cl54�����F�@��or*�Q���63�7�Rt���щ��`��V�����ϖ����x"n.��V4��U�u�Z���32���GK1��$u�Hv�����s�Sc�w9�eZZ��G�~�A���FM�����/��l�pPX�~�IL���:�k��VAS������q���u�ڎ19�H��6wM��	a�zɐ����>�	���B�ϻ%�J�h�*�e��'0�z��=|8�|�0P���`d ��vM��0�&�t���J_jy~bS����
sof�vyH;-�K�h����od�S]��
����ϹB�=x" p�A����]���Ӡ[�~����KM����7�d+o��1�t����
�1��tK��d�&��Ī]u���c$�"$"`�������+謤ڊU��8gw�z��ٝʻ���H��^I�ϸ�5��糙�V0E�{�F.Krt�OT���/?� ���P���tb���q,Q��)�c�����S���I�#�ﱰL���l��˗>�0@ I��5p_xɬ��<2��P�nff��[,�8w�x5�B
��s���CS�t���z�Re0璙`|?�s>'bgF�'�nj�����(�_��"�2w�KX�΄0k����N�0/w}��XFu���t�13��T�_��jr����/{ !�xzŤB$:Q�o��ǲso��{�eu���Y?��G��i�i�7����^�$S�P��A���d��Kk�G[͝r�S�7
�������8�u�y�]D.mp�����4��e�Q�v^�N��D(q����0(�wip>:@�G�S�n�r��^�7"�;�
8ّ�C�E�B��AT�6KM����M��V�{m�T&�T�~O]Q=��uW�lC�l���[K�Z\�~N�~�:O���Q��R]_��饼/iX�ءHg��n�\Zl�^�-T��,ә{��|���[�u�KV�������R����Mk^��s=d�%�CS1�09��˴�T�b��{�oy�<eZ�`N���zl`5��om�(���ܜw����ldB,��kH1�[G��O	��  W�K9����+�*x�����Onf���E�	J~7FW��5$_�7�n-�����g-��uM=��Ҵ���� |�(�Wp� ����6���<���f��D�u�f�n�=I�0��L�G�`��p��.�G�[E��ay����a�.'-q��-���R˅�?��v���-��R.���˟ '
����/���*J d{ۇ։��!d2hnM��u���/�:�h5 �S�ga�Q,���'}/k�,�WDb!q�i��̠%��m"`GC|;34��_ޣ!g�1�2U=LR�A��ԥч�҂�&r+��:`��JI�gN�B��c%N``�>��+���E���`9_WD�iEk�`�gp�H�lv�PVG_�_ep��������[j(㱞e���]�x8i%��PzbV���rv
�'�l<>��.��@Tֽ�[��M�c�p������Y�N�ᖆ�Y�?���=�^�U��;y'c�˞uu9�����|��Kۙ��ە�5�����L��z���uaI�Sdߥ��,ࡎ4�z�ܞ�_KqX`�V#6+	��~w[��@��F|��'M�(�P1R_��	�\���]�pu�k]�;q�P
|��1��Z�d�D�@��*�d�J���һ��!<{\z�� >������K����r�n鄖�뱞y��-�Xe�5b$�p���6�M%.W��kڊ{�ф+�����*U�� �K�g�%pCS�AtŰ,W��u8S% 5O�������ücHY�x���5D^CG�	��l���)��4 lڇ�1;�����&��u�rz5!O���}NQPd6���"aܸ)W�u��)	��Q�G�FJ��7&O��0�_�`ޥ������8�F%>0p��|,���H��Kʳ8�͐"��Tj~X|֒vI{�}��7�B��LhL��qx� I��J@�^�"���}�~�ɐ�`P7\�:v�l��w6��o�{B��������w77�N6�ΐ�n��n������E�J�_��p���aA�hF@�O����i|'��6:�/z���j�����ñu�RrN�ɳl�5>������=E;�G�N�j�
�G�3R#gh��i��� ��n\�p��.���v��=�Q*.
�X&����������\� �!c�R'T`��7��.,���yʛ��Y�G?w����a?��~y�5\�m�{�r�^�ls�A�<��n��~F�h���xJ]{�z ��Ӯ�lQ�[�i�l+P7�����<�J�#��g,"+
`��,:��F"��Ϸ{�I��hd���	[�@�@3s�Y]l鞱O���j�&�o��'Y?*޶�R���ٻ��3�$5��<�M!��x�[U���G��q[��.i_�]�U-]�����?������|��z��0�*�A���?N�UV<zm�R�&�k��㐐uq��J��w]��t��I�<'B��uj�W��[XMSݑ�x�3X}���l�n�$�El��j�a$eh[�ݓ�QҌ�mW�天�e�l��g�kK����R���;���0�}�B3�S�(�"=4{O�1Zj?��q��e<�&@�U��n�0��*�.���h�^b���L��7�s���������`w	��|Y�wM� �.�0����I��4����Uʣz�ne��`(��4hJ>�|.�=mA4��{���]ae�,y��O��4��.���]`�w�/���.��D!�ȭ��3�L�ǽUW��\8O4n6��G�H��?*;�1�>J�٧���!�Q������$��k���-����b�L(.��o��;�#�(<gr�g/�<��%���͏= �R��qk_�&ڌ�qZ�ە({�E�3��=�|����3��E�K{b���+�Ǝt��0#�ԋF@v5T2qn,x���6��v�q�(p����
��N����=�z����H]��?I8Ľ��JFn'1���֜��i����]<�^qg��䅉�Yd�H#��	L1�HV�I�n]���U�٦	�֢E�u���Z�j�[���J���n}Ʊx��$����v�5Õ1=o"�y2�^s�U�v̊�n)jzv��J�z�Q$4r۫���Zt)2G;�t�����cB�E�e�a��$�Ծ1`��ʣt2�� U��W+�^�!�p��GŹ�s����߼�R�B%��VCN޿�db1����H6����c�Z��I������VVl��q�L�����3*X�	5�є�h�v�&/�������U�㙳4p�ȝ�ߣ��Χ^Eѡ��9��mJ�p��:ui��]���b�� ׭VNaL_��칷�=����EȪY{T�>��b�	(�\���|s�NJ�K�U����MЋꦊ��#�6�4��G��G--��X��!o�j�"��62i��c�p�:�A5���6��� 貵�ڌ�7|�)q��X"��&5P�;�^��Q�뉯�Iå:���G`�5&�9����	���E7-x���m���݌����Y�E?�J�惟P ²ly\�"���ۦ_*��<lS[�D�7��t�,�𡍊;��?��<Ӟqe�͔#}�o ��_�_LT�z0��e!ObrM:��	����v��Rd�G��|v�V-^��7�R�V
+�ݚ8kV�c����������t�fsM89�J�g7s�c��4��v�7m)�[�&��HÔ��;��g%�Y��;M��s�dU�"-JݐQ��ͿT��j�c�Xʗ^'�c�����`����HZ��ݨBO!L6�ƛ���	�~@&�
�Q�%�E����lӀ+Cתl(~ƅ̵�����T�]��do�����H�~�	HQɱV�֛�ҁJ �d����O.1Đ����̥O�����O�U���N��%M)����V^[�"{�n3��z)��D��@�}/�w��Q$�?�V*��6�g7@��g*~���<Ts�yB&���ʶj��ǌ~ж�FDqd�~wA���)n�%_�����Ӯƍ@��C�	�뎖��.�z-�r@��#�$!�9�W o�������F�`Yړ�9�v�@�_�rvgoR�}�K-��3L�G���;sv�a�J�h\8�b�	M�$`Q��5h({��cK]^t3pu�w���p2���m��~� ��u���=���X>�q	�T�D�Nea�-x����V�Z�� �k݉?"<�l���p��N^���Y�_W������j���=�ըO|5�Ō��<��A� ����B�Ԃ{w���-� ��-4+��΅u��<�n'��M`�\�X�M�(����7ޱ�J&Z,�+�t,;SE��kྴ��#�*�۲�y���Uw�Y�TQ����^�� 1}ᡫbn����ɟ�B����ex�ovak�|�D�BQ��b�g�*;�bv[gWA 5�Z��{�R��&^A ���K3ΠzI}�j���U��-G)^Q��5�6�maI-S� a����p6Kg��i+IPOMG/~!csF�o�E�%}�U�Ļd��K�6�x�V���g�֩�'�J�<*����7��zi0�F�lx��C�`cI���̨��J���8| S�w���}O�>��u�:!X�B� �&$:e�7 !;�������n�0V=<]�G�&b��^A���#eŪA4�o��]+��0�r`���1dhpI��ӣ-�/,�/�}V�ʛ����E�S8٘�����e����o�^��7%�n�R�����x,��3���D�OO��o���]3R�L��p�iüp����ŝ#N=�!3�7q��"��UzM���À�_����?�u���y>�T���(�_�BK9�Ӫ㏛5O�A��R����$n4�"�"�	g䵔){�wH:S䩵 �����KE����ާ�j��b!}�=�h�������MӲɒ�*����.�C�ڍL�q��K�-��_�'=B;�0���1�`l��&z=�T���W
 �k]��#�T�t����e����0m���!�t��c�mI�ʪ��1NaEO�!,��b�n5�N+�~x!!c�\�hkx��V7}�e�!����Y-=?D�Qjf������è�+C�پ�a'+�P��v�!�����yc��_���Xy5~��Ʃ\�g+M��G��Z�9{�g��^��>M��m��ݎA:AEַ���:/_�/k��=��Z� �i�&�%j
INs3l���@l�}>�i�/�1Bٯ1�o@��!rc�2�q��m��	�w���?ϴ��ة=��z�>C���t�F�oO'��pts9�r5�8L�{�e&j\�!ϴ<��]�O3
�Á�R�f�P��^B[9��-�M�j��_N%B#F��	��_�2ӠM���Ҿnu˓n�/���xqSM�qB��
t�����cw!O���������z]u�$�se���^��+p��=��lJ�]c����_�|���>�Qx8��=�\�G��qb/}�=�
:5X�>�� 2tk�שET�=�T����òP����\ 5�2�#9��>�N�5Fu*{R��,M��Pgx(����\x��;��>���:�`�����=��q́R��Jv8�(�.�\���쏍�d�ol�#�jܔ<��[N�O���'������gWsCjd�F���^�+�e�KFv�tWN/�#q�Fv���He�\v���E6��g�
u��,�f� �����ד~��������vZem�	���$�Ӽ�B��ڔ̨9%�������;���c�� �����I|�}�Z�=�_���1LZ�d��{��u��k"X�"�h$
#�G��.�'�&���-MU��5 �#S���$RyJf�x'�#s((���ܥ
j�����j���&f{��-��-E��s�I��&? ��L	��ۿ�1�@�c��B���k$Ѥמ!�L$�pf��P��Fs�= ����{r��z�\�3�{*�*g�4������^�[������s�����2aw[�C"f(!��4[{ѐ�����+I�A�'�����$���&\D�l��|�&��ς��ӎz�p`ܱ��a��X�?�L���?��b�n�?������ɐ>����|56H��E,��/���g���Á���`��T���I@q�TR�\B� �x��^?�Z5��2�Q{�4��j�ߜ2�g|�a���J"!D�)s����I\L��!�dj���B��Z���r�8x�ўf�26xU)&�I]̑�R�u=JTa�ʯSw�D1]H���o1���$��Y����#��`�Ly���!��Gm!�&5�/���ۜ��P`�J0A�!�Tt~���$��"4F�
�uE�V��*�sѡ;?j6�U9�%���Z��U�X~�M���2{����C��������`�����V�j��ݭ����]���^j�8�Ǯ�xud�q0~��o�]�D�+V���3֎��Z�ɦK���+H&���^6�rj�y����c V�.�jP���[9��R�r��ut~���3�ͧ��)��;�Қ�j
.�B�kkl��������Dy�L�M�ީV�c�#4�D��[�x���^s�n��7yB�uT��xK���ȏ�=�5w�J���ibV�>�FZ��`�Z�������pFCC�Α��ڙ�9�)h��1Ӆ�p��o����坄�c�;����>��G���Z~G��|�;�0��@��&�_\���^`J
���75�*��E�����BN੆eޞ�e�ڪ��*PU�F�/��~	�5`���uy������g�aN�(=󽠶�����-���K��%ZlU�~BkӴ?��������,Q�?X@ķO-!��a����2�D�\MtS���U�_=�tR@F �Ċg]�}���_j����ko�7MY=���5I�7���@��% Y8ẗs�f|�],5�'�ͥ�u��D��K^N`;�mP�=�f/�y�x���XlN��H6��ի��
+KƑ;�ۼƞ�����|N';ThVwaI>�������ɡ^Д4w���Tu�\�L�Qd����(�(��˱����/!��ۘ�[��O��b���=s�4���v�qڱ��)v0�!t�u&a��݄۷������Ts��N�F!��؊��ųBҝ};�x��7ɕUډQ2^U�r�)�ὶ�-C��?,�z��0]2�.����]�13@�uS�=1�.�����. A���)13K�5�_�l�Pkiݒ�/>u&��^��_]1��Ĳ.�qF�o�;����LG]L׬�w3���½<+�ھ.�KZ<��^�[xh@��?��R�p:���EX����9 ����~/������y�8^	;zr''
�Al��^0	�;�8�W^�peɽ�i��P��� �B�,^��<�˱$E���ky�=hೃJ�O�L;�>"���`�U�)�y���z?"d�+�
5�k�6�"	P5���[�#���
�0֍sm���3L��ʺ+^T��,`����(#Af��K'>�a|M���m��w���nR�j���-� ����(��Y]�3�'��t�n0���o~"�c�z�v��~��p�8�eA<�#�D����&�rҚ��
���h�e��ʯ�o���^`K�&�1B����8h�/<���}������~�e֫�[۞�Lw0{�z�:)��?��>���lӷe��=�$�3]*y�9
C������+�_O�y�M���E4�)L4m��sـ�J/��]O�MnP�ݮW@�[�1+r������0y	2</4����~�D�?A��ۏep�Dn�۹��d���X�AP�چؒ���`än;<U��� G�y�EX�^M��Ԭ���<kD��@C��o�1v���z��L�bmw"���}��	�L�G��6A��SAq͞?�%�+Y �I�o��ntu؆z�2��S;Jx�?������C���6)ȓ�Yu�-I�wy�Wx��Z�eCR����>+�{�B�#��iB/��6Jn`ܙP�7&�I��[�#�|#��
Z*�@i-n����xG�i��v�3K<�p��l�V��6�Cؠq��K�(�cZ�vo�f/�aڴTu�-n)PGJ�w��OSI>�"�&����.��*��>_L~*a�;M"v]�-F-��x���5�.�;�L�U��c�X��k��f��7:�=�p6�NE�p#�Z��3�\������`��ù�������(Yb�\qP2u�;C���ڛ�I$�u����۬�tqƿŵ��I�Oc��x?��hLc8!�&�e��g�-��.�򭓍[{�������B�� �/A{y�B�o��Dv0�Yɜ��%k~�۵����=�'[���,i�9Y�����E/����~j�+����R��T�o@�]����QL�H�7�2"�]?�+⯺sn!��v�oăjf����e������:��Y�߷O1/�i����ƲQ� |���/����5xG��$_��Dڏ/�KX��`�gX����ӏ������;����?����IT-GvC�\��Ҍp��5��/�8D��DO�`�T^Tlη��@�!Щ�07A,��V��.V��vSXը��Έ��e�����U��_�tЃu���u'�H(����*?�*�3k��Q�v�] ><Y�Fo.a�ʱ��*�W�J��.��V��<ԉ�
)5Z��m@��	���;�\��Bk���$&���4���b�\z	JKO-rh�&(����E�������L)�j�nU�H|�<�r�� ̋^�?3�A�=�/mt �+[5�W;��~���Q�����,��k�J�������{�3��O�����m��`��s߸0�lFwQ@y��&��(��M��Qا�`>}[�G�!�:_�?A���@�E�Bz��W a���~�I��k��ɦ�LmL���qóbp".�	�DQ�܄5D,/��3�T�r����V�`��լ������HUQ������L�l	A��ᷣ��|��[j�6h����b&0��<M��O0�fO�,2=r*u�;j�O��i�y��������+�z[�wnf�W�f&Y�.�9�)�k#���;����'�S�҅�@�5`<6��>�o���м���<��L&��PR|���H�ѫ;J�6ז� E���$M���b���jC&y$�>�OS����G��>IC�sׂ�\H0�/(���1(��#N�;z .#��;N��(�!m��˒� ���s&�= ��p�?����v�+kp�a�g������������	�6dg6V8��B]"7�#L2��n�vF�5|b��W�6��m�_����j鳌��8Q>�|82`7:��q��T�_�0oR"��~��=E�@t��`(j�X@��hΓ����x��1�ȋ$�̕s<�o�r��w�I��d��0��"�^��k�N���P8�H2�CF��nU�+Ǝhyܗ��3`�xk���9W�Q<���1]����LಳF�69K�dJ�O�V
�	�E�Q�D?M�c�9�4��ͦ~p�6�u훒ʆ=��t������o,�z�����WE�_��+�#ݲΜ��5
���_�;��QéŎ:��!�g~fˡhÞ(F·VS=�?C����2�	^��$S���i"'�*k�J����
�L w����Ib!�d.H=Tȃ���.�.��~���6<��q_M.�}*�꼗r����w�;�v��e�[����t�o�F�Y�^�k�=���m����~}y0���>�q��ljp�TD;|P�Ӗ��c�z��������jf���o`=^���fڨ���8��MHB���
��^k5R%����E���ف�u��l�F�؇��b�>�����Y�,���6��7d�w~��;���(�����l"
�)&���?`�7��Ǟ��a�$����qX70&�]�v�<�)�͋�_�>�J`E�Ԗ���Oi��%�3���&k��[�T�
��^�������pY5����D�^��������^i�J/�Dq@R���y�����bD�����*ZA���W ž|�_�u��pό��ˊ�b� 8)�nv>by0�
S��8���7�bL.]Ƽ�7'U���I�����dK�o����$�|���)��J�k�����R��:l�@�|�&4�B�Οv� �
e8ݛ���}
��)��w���B��T�p���0,6E�+@ϯ���/�����V�#m�70���ݼRv6YPi�г֐J�Q�Rzܰ��ϩ�{��ԙOAmv�j�-z����<0�RQ�B�p3O+��P%���50T@~��/|QËC�$���9h�Z_����Wa�~6pLW/S��I��m��;���c��c���Iu�K��p���
��PjEn�y�n���k��_:8�لo_�����xY��1SFX �`��	�����z�F.���W� �;���#�L���h�;G�xWq9
�P��� ���,ð�H֚�W\���*Ҭ]�� ��~ �k�gl��L8б/�S�z.)�� ��3��3��c/P�%J[����8I�B],���+�`i��C�Z�8��.̳�z��oXc���*j�G*ی���(v�W�
 �L��p5�.��V��`���e06���VY>d�X}+�`�)������#���q��ʞ�l�D Q���E�ӑ�p�+�c`��g��x8D��p|">���^��X4ҝ���ߡ����X�J{EY�1�S�w�
�'w[EI��w�Mֽ65+��u�HZ0�˚��q[�>yQ2���@�挊�-QO���O9�;��:�@�ýd�ǊNJ������Ѧ+3��{��.|}����-�w�]7M�q����N�����C���Zfˠ����K��`"����r�iy9��oh�8�N�h&��-j�{!}5�,g> b}_��04l"
��H/e�
�PQe.�U�N?<�۵:����7X����>�X.�LO|)�!#� .~Q���r�Y$�ĵ�:-�&�]��7` �����Dć�0��َ�냉ߨʱ��Q�$�B��;i#�a��#&ɑ�0̞U�';#]EF_�@�ᤖx��{\(_{��4V��x�B�Q�q��y��z�2�\��-d��aDO�>�2�n2��n\!�ǌ�j��.�lq�)t�<��L��~}�[�hJ�=��уBN�,ǲu�&']Cۼ"e��TQ�䭻;x��)CM�J"��|�J�e��+��x�4�i����Ü��>�0�ʟ��
�Z�o����Ѽ �U�e!(۫N� _�'��Q17�Ȍ�]mP�vLF,� �&���'������m!���g�=!��?CO�hi����eA��#�
�X��2I��m�P�~�GBz
�����A]�@T��S#3G��j� ��՗π��X��<��1�0&&pE��@��u��I��C�M/9q�P �r�ɼŭX�����;�RL�I|b�~��G_�yp��*t0���/����p5�{�{ �)m0xY��t�@$�+�d>�q��-��+�����i�GC�bv6%D\�������]���ܜ�Vc���U�
���^<��� l�*:.�W+������D,��_$�9`��M7!���KȾ��֦��[�ô�P{H퀔mu:�+��^ /�w+\�^����=�����o�+��Z6��p��?;��|�RA�D�6��!.��ie����XP2�EtQ�\ ���r��`;�Q�#�	`䀨�f���݂�=J��o@M����J�`���3���4r�a1�J��S�����L�l�{��NT�g�0��}�Io{���|f�y�_�A0�q��Y�炜tO2�ЮZ|�����p.E9�A�{�1��0D{�C�X:�+}�s'��H�F�6�K�@��U���ḡ����U-ܾ�>�F�?O#mfb=�Z�P��d���W�h����k$@!K������͐�i��P�� ��{9���.�z�f��twQm�Q=�����x��7�С�`A�F�e� �����d\]ݪCf��t�k+���c2�S8�ӾJ*�蚾��5��<F]��Z"��+1��o+�<�~�{��[�~)#Vn[*s��eR��#��3"���o+;m�9w���a�.����
�v�
�b��b@B�T��.t'�aP�A�s�/Ķ#I��Ŏ��é���״L�sM�n�����ɲq�)�X#S:�Y�*�5Eqݲ)ި�@:E�.������G|�����%B!ԫ�=Vc1�\$vTxM�u�mQ�^���Ӡ�[5��
;^Ȩ�u�	�r��*$#*K��J���!N�PlO�D)K'���ǯ�Ȑn.�a͓pm�!2X��e�@��M�u���4T͋9)��٬`�3�d�;��O���XT-]XB"�=�I #�&�Gy�X�Uu��~=~�7ԩ��?� ��蹏�h� =����;�9Bܴ�������h���{������B��#�\�gSd�h#�X�5 ����?$�:S�fP��g2/��䘫���Mђ2����/B5�wƁ������_���-�cB<���p���1D��q1��M�.��lq�K<��L�A{C5��ֱD3���� �0�M�?qK_�qg�����Yb���w���)�U���'���4��Q�Sd���z؇n��u"Dg�,B���2ʠ몦��u���&?���Fi/g�-�Nz�Ӯ�_�!cr��͒��z�T֋ Nņ���4��8*0=I���v��}L�����	8}�j�[�WQ��)Kk@�Y!����)3n���wS�|r������V���C^|MC� ��c=�$V$�}���F<�� �~�.Щ9�0�Co@�.�J��?V�q�\+4΢7mX�=�t��L���
E����S��.�c��-/�ˮ1P��,�֛v0�İf'��4�]��Jk�!�hˉ�3����3��~����~7��d�I�R�Q��>P�~�<{�z�x0}��A�]k�J�g�P�ՙA��.�L�a��[r��t�T*�s�`�Qp�n\�tO���]��c�w�zݷ���A���g3�P�}�����[�&�����I �~2��f�}�t,��e]ߐ�����c?��C8�'CwTf��_3���eLA��P��I�R934Y��~��������8�E�K�[�h�st|�A^�����1�7��яmȶ�z2��6��~#1q���X���g��U�g�3�0$�s�X�:u�+/@%�����[�4'/:ғ�?meP�+Rm{���2�� T�N׉����u�J���=Է!�9��Y��7�|'��O��U�f��	��1GyAK�(�v���@ψ�	@�I`���!�kr���A�;e~�x�Q�� ]��1L��r���~Jr`��S��Y1cO
K�s�!��R 
�N+&�W�-N� �9R��s�U2Q��U��R�\��7��;�H��q��{l�t�������h��&r�� ���W�b��Pךs�P�Έ��FA;���(���!��F�|�������' �k�sSQ��B4��H�o���m��I�xҪ+�pu��8E�d�+G������xu ��β=5B�}�I��h����J-k����\���j�n�6e-�Lس�LJ|:h�Ȏt+��x���N��H5�������k|��ɷ�K�h��MG��7A1 #M?T;���8<pC�����	:r:a�Yd�ɬk�
�Jk�oХ���M�_ͧ��O��g�_��a��!b�~��H�/[{�h"��Z(�*�q���a�􄰔 �*��+1,���u����lJy���ŗ��B���:h'FV�d
��J{���\c����$�AˌJO�m�8��x�5&���J>#^z�>�,�W�����F.&4M�#H-�k�;%�7����09���WW�����S!�ᘇ���!���3����
��{�r�vc����M���&�@ڼ��>]�e��0EWV팶@')+�)��kq�F>�;���.����Z'c�#�ʀD�w��j�h�f�*�)Agˬ��qA~���h��H��s��+���l($��K�܃J*Osl����#�ZF�?�¦.q��-�W%FD���B��
XsI1�h�?G��ɥ�$lg�֮�1j4NR�(�:�24�R$&�;cB|�����)-x�e7uR��I� �Ɨ �J=���6l�XwG�D�=�3�8�o�
�����C���R�l`���@Q�[����%Չb�M��n��˟�g�� a�MM�t�rM@v�q3%�殤?K�Y�\
m�~�Ӭ�fG��Өx�������Bw��*R���~�b{>�������ϖ}i��M^���Z�O���7�B�1�/3O���Ro�����®�
W�2P���	��aZ�v�LC������2Ur5�D7�p�$��C����SjAE
(�G��|��>,rV�N��<�r%M�Q,��3�=��`�N�4�:f��& ��M]��� �j���)�!wb�IhG����E���ښ5&��iǊ�x�
w��K�~��g�B��<u��}����p�,��(�{4���J�%{�d�b���1�n6���k�<��r�8(-�8.N��dT�T��e�'n�x�'I�*Uj[��K
ֵ�_<�^�Đ��t'8�N��#�+^�܏�.�����x��~ ���ݼ�S'�tg�4t�� �%h������X��@9�FL���d���%9r�5�<�q�����D5~���hB�� �ݱ���I�H�b^y#���Z� ^�@Fn�.^*�by)��Aw>_��mS!��$ƾ�q�Od�sD����b����3�����i�se��8eM��;�,o!c��T�qu�A�*!�i	���:�*���>��f��/��o���2����\�7���6)Z�����rǙ�J�w�J�5v~Fi�"���Z��K�._��!>I����e�h0B�(���H�)�].�9K�28�����։p�`[��z���>�*4ai�Y�t����=�P��6�?�K�l�zmd��׼<)7���G�,r.�2�is��[�F�G��!�����V|�+ԋ����϶k�n���W��R��5�׬;W�劥k��\�i0��/	�N�.��Y)�.n[)�sή��������x*H-r��%w��|�8����I˄⚙��>���0�����W 3��';��b���"�4�˟�V�Δ��`}M\A���fH��boqi�juo�1�J�bk�o}vgB�w���5��N�u�}>�B(�u}�t��=�iN��tZn���d���ywHl)��h@b���"�� ����h ����4�������ۂQ6�<�u�-�s�p�� 'yQw��X�7�	�S��f�:�Ң*(Ϝ���^W%_|�]g���Ŀ��NRB�@s%�X�U��FX3 bA�}���;{���+��v��J�&����Gtn�a�.榍#��Or�*��g3�e�"��U ��羣�sd�"�%]1���M�9 �Xq����lC�},�.�P�
��|Mf?��}�uΞ������1zĞ���4@�q��D�;��R�^�U�b8
�����A�*�q�W�+�9q*VC[��f3K&ċ���Vu~uhT�K�P�o|�'��[������ȟ��Li��0C�����BQ�L�Q���M�����Dn B��w ��ݙ�ݏ���&x��b��' � =y	���"�)F�����.�� �r0_�V:���񉫔k�g\J�s��+V_R	z�&I���zUҼ]:�QV����{���w�I%쮺v�{b�H�6l���Z�,�����C�dF:nѸ9�F�E+�(D�%\�l��i�34�X=:�F� �C����n���k�?���7�����B�\a�%K$Ul���I�m�ˡD�]�sT�Xvo���Ys!�8{b�uND���'��Җn��0p�k�`�%%,4	�K�'���=ο��,� .��tJ��_�ȸ�,�V-�G�t
���& �Ԟ��zF�ʵ��0!4�-��O65��.�d���HZ�+��Wy������AސM�o���'�es����$E��=c2�>��Г8��S&�1����U W���ٽ_,f)W�-pO_+�"�1rq��xEg�>�o���ٸ�����B���~u6�=wu���=˟ڟ(�z4FB�m_�2�ꫛ&?W��O�=,d����/f��z�L0�S����ѕ�m���uU(o�r�G;��=�=�[����10����8g��,��(P��p��f��?�0J� �^u��X���c�a�����+}��6z�`��s�,�b:���M�v+���½p>�O�O���t����NV�rn)W�wk����z�ϐp7cΤͻ��:��a�����k�J.����1eK�$��#��HA��?���c�з�l��=
`��u�U ��N���� ��h5K
�&q�R	�4�!N��q9$ti*���*���)���V��
z!�X1�h�\jvx��DOu��E�z�,�������x�a]��Y���w*]b3ƪ{:�����L<�m�ZM�rW��.ƞ�Mnd�,.�J��&ߑ�L��w,�!�@L.\֝{�y��T�iQ����$^0EHn�e@� ���V���;�:��Ƣ�(�jg��:����9� 2��M����V��� �H�e`~n�/��a|`l��zRcYa��vf���~�c{%��x�W�Cy�m ��1_�,�q�5�Dw�H�=�j�aᚘq�]� C��7�eǎX�[E&֦�
��Ùe5���ĤR6��� Z�3����7��Y4�37��� ��m�z��QdA������ǳ �`�!�яF�t��1��OA��I��/�屮�)x:�zB�~�]ze��9E��%�W��������]☜i�O�܂��F���Fsԝ��h�����{;�<	�T�����~�����%����A��i��sg)�b?C"+�=�v���g`6�������,�Ī!�U�n��3�2�i��Ӄ6 8�4�0�4�ܘ�u+�E�~&_�f�o$��k�cb[��4U
,1.��/��MK6(Tr��us�R$d� ��f�@�����E����T>�̑M����ll�s�gu�D
"K��K�g>.�����/b�v7cnjq����5�_Z�yI���Ǣ��a΂鉉�D��cUC>�`�1�9|����B� o	%e����#�b`� x���M���a��Ț�2[��)�%Ǹ�@�X�5�m�15����L�Z
����a�T8Q��\��֣f�]��^���M�u��aJ�\䟲*$�!��73V�a��Ȭ���p1��
����Ƶ���\;�y�	5[�O��u4���˨�Bo�����'4ls�������񠯙��b���,�-��U��H�۷H�.!ua�<�WPG���/�ܵ"�Z ���U�6�Gs���}�)u��a���c�]���A��X��H�����ŷ��f�7=:���r�݇H���a��¸���[�&�JqJD�ħ����ӥ�f�-Z��'&ùk[�.i��s�>����t򴿟x�}�1t����hX��q*]��׉&Bľ:�Zj�zi�J`!��{V}�u��I��<|Z��/��I
�W��g:�(�����p�^�������q������7�U���X�XA�E���|��P���u�`R�a� "L<��-��%:�(���DF�3�\��(KNCpceЖ��6xEq� �|@A��u��q`�'Y�?�u�̋�t;w�P�b* E'�'�bE��_�������1��r�ͮ�kU�|����8�-�KU����\�hC֋�2�]�p�q�zZ�,�&�ƞ����mj�r���I����u��Mf{�S���I>aJQ�N����|~�u�E�k^5"��]4נ�d�#?���}�_�[���eH 
Y�YB�Ϳ����L^���?���\�s<36�p[�:k���6]s��f��Ofd�
0,�r2��@�׺�J�uv��$��+����U�M��m͝ƫ���	�J�[m��qj��|��Gj���	�bC��6���@�,	��dǁ`�d�
LN�Ĭ���W��,x�H5�ؓ�
�IDɵ#��)#r�Y)���(������;�%��:C﻽��������0V��ڼh9���d�_&�ͨ2�?<��}�$�;��P`k�$��k�3K�x�4��~���T�2���+)Fk�Wc��S3V�Td���1�i�������'�Y�AH9qq�h�{�U�X!��zӧ�H���!H5"��4̀�U��� �1��_R�RC�K��@�1a�F��5��%��:��b�s;{S��EP36	.��49 �XYn�FO�m�I4��A��͙'&$�z�zj��p�+�lPx��m$R�%��O'K?�3�bO\���a��2t�k$Z%�Ý��d�N����wH�qͿ��(Pn&J���u���X� �W�����Uk}�f?�&�^ב��#�VY�}.$UXj憥�9�n����&2�"U5^����G����@�|�������?A�����/�%e���ɖ��q`�x���m7���4d*E�ӜrF�ݜ���k�wOΡ1o��dݝ�َ�D/��}�>���ꙣB�@�z���Ł=�|99��G&��e��Y��o��������e���M�g#Yi3��$>���Zo���ʻ�wI��v~V����^0�@i}��12��Q�l���wd! �L�rTl�M#��%�'��a� �}z+���$�ȷռH%[�;�� �>NDl���h�O�������N\�L��pc⧅���y���
�ʇ+fG�=0�V-3��订���H�fxhFީq�܆a�ugM���G��� ����@�w�g<5F]4s9c.
��-So@n��B�lC2&/���E�Ci��v4-��z�,���Z[X�s�>Q�MR8R!,�I�ގp�k �y =:�+I,m����$��<PP$ġ�$���V7
t@^ՅC?j
��M^��V�AM�z�Ѱ�D1��LW(�(�r�RJĽ�����j��Е����%�d�rd���P��T�뉴�������@��� n�����6J�>Y���<5������a�a��ڲ?����q��k@'�^�g=/����k*��:7I$P%�e�)~BB�_l䕿�������kY\���R${���7*�&��!�{Ҩޒ�i$;�/���B��X�@�U3v�;�le���L�r�M�ғ.M$�ۛ�h!���/&
m���^�@C�k/��ɽt���qdT��I��bm�ނ��D?��6�kK!!�ng�R� �� �8wZ���lS�2[UY��o��p�8���^�mw��ӎܑ$�a�>2�c��ﴳ։�h5{�a�$��$��)܄3o�B��U��nɭ�\ gԇ�!�@�	��u����R�kV�k{� p�.���t&Z�)�w�yl��L�qr"���C����9A�Q݁�]F���-A�{�"�Aq��9V(�|��%:�ɧ?^�f�Q��ݕ�����{��h1�jA�G�=ԅ�)ƛ�rh�U.�v��:����l78`�,S:�Ʋ���̧0�A/�m�Ad%`�"�%P*/�/7DX���mNb���B�ep��|�Za$�/
�ǋ6G?�@q��S,���\��
:�+vۓ��'� ,�j�F :5)B�N��|�ڲ1(54�zۘ��t>����c�;g�n���19��^�H��)~:C�W!��.�r�bFo��W��|	���������N�őr��OeL�o��K"ޚ��e��ʁ,o�=C�lN�]��=�J���g�ņ�z��� ��!?�E��}�Q�J������d�4|b�ma�j�}���i�v[~��e'��!pƄ�\�Qe�͛ũA{�L��p��(�e8u�G�Q �`r�d ���P�rf�V��=��cp��[0F�\qU�1|ZR�0ݞ@
��ݓ?f'[���Y�&�
3nr}��d��AI���	��j���b��ՠ
F�bys���E�۸VL�����Ql�d���&ޫ�/��9�ؽ}F��Dϭ�&w�B���V-k��ґ���E���#01����҈��<���٣kiuf|ϳ���)@�r������	e6��� C���*�/��L�5a۩�i��~w�}�6�Ɠ��,��I��Y�h�DY�ׂ$��-lB�B*�H�}v�P���+�ôI��|G��aQ$��`��(��[�PȎK3f�N�	;��hʇ9�I�]u:�����3������@��b���r�"�vbbPa���.��)[j-�C�-G��YX�jv�nf�� �,0��'��N�:����v�B\���	'�m�U��q��8�Tȸ�V�U�H�,��ꤑ�ٓfAԨ���z���"�PN
�8��2�3@���f=S\v4�l2�lV�C}+%�X�Ԕ�B߲j+�у����!�Ƹ�>GkX~V+Y:�W��ʐ�{�`q�Q���<j�sw����˗��=D.Q^�Y��`^̨�3%����Wۆq�p9�?� E@�*�6��n�A�a���9��/ �Lc���Oz��[����߉��*�K��ړ80�g�f�/`J��@��V����	��q��ru� ~�Y��`:�P�a-TAe���8�[%���7���E�q����23�[V�sa�r_���qZ;A���S_�j�pY�hM����K��	N5��a-���9�{���@�����!�2���6�J�)|9_ˠ��I�3���j�qqH],kp�ӂ�q�?���kb��4&IZ��3��i���?)��2�[��j�*���Й�B�����sJ����@��>RI&�!�iy4� �
���̷�l��V�>%�1�B�v���ߊ�p��3C�,X�$�%Q�Q�ߜ~B��,%�CC�8=R�'!� �,�#Bٜ?�y��h�X/R����8����!�z�Y?�����Y/;�u�R��I�5X�wsWZ���sc	u�J�i]��5[�����z�<��Mn;&}��n��ͲdL ���Ѱ1`)~��
���ò/�]���_�z��a�C����D�P�<L@O�h�
���᷏�he{|b���K*Ȁ
�F���e
b:���Fn��mQeY��(DS^�4m���ϦĔ�ӆr3����*U{���]��z��KQ
s�Ih��%�Q�AWxQ}�r�~�����Z���vJ�<.e�1Z�C�:,�)���G���q�>�׆�;舨��A�Bo� ���������W	~�3 :�q]2Q�Y	4Y�2$���"JmcI�zNg�K<�����jDJ�.ߖ���+��h�KiE�tR���v�F�g�d��[g�Q�@��q*;�ǳ��s�ύ��qm��:��_!���9�9�[��A)�e9��t�Cԝ��	��M�ס���m+����Uw]��y���*ΨUM�� '�f��}_���k�A�u�i�c�*sv�����2Y���6�RM��?k�3bu�t���
]>���� (��:�hVq�^� V�ݳ*�hV<��(���K4Y�Zd(8Q�`��hL���c8p�7<)?������9A��Ђ��MM�k(�r��>>R{H���Z2���܃����1���~�=`�g}����K�`��8?���x�SwvE��&@(��ɕ��k�(�7�Y���6�A0��Z$�L�3E�}�!���u(<u��i��pIG,0F���ʈ�h�A ����ۂ`5�gz��-�@�.j���ȓ���l�.�jْ�+��|}1!qcГ%�v�bB8uŮڻhUmU��Q���Z�쮉���V�I��������B������|Z@�f3mɕL�8ݐ��ow��Z;�=��2[�T�~o����qP��A>��C�m?όg�+�а�h3��.�|�v.�+b3�/�c��
����ض��MN�~ǐ�CLRӣ�a��'	��*��1�}T�3IލU #خ�f�����ӻ֐5��@��.[L���Z�GM�BB/��N�p��p����ߣ��{��%4)� �,����R���di�v|��˳�DZ�g��Ѭ/0��gb:��9Vx&�����&8����q"�� �j��q�c��׆[
�bTE���gF�d�UP���<p� G����y ����o{$_\	��q������cx�&�~��/er ��I��?D
����t(?)0�U�dHδ������[r8V����a�Ҋ�O���;� �q�<mw	8����.�¹����tU;ż�qGQ�����}Z�{sCv�t�T{� �x9�F��c>�.]9w#<�m����))��=�u��%ޙ��^�(�`�k�i���������2��nS ��m
*Ѐ��>���ґ:��]�~�O���1.li�2�'0�n�����p!����?�����o��c����ǻ�T��d�Iz0�Ͽi�f%�3�SIY̵-�yb!��״g��\���8��P9�#4F£��(��n�'��l�i��yw	�	�i{����I�*��GT4~H^�i擄���zaE?a��Kg��Q�u��8�A���W�D�����ݪ��!խ��=�ε(�{����BE�#���h�|c=
+���Q������/�f;�5�����ixQ��]���P)=�񿡈�P�IjZK������'�߈ֲ=Ҡ�)EV�Bb@�KJ8�w툁cՂ&�EJ��1�����mЏ�����[ǨKG��H�������9�Q��Trt{뻓<⅔�%��wg��p�#+�S�8?u���~����Pk(X�`8��Җ'�X����4��Q�͂�Ri�*!M�Z��2���SӤ۾�����؏n]�B�="$�ߵ̽D�e2�I�ܔ�<ײR���;ڌ(a!
�Q�����ϚH5�^@d����I-c��x���1(�J�!�_>
ܯ�1+s�zJ���bH���?�J)��8�����f�]%|�[�^�f'�ŬHt�e�=��iX"!=��.�
���8��57J�"�����3�^�AjG�sCs�0 $٘��v��� ����P6Jw���:�,����������tI?���>d�B~�DՍRI�7�9�i?Tq,�M�,��2?c�=)h�"����-�l��	N~�&�i;w�xG}�{�+I���ɋ�X���!/����"��>�l�&�'6��0�(�n�O�S�@�
�����W)��Y���*��,���@'Jr���z
�1�u~��"�HYH�M�O%EWx�G�J� NZ��h���dɦ���F?�x;��+���i>��� ��E����o ��z�7�N��ڜ��I/f�Ȱ�E��� 	#.t����l�u(�b⚨a4�Ԅ��3?C����Wf�����0h�耾���F�w���*�O�xY��vZy�:ky�m���-��
P�Ft&��@/��4|�g(s�&5/p��G��=�!�_���R=��<�ۇ�U�(���2	�b����w!v�}�� [���	���Q��rʗ�왷��e[mK���@r��<���O�gԭ�;9#-<;^�,/o^�k�X���W�7��[�<d���T���]�Z��"r�!�U���_�U���Y�I���
۲��	&�r�A�%2I�a��^b\�ԇ�ɖ�kP�W��� r�����VS�nd۾e3SC ����( Z,w����F�P,�/��z)8���Xn]�і�(n�e�����������L������NZAΊ����Wi��`q��t���TI�3t���6��6g؊E� q5�.� ��HfY{�Dߥ0b���~�\ q�a�\?�X�x���g���J��U	�8c4����R,g�l�2n����#&�G���N���,-��@*v�)���f�Wt�m@�\��z(t�|v��--)���D�0��`��ũa���D�H����>m����S��u��	�`���S���♕Zށ���k�Y����|̮2�j�y~�ٸ�k��������)Z2�D�����P^-sľ�#���(��D(=3�C�o�K+�#|��;n�����<?f���g�F���7Ǝ(�Ɣ�#�_��Q���]q������JE�O���8cg�P%��D���e\)�o�# 0�$�Y�b���9�`v�f��s X�ږ��'���v#]{�_�� 2��I{�j��{�)WA�Ms;1�ɨ�g�tX��44~;�(��%_��Xӈ�^��RQ}�v"J)s�K�[������@�׫rl�[RWP�`���B3�J]���	��Hh�f{ۭ(V����:�7eú�܍$2rȿ��j���1Mʿ�e����q����]ϻlXN=C�[�ºi��l�>�y�g���"�z��}�>��"Չ�4�(��G-� ��V��!�[p��%�h_���S���ֆt��ϙx-��翡X�bkS��O⛂P���]�e
M����ʧ4�az�W6١.~xa_��VpV��|]����5%���щ�YD�%#��QDΥ��y��$מ&��0�a�ff�$�	e*$Ӯ�- ���\�Mb�`u7&�������(kS#��5�0+��xn,�n��_~1ˢ��Rn�����9�5�##���}�^ТoF ���g��(Z�.[>�t�#��/D����
3�}�!ޟ9�^[!�;A�1���s0��Z��9^(^�+�"��� �<B�\<�ZȦݗ>�0x��u^��a��� ��{��D�.Ob^L�+���tuw���!����_�U�(��M��tҸꦬ�h��[N��~��3�dL>e���%C�l���7��*��H9�A���q�R�)`��#|� ��>���r�rjr�D���<<jn!T7kv�0z=~��"r��4aS?���T�����s`��ZZ�n���h��\���<3� �O�(f1���@7����V�i�Ӕw�g{�;2!v�rFs�3���<��x.���\�Qګ����+��9h��xd�#��߯1���hj�^ �c��l�''�l���T��#[/�*T�3-�Jm{7K�Б�y����`Z�mN�i�?'&�Q#�)@�l}:��n��$TU����J(Mx�n���X�|�g�*���x�F��M���Q�!]��7CTP_� Xƨ܂�E��v=y�JF/�k k�s��b����sl�_�U��b3L�w�d�'a �w�i߇�N���
[�@���d�Zi�;a"6ץȾ��F���@��s_��ݮ����%���P����d���7Ύ���E�F0�� �͹JW��g:�X:D�R��߃����AH��I��;+]�����w��*�a��gL//ة���rWTDQo�)��˯<Z��=V�4Yo������D��G��]�J4,���D/_�U#��rj8���'_�H�3��T�1[�LQ�l�$MX$����	�

��M��ӿvJ(�e�� �'K:>aF�ScM�d��d�m2;?)+C�� !ܓ��;�?Q,=U�����/"���V�s���c���l�>fDk�{�f���l�WX1�J��}]+���7�=S�39�Y��G��:e��^�'���>vI��n�Az���OqEu�g<�^Q���9�yJ���m�`��I�ӥ���p��i�[�!��IR=�2!WВO��]�IGD�1 �v��{���^~��m�X�8�d]@�R���Z%�л�[�{r��ւ#h�z��9e�qA>
.OC��y��U�{�X��;��^2v�>:%��G�~]�<�!��a�U��^Nȱ�:#_��Xc�.�Z~h3�&;��'��x����̈́f�`��ݸ�@��]��ךKo�#~��	�D!�SJ�J�� fr������}�~���n$�&��2��!i�-����{_�|=$pm�E�o����uJ�O,��ro0�AW�_0Ě�+�����$YK������Fɪ����ԩ��?�f��մ��9��^��Ĉ��"v�[��m��Θ�QG'�\�a�
=	]R�Z�m�T���^��j ��M�����u!|3��MM��Air�A�|X��"����; 5?�	:#cl\I�%l}���$��Cf����i�	������ѭli9�e���}/GO�L���'74r�w,2V�@7t���#�(��_�Sj�\�-�j�i���_�C�˴Ɇ#���������̂�Ǽ�����h��l��n�����*{�F]<h�zJd����;���W�V@.��Ťt�����5�à�y�'���B�`�h��Q�)�(h?���|�m���$A�G����`q\'[��M��D���|��q���u��qh,Ⅸ�O��Xw�κ��7��Un �K�v�Cf��lBH�e�a���y,���4ڢ�/������;)��SU���m���qe�����)G���a+p}|����>ffp8 ��r�����Ђ\ؿ �H�f�t�_�&��-�lq��:3\�mi���p�yE��۳����B�8$�A�t2���/X��K]��MJ/b v6�Sa(�h�i�ݺ�7�w�T�y0�10��a�K�7^3̓A�+e��
7ܨ�N@i&)��@���`�c����嵽A����zUܐwByRC�ǉ�#���ŉ��Ӈ�22�D�Zq�zi_�)���" �ͳ�;�
�	5C�g-��!��ܫT��4�Kb�S��b�,_�v���v���}��8���WI]E�V�C(�m�|
q�ĵ �_�˃����S+�#=։$�?x�\`~�8�Ń�wA�C��|�ö��ۂ��Eț�Pck��T���۬�*�2�d`�e���I�#n��KU�?PP}�>,H���^T0�q��+h:ŸJ�&Q
�}ɸP}/������ɯLo��͆�Ơ-�y��:l�΃���n�1�e�_�j���*Fh˺��2�J��a�f�B����	N\a�,�.A'$�MF�0N�)�U��م̈́]ش ѐ��q0��į,���X�UD����[�ٽ�Mڲ+u� �n`���ڬq$���%�/�Ne������پ����f!ɴtͿl��̲l&Y�v���
����gZ���-���̾���N���~|j�Z��?#a��c��b�h�i�fUF��R\�=�o"�,�[�5l��|	�/�壅��\��Ќ��ؓ�"�9�oQ�7/��n��S������[p��}?! l��҂z�03�m|�~��C߄|`���@ӏȤ���C�N��P�˩�cs�:��%�������2!��{���*g���d�/���&T�A%����2	%���l��w�����7(Q�D��t�Z�&\T\�K8�k%�2��Q��������O���.ܵ���H{�Xs3c��6�j'��vR���5d����T��(D��{g�b����Xn�����ПǢ�^ap�g�Mz���P۴}� ��Q�B>B���s!G/�9Վ�F-�|����-�6��/LxY��a��;�b_0����GlR���i��]0	����{xp��]9������ϊؠ���btv���!�E���x�ix��#yӥ�J��,�1(�9b3_�"^�Jq���I���T��X�Ψ"�7E"o��
Pd��s@�7Б�f@a���M�]����1�,0��_�-[
�����qjކ�vz2H�&ş��Zq��4�s��G&�@��4I�Qgnr���/t�4�-6|�d����,lT���9�����f��/�[f}�]�H�#���"(����K��6���e�6�oxkC,�NA��U\ �����6�����5�_+˝n�� G�������C���
�x���Z���_3�9ڙV�)$����r,��
�r<��5�V�LwP�|�q���1�#�e^h�W*�.�r���� ���pz�
�Vp��BN}�t��_�ٱ���/��jgא�J�T����:G��4��jE��ꀭs�5�_rȷ���#�R�	����7ػ�t�w��=��s�#6A�@ăl��w2=���v�s8�X�����BbnbG1� ::����pdky���k�gI�@`���~#�}lu�\6�ʵ��!-�Ь�YF��mqk��dy3�h�=�2��
{NIO�P\�O�H[�\�l ��:0rw0��Uƾ�!`��/���_~2���Ĥ|���+��9:��ːM7"���B�2�,�D�i��g�{�?��Ӕ,hYL�N�3G1q.�׆����u>��7�~u�4��/�W#x�,�4�q�F�ԥ��+ A9"�-�-����$1ܑ����� [|*�%����-��d^<ұsJ����km(bRG�D�C]��p.�^���e����-��R��.S�U�,��p8̄�����Ȁ�&���L�S�s
�$��fZ:�|�`�LG�P�GQm�pʫǗ��R�@��≌��Ǉ�/*z1�jFO��%s7����.߼�,ms-9.����lUv�*H�� �#��L�e�s�������|�ֺ���n/Q���k1��X`�=��\�A�I���m��&U�F�R����_J��[��#,I�o2Wg�+�]�B����r`�4�������o��R�����A����k)؉�n��f,�[v���pa���nx�4.x�l��w�a�b�	r�C�]]���}��I����WBs�q���2����>��6g%S�Y1D8��-���xH�;���%���l��i�-ZQ0Ǆ>�T���j-`��K�"C2��%�����E�K�h}�s{v�W_K9�����xo{��#G}	�f�@�l��d��.��nD:�}�`w8�9h��s��⹎��
!G�0K�_/�a��-u�;��=�Ŭ�XS���V\p���K\{���V�i-�3#�`�C�[M#����J� �X��pt8]����!��5S�5�v��Ģ���b�P�F�,J�>-�	��ɘ	D\}������E8ln��'q�zp��yL��f�Lم��3r8��B�=!��k����i����%����������1b�%ޖI���y�eJ����F�߹�O���U�熋C 5��Cu�p}]��r�7CV��V�H�ўیm@�#A}3��i�߳/?�p�0�:k㱣@��}�J����Jvk�!qǭ�δYQ��Tę7�O�$�T�����a��G��2Z��Ѻs\y ��Z���#���.s@����+�+W�pi����ĶF�W#{|�7������ay�4��,R�ʻ������D��7��������H�No�'���Sm�o�� g1���=��(n����7�3Ĵc
Z;�����]a׸4ѡ�x�wy����Eu��wz<�kym�3R���lż�,��8�}<�@���� �ct/��+��h�FXW)v��6Ai��A�r],;�4�m?F9����%B��MxLS@*���VD��rˣ����֎tt�����A�����Wc�EO�_ў=,'���G��WؕoÌ����$O[��o��./�"��vr��GZ��[� �����f�%IHفf�s�����39ۙ*�Vj8}���S�Ե�f@�|D����`�6�R�G�!�!�X黲=����� ���\ӭ��7 [䮢����;����5��Ư.J��.���R���'0$��x��%�]P��mq��qߊFF����B���l�%v��xhm�$˗�W)��$	lkkt��/|䭎*�Ff���#�.���ځ���,��>gǥv+��0:�8���GC��Է+w��c�˕��X9�4j�1.�U�<8*]��rC<qU��1C�3�M>��� =��Պ�

���=\��I�J�d��($�V�'� [��r����Nn����qeC�.�*����M ڱ�d}����;Q�q���]���o,GW����4P��W�Z��'o#>}-�K�j{�ib4�y�������^�v�vzX��G���f(b��f|�� Νb�iΏ�
l��cd������̛i�K�Hs��дә5#���,�34��Rָ���H?�ae%�>A��;��gQ��S����Tp�+���u�5�x�+�@d2g=���U��g�k�My�����V���6�$xC=j��P�B�f<�����0Q�Lhي62CG��m�dc�U������}�h#��q�	�/'���]αK;q�;����AV��n u�C�Ty��Q}��Fѥ���0lB��ļD�J���v���z���l~����4�������}e�z��5rӆ?̝r�����V6����\hlN�6�eC��[ZK@K+y���lG[��Y���l �l��zV�ޅ�0CDFk��f�Z!��D�ͯ���I�!]��_�m=6�߻Q��w��.�^��2b*͎���\���2�0��OB�ԡiU���t���%_@p��\ὁ9��2"d�b*�ʸ �~��m�5�ȅ���>kv�3�ݘP�('������狸6�W���G�&���f���t{�bq����.fB%��Y"N��.ΌcR�u�]�Al���'9����;CV[J���)���p��a�+� �S�>%���T�>z��ܿ�i�H>��y�qf˹�<6Z+�V%b�B�Ją4�ȞM$�ຓ�����k)�&���M3e�='S��ɍG�+���͉��3S�'���hS4߮���/m~�Y@����6���4Ļ �D���%o%�o���D�4vz�PKt֌�-��RJ�-v�Y�ePcV\�4Ţ�I�xv&>��NST,�b�cP����$��$DV�u���w��e;�)���ʝ��ra�*�{�u��9,8H0��0�n��pP�`n��!���r�h>��M,���2|�:���}:v�a�ޒ[#�"pyj-���Y#�ʃ����DA����^�Մt��U�"�Qk�	���*���}���2��m��#���5�އ�q��������C��LK8��-{jzH�j�#��Ch�܆�?���|n']��ne���68���I�6�E���90u�a<?����	����LT���dO�Aq��j«��v�}ń�B�}��Mܛ��>� 2���(G��ޜ�9���zgmi`TEOSe��Y�G��c�II½�G��x��'���(Y�X���R����t7w:1�g�Ϩܚ	R4BX�Q҄K�[F�e�$�pW�)D�F�ƾ�y��l�	���SM�FuŠa�t���}	��{-7ɚ���>K��I�=�s��%��۳����ANhY:�=2�wˋ������֊�j�"��*�����ٯ0)Tе��:u�y1��?gݨҩ���~�	͌x2�s���g~6x�`��^�x_�>�e��	5 n�1�=����LG]�kU�"�NUK�f�h���9��"��@���A��M+*_׍ �� �VT��ܙ�bN��5��MD>Q���;�I�`d"���+q�H48m��b'&������i�ӑ_�,�	p�eƗ(!b��g����Ԍ��|8�|��^	�Xp�h;fډ�}s�"�8_�#>���ȗ5�N���=!!��m$���m+��y��[�*�l�f�5=}��y���w�Н�y�N`�����1-lM[���9�:i�Ѧ[r >yl��@ԓc<���v�J>�	���3'P��^�t�/�؉�U��+ r�R�	R�{��.���)��D��9n��T)	kZ'�_d��=y �0�������S��T6+},�8�T%��8��Śz�ܶ�4?2��E���n
�=�J#ta@���GX�aR�|��d/��?�/̮��	����T�^C��a)�F:�$O�V��*���{+\�/���0棋)ʹեLSq�����{:�ǴzЫ��SZÀMsN|�N�J�AK�I����+(������N6�COf���:8���ٗk	!�,W���Ŗ����&"���>��ꁠЗ,��b��S���o�,`g�����U�����NX<�e0�Bq����!3X��d��޺;�v��h�N��~�3}��C��.ϧ"��J<��[��������,E_6�~ ��->�l�/�^f����ߊ�j,KUs�����$��s_��g٫ߋs��u�O`u�o(\8X�]��#��͞BʗӘ.�8HW���'��Sg���f��@�"om2��-���\���^ZJ��1PQP�8">g]F�ɫZ��h�Y۱��+VتT��洋����F	l�nQ�H1�x�sϩzؠ^W�e$g��7�;y�"z�pF���f�`e��I�SP3Q��� ��H�R!ULo߁��A�:�;���R�G]��rc�^u�;����:���ǭ���K���o��V��H�p�ϔԔ��!�bCQ"B��)T�V�y�Pf�ȣ��aן��Y,�%z� �;<?�ވ����e���nP���:u<�׸��Pɍ��G��nl��8,t|�7�(
K�I%|���HŔZ
�I�Fg��.�`��,��Q;g�d����4"�gZ�cV�i���r���𬡷	
�/���qq�?��<�(��vGy�u4Z� Ӣ=�V���?�"S�x�%�=�ʋ n��e������c�kFW<֡�*������A/��i-L�(��y���o>|��z���;�%@o�;�K��Rq��v)����LY��}_[�=n\*8�a�>���H�Gw]��gY+�$s�T�6Rr}���Ѷ�ڞ�����A�?��|�
g�O����4��D�9i���cx�6�m�xo�蟑T� T��Ϭ�R��y?��}��創��� K��a���Q)��?��W�q�@%�@+�cA�!��:�S�N���T���"PӈY-��lC0U2�f8=F�S ���ј�=�сG`�|�R<���]z�
e�������d�L�h�y�7�~_f#{-��Fot?@���m�|÷<�3�Ŧ���`1����jq+3�^�S�?�4�^���	�['wޮ:���-�+6S�m�	��\�,�����I.�2��A��Rķ��o�� ��כG�?`>jÌ��	Ɉ�[�Kaϡ�#l�	���V�z��;���<p�K��K7c�;�j�c2�d딱�nPm y��j	�_~��Su�W9i�RBc�g����';�}��#;��h�ʒ��G	�����ȝF�N���Mb���xw]�p$�}_�����\���3r�Oa�����a<o!=7!����ૐ߅,��י���f>~�:Y����&k��5C�Ho�������������RN&��g�:z��V'�AE��Jj�E�,�#o�h\�]7ϙ�����k��v�+�Å���D�Ǩ��Wm�!�h���v�η�yP�" 1�z��K���8����7�b�ַT�˫�k���A7��uh:\ps����'�v��EZ�D;W��i�^vꂄ��|7��b� I�14���o��E�{h�;��oX�d�M��|'����^m�.{B6��T���︓�(�5�o�~�RY�1�.tf�_�?��αM0b{NY}�������m�yV��0*s������"��!���y�ˮ�R%s�����Cu~���lk6HD>X��(;����~���H7�Z��|���BQu���D"����kMH[�:�8#֮a�@a������mcxe3FT珇��ja�~��r��׉�|X�*s>�o����]KәKP[����J�Y^~W}��e���)s�GEMy��R�������ch�s���נ�_1�:�%̋Kq~C��F��������T��x��P5D!];���9=�dRFM��b�\S
}���=�I_����W�O�"ܵL����3UeYlӋ0�<@��G��%��O@�֎N���"Um��N�S4��c�p�]�T��Dj�Zi81�	4��qu�hT���2n��g�Q�T���c���C#q�����2UZ��GҮVw��޽�������Z�@������<�����í}�ld�Gk���}�f-7���-kD~(�Z�[z[q��Q�{�����OF��K=�K������������u0O�;�}_ج������WMr1'�Ǝz=c- ���H�A�� ���������nU�:9�Ww��+Bb��y�ɰ)7ի�^��"�:B��v�F�Y_�
�}L��'2ED:MB �<��+�kOL����~����ކĺ�����FZ��7$�)��zg~�X܁bKY���$�Fz���Y�G8���%�K�wg1���?������,0�π�*��5Tq���D�왍�B�Q��N��Eu7=���C�[�~���a��ʒ���Dvr/�s�j7<)&��9�xnN�$
��}��Jl5�y��*��8�-�]����B�v��,�@ų� ��L��}�Ktu7��gɠЃȴ}�wh�p���l��n�,�<�<P�S3@���`Z�3��w
_�[:*uxGq�o��)�ϴ�M�z�,��e���j���w�>O(�s5����;Y�X����/H�=�Q��y�b[���˷g!͠��la�Z�4�8�Xn�n\0�
�{J�?�W� 6�2��P���d;�+�P����Ts�O�<�k�~g�D��ϱ`P����r�J��`�L}>&��Zխn��ޕ��1?ҎW
 �M����{�x�5=��PO}Ǒ���3�����d`'^z�|���PDY�#��O���_�m���W4i�G� �`Ae0�c�m��VPM�6���xJF[��v��d�[��/	m��@�p?��~p�Y�#��H@ǹY.�/W�*������7�h(>	߻��,���@\��+T9�^����y������[�T�Wn�8��6�a�c�+`;o�Bzĝ�M��mh`OA�J�n����\�$�uXz�3�8�<n5���M�h���-������iJw��/�3y|���_��8-LI�j�/�l�9-������_���a%#� Q��ųR���]稜E���
Q�I:���'z#���"�$-�b3�Ow,��j�i� ɆH&�To	�c`)��iVW��<�0��Nq*�UV����_�<dyD����oe���׻\Rɚ�d���趀��������ŵT�d1N�E�:V��M�Ӓ�Ee�x����g8d��*��m���1��j��ϫp��%���ea��yw�ql���,	"�o�{�	�� ��sPwQ��$ ������i�3ۇ���,6�Rz(�.�vq�*,����{3��!Gw�<0��N:��>N�y׹�j��go1wͭr�������o�����6֎y?���ꇍiC���B!G��[� Np���T�3��7�,�%���n�^�Ԣf�tzy�m��>�Z�n�cb�u���m�B*���=�4����	�� ��F��1v�N�Q��f�e��Q
�������Y�~"���8ea1F��+��ã��+i$�{���g�P���ɚ%jt�`Wq���]����.C�I�"_lH�qPQn�aN�Rj���XF�!7�W&v|a�A� ~z������E�؅��ǩe�r�3�Oz+G�.���{�j�,�>;,V���{Ͻ%Me��&�\z�L�
�9��}�tH�>�np�,�bI������uڵ���ή&щ�l���7�'@7�Oz3��l���(��'�e��S����o���KAH�nh'ϋ��*���cZ�a6;��!ݎ���5�����PY��M6�	C���@!O����*N�\�&���q"��������)��^y L��@H���l�썐Bko�!f��[�]�Y9�-���[�n]3�0�(V�>6�[�����w�x��8�&E�tk����Jw��7rN�Kin��E�K�f���.�BKPƶs�فC�y4�7m�yHB40'A3
i��s�Vh��|�}�sY�I�+9l�*�'4a8	�]Ļl���B��$R5�	�Խ��s���N�Ɯ	_��Z4[�]A^O&[WjMG��(�h��ŋ�Ze��O�����g�m��>��nS�>����L���.D��GJ�.�)2ϔJ�yf�����8P���"��� �=Y[��\�S�Z��������͸���^��-0��G����.Q��b*j��s�uVPe�(9�����3��ܭ�u���̲k�v�����Q[ĸ��
k�a��k����3!Wn9?�2�wA�~��o��M$L��/�![��7�Cȗ��j<1��׌YD�6i�!�u��N{���Ȝ�1�,S��|�r��BpA��'���	ѭ;�i�{�7߇�kJ��9�:�t*�6���E��"��#��1|��������4��Ͱ�ʆk,�����C��T�f��&�1<�i��O�	�y<q�mq;8�6	����b�Q�q��f������,]�p�ֲ�E`���	D�) ���Ƽ|��v*�����6d�������*C�*�WOfoY�U=Y��I,U$�
V�6X{2�N��_d x�Wl`R����2c�j�ɇ���"e�ߘ8���#3�͛���lK���M�.���7v"�k��?���=���N�O�BK[Pl,�,�M�Z80u�~��^�+�Z���֋N�4�D��2����jf'�1���(�>�	�V�7..|M�����s����2ó���2�j���s' �VxQ7��f)	�u��5���� 7�:C��-�m�8�_��!i�
�i���:����Ə
{������H~�0ھi�j?��X�MP����|<�x���kV�`.�^��^� ���3<1��庈�D~���o�!�&�Ҽ�+�A��\H�q\�Щ��v�Wvmv�Ң�8 d'he�����8����p�+c�r�>=h�GH*��qL�[؄���_��F��=jNH�AU��Y�G�
���9�n�zG�.��D��q7��9R_wT���z�;��3�T�����"�zY\
d)ʭ����AQB	�ss�!� '
յ��LJ �ZWW��61W�����7;l�q{�㧗���{
�b�#��s���
�t����d�t�G��A������qYl�,�W�g�%Rf�y�mDJ�4��w�)�n4q�#�z~+�/ayy�Z� G��C:=.�3�)i
�c��5�R(��H$t�`FH����3�����W�N��!�6�֣/���ѬM�����$��xo��[��{���	�'�D'�&�*�m�ή�63U4��y�9L{��B�<q�� �U�����ӛ�Ɍ�K~��h��b�$,� n�}�% G���w����]�G..E1���>���[9d��L�J%b`*����ףA�mr��X�V�<?�P�h�ڞ[�/��n	��=��#�[�{�eOP	��&r̹%�T'1�*���1KCwh���ۓ����h����6P�Q��#3rW� �p���
}W}|�P���龗�Q��fp��4�,I�+t��e8�شw���|�I���9PQuu�4W��VD����UU�+?W��"��c�6��-#-���I>85H5�`���mF��4�(�Уr�����[�sGD�B(�ԥ��=��E��"ǐ�G������,$E�����<`�@���a7^o^ڦÒ�N�A��Ƀ�f�Y��"�]Mu)9��U�Z��=pWb�5h�EDV��e+��`�r���>1�sNlc��rBx��󛐱�N��U\3���\��V�?$�͠��R��_H�MuM�N^=��{u8"��,�}��i�Y�rt�u/���B�ݲ����w/��$,�2�%͍�Ӧ��yDT�v��i|`�/^Q��I-3T�k�Q�}]uc�c�"s��vC��'驚D���u����q�{
�&���,��៛��;>��)5��j��ds�!\�خ�f�"�%k�Z�i�}	b�4~�mc��&6n:��;�ws��	�ټ���y��u)fi[��2n𰧪�-�3d@Lf��a͈�r��\D^DQ����HLf[�C~U�⵨l�;\��ҫIU�^��9*��yX�nO	^��K��+�\�R����{�V�PO�X^�s_����~��w0˶�����ds���<�C���K�ݘE
A��+��5��]���S�Q��Gz�܉��������oR��"�M7���c��u��
Ҹ_��*������=�P� �?��'H���Eg��`�_(�UC@���'�4��88�k����aJ�c�S���>#��d�e@%�zU��4	0"	y:o��k<B��f�ii��x!�.���a��8��WL2��x|�����xpM�V�O�p���$v�ԴviA���Ri�]A ��S�>��R!0�� �(�vkDVW�����%Z� �M�+��<ў���y,9x�&J�&����i��?Q�[O�ۄ'��K>I-��{O`a�g{�]6@�p����7uN��=Ά� h��|�DF�
*{�m�y���������GV�x�<���t������_.TJ�[%v�z~�k73�\D�	�{���Ug��� �
R�*���z�X�=Ӛ�RG=SZ��_�`�au~��mj�͍"zVEX~=�ݕ���L;�+�z��m����ό$<��|Q�/��iy��j[Y ��_�� �R�H�z���5��լ�a���S�p���ƋH	�hO�D�auuJ�� �1/�'S���P�ۗm���Wʯm��Kd�U���d!\s�u]����n����n�1ث���]��)��Ge?h�a�)`����W�,��&"����[¢֫�_*�T^E��]ίm,6[	������%�ѩ��*}f��v�d���N_kC��
���ql���,>�Nj��N��qwME�
큻@wN���7&����s�8�D�D8ڑB[.��_�2�AZ�8Њ�H�l�b[�4�$"�ً��a* ��g��."�Ch|�W4��_� 9���p��稼�X�kP'u\�AWb�����S{�M�	�nYy�ʋ]���D��q~V<%�����3�|k�4O�)�����ΐ��޼�R9�����<�PH6#e-{_A_*:�;Y{������K�&F=W]4���__E�d� X9�MT�W�ۭpn�	=��J��i��pP<U��ד��Jp���=��j�G�p���(��%3�.m,��� �壳�A(���J�#�	�F54�=]�qa@��xI� 3�΂��6�BϠK�~X@�O��	9����H2i!J�E[ܭ��u���x�"�]^=.o�m�!>5�'rD��)�kT_�zg�[���LM=�J���]�x���B�$�ݠ�K�h7r�#��h��TUD�K�~Ng޼��s����s|2h�#��1�&�d��_����A������� �]-h�{�7GH��=t�w��oM<p7V�`W��p�o��������d%�z��!y��)��	�秷*�w�F^n� R��H▛����D��Ή�Tu���:�}J�c�[�Fu��+� �֦H� �ې@g{�<��4B0��"R�	 �D.�J&�$,��"��0����&W#������\0Sw�*k��-�_�֜�2�unW3!�7���_���tw��PA=7�cx��l}��rH�[���4-"؅{�'v%�nm���+��]����>��7G ��	_����Aq�O�@{��E�M���9�y��N���7=�"��iȄ��?}F�,D� �Y�k�����-�hk����pl=�敽ς�r4a�u� O�C�'PN�e(+濐ph̹r�Dg@�L���x�E�%m���m���ߐ�b�!l�n���
ԙ:
#��$ه���,ح��	�1��M����IZ:똞�3Xwo���L).��x�ZfZ�f��Us�R�i>�i8����i�}NO�0d����4�Ѵ7�=� Go���*�{^���M󇫈��\.�O!&��,�^7�C{�3��H���/]ޝ�rV�(q8���B"@D�Ά�	�_�c]�����nm�d| ��f)�	��M"^����#ӳ|7�q�nw����bs1g| a�Dߓ�j�M�=?+Td���O���)80���UgU���Ő5�(�A���-�������5�B���7/=NB���v��VT^�Oq"
Y��h,���皆o]�`��ޏM�c2������y�沤�P7R9�[�L��u�"�yh0R�%
Z�@M	Bh��d�.5���O_'q��(<�&Z<����P�Pn&��`�dz�����ƍ�7+��E��~���)�dq%sa���#�6DN�j슔�Y�X���Λ�2��}í
�t�yF� �WFXǋI���$\���f���c.6/��CǶ��)�V� �;aǄ��?`��{��R�׏M����٨���x�bm���%���t�˴���@����y1���
����;�7��hρEv,��Q����ʃ�r��؀fk�bġ���)@��p�̩��nׇC �\T/��D5z�;`���g*��ZX���j���>���$%�� W�_ ң5��L���caN�Z�e��UE�؉Tc���ւԙ����҉����7>�Bxq(�fn"�{�P�u�(��@����̙��O�Bx�V�5ԭ�P���U�vF*�9C���faMqAv��މ��։���8f)�ĺ��Rs�c6
���X[�%Z�.�!� @HM����(M�z�E�wu�����w��1+,���Bݹ5�Y�.(�QE7��g��^����� ܆;��X�a�i�G��?`����Ӿh{��m�����'���9l�B�'��m�ūO���YQ���.��4k�1l���+�\�5�y{E��b��̀�����"������߿UO(�<�1Q9?si�E�aNTEb���&�s�0z����9�� ]_�����Jh��G���u����)���9
��i��mBnD'tww�|e!�����V�&�����i8���9�MeM8��1K�`����!/��n֦��q��H�� ������C��(�I:H� ���B',���7i;
�+P$��?�&���45�����PQ�k��UF��˖F��v���z���-C���]���)�\ ��'$��&�QS��6��e�Td3	���ʩp�}�.���^��8-�W2�tw�B�|��Z��$&vZ��Mi��NL6���m[�=�
�'x��e�aMf2�t4ֲV��x��Q��<�|��v�Q�FD��e?�kzX�O@�(n�[�{уlL�e�a��Mrm����3q�#'gv��1]���?�G���m���G�杶���;��������w-O>���\�U���Sv���=���xe�@ a7���_��Հ�+����;��h�U51��Q�LrEd��'f��m����?h4H}[�v��U�ODb��+4v���np�(�2��u���&'к¯��w�
���y��M��
2һ��J�����P�P
�����.�j@ݾ��R��p���.���7�I���gL�r$�k%�lN�cg�� �'��޼⭈Ϧ��1��bگ.��P�T<y.��I����D�p����!��n������p9d�h�'�d�< :�[����^����LW��>؋��i���޵���vK�O�K��R�'�1��]�����+�"8K��Om��2���K�����[����?Ќ���
�����S��Dۚ<��Џ����P𵉠A
J��0�,��۽���a�3���l����q_i�3���_�Y1c���s&B��V�P�	`�����+�qZ�4����d�+�W�� ��J�5 �ӬH�й�0>u:�����H�r�
�'��#�)��1���w_.����8������j"�31K;O˵f����7M{K�>��,#�;�d����1��EB�#������4�]K��p��ſ_�iw�a��{���� ��wP�|=�Y���@il�ʻ_17�\W�k���e�|	��rs�i��L�J���"���
���gIĉ�C���	�͋���/3��,�hD�IޣȊ{%�j���t�0X�:wQ�&a�c��ZR#�ݐn�\1M)���@F>��IW�Q�`Mu��V������,�V�C�����O d��[,�sr���M�
������Vf&Կ�=�B��ߜ�0!�k%΀�	R���Ң�/�=�|���]`�)ʠ�U]�D�k��9���7�FmlW��p���"�h���VB�5��(u��%�b+,n�>��.�T��q�7:�	��t�С��䗞e�ƍOl������eT�L�B�����]#�Yat &��cC��AG��o^��|��e(E3��u��>�A��CJ(X��-j��⃆�ӫQ�Dh�С�XªAi�~E�Cz#����b)�;��M �u��U��Cz�?r��x57��GĶ$42�E����G�����1��
 |mH��Y�����{�"�p�"���t�dQ/�����%�q���Ec��Մ;�!s��}g lPSO��T��u+���Әd �wy>��RMA��(CY�Fj��Y�N���L_&���h�.���t���ݗ��qZ�`c��� ���SGpq���+�'U�� �FEr	��n�7��EQ��-�gdA,2!n��H��m)n���^�l�ޚ�����Q�L�h�`O�o$W�������{�^4E�D<�W~ѥ�Iɾ��w�������Qjiy6��Ŧ����c>z��ak���Փk\��v�=��ſK���@N>۶���	���m��%�7j�]k��	]��^��� �Y}z�3�7�()��^t<�c�2D��[�^�y��>,K���֫����1���Z�*s�2i�TV���AO��ҕӘ�7p��-õ���v�i�3P&�M\����hE����h��^�Q�m��J�1B-��$�@�\OG��!�nc:iľ�)Q������.r#w�Qe�p䧍c�w�Ś��Yf��Q/A�Pz���æj��NJ���3��X1��x���-��9��:'b5�'j����&,g/r�\��Q�Fg[���a#�s�	�g��5r?��7�#D^�-����1s4Գo���H�)��R��4�;&�5�DݤQl������3���#�|��,����,�zS���ƌH��Z�G s�Fq�_�[䛷�0p\{ǟ������|�{�[{)�h�XV~ݔ$cy�D�ޥЎ������?o�:�.z��D��r*�
��ً��8x�~@MMr�D-|�bbX�_�z" \�qp
#g���%pd�nR���9+�!�u�8��}�[���i��!�E���Q\x0��	d@#6A���m4������t�V)Y$�ApGkI�J2ßd�`�>)���+e) ��W.�yz�c_�j$��qyg�w6��d[�Y�Ҧ
m&q4��n�߳���"dd-a�ږ.��Eag��A�9uw��&��B$go�����i���॑�r�(�}�5A���v��!K�*Mh�[$�K ��|5��s1z�K@�H��x�k��^��%�ut�ʂ{�o���Et�1wԀ����Cf�\W?X��N��\�=5eYl�X�Ѿڼt�F=I3+�
�B�n�s��Շ��`��\�s�OJ�73?c?EZ%Pʨ3�<3����Z�e;a�K��������Ϋ'UY5��zEF����<#t�a��j� a�obs�A$�,�M1ɏ�������P[(j�1|waK1�a!	xkI���t�jHn<A�$�@��bIOE�>Lb (^̚w-'QO�S��0�N���g���k)�6��cv;�,�25-ϔ�Bn�~�3��xU���g~6�����%yǓ�u/&C�dm�5�^u�޿����tM�
;$zn�e&;X�ܴ��Um�,�GC���~s/��5}�f��"�,�<�`RE��i�p�<H9� ���۽����yŰ`��%-Sc�T�l������/�J��"���Q-q�C0��p�i��2U�����"� 3�%���r�6�� !Nk�����b��!���ھ/AEI�U�����6?��&�V�91ay����o�
~�N=��������\s6���r�R��tt�6�ƑL�7�����Kә<��Iy?�X�~ǥӜ!ټ�nD�1�Q����[[���r�K�+�˝�DR@�b�����)�4��7*掝�><��U������ɒ��=�~Zvǈ2*$���[���}((���A�j����-�_%�3aޯ�]��&�b��bODT�f���C�c�����Cg�	>��>�ޞ�S���:A�`���"p] �#X3�U.gBG���#��/Z�1�x]��61>K*:�#���K����v��Y��ӗ�H��W'�����+�ܦZ��_7��@�����Ŧ	S;���ݰ񅶨w��)���@t�1�|G|��m�!��@�\ɉj��C��j-M��Ot=��E%�.Cy�[��|��G:��S:N�s-�����88o;�����#����t���H��b�m��s����Ԗ�o�nb�ٳZ]?������q/�w�2A� ����Q)M8��	�ՋtБ�|:��*4�;�k�x<�p�#ʢ�?�\�9mw lRkC��C�� �#���R>1I})jAi"�~J�NbhX�I�������y�f�o5tlK.:������ש���{��at���<ծbi�J�?2��
�j4�a�ݓ�5�B�Đ�t����,�]v�St���M�,%��C|I�/*���O����f�b��c� ���o�5�@�h�^f{�0Y}�����Sy�,4��/�n�*��1���(::�E�	�¿�'B�?2�(/�k&������~����h��D�ggoF#}�0�9�}�Q��-�To3L/��Zg@�y9S���@��Ҳ��@h��*ls�Yvw���zLΪc�Я� $�R�ѐԇ�4|L*&����FFKjw7�Q����N>���'�H�����76���$�e��im�a���uI%��C����j�AT �D������${�a=��[xjJ��B��㹺�{��mO�@ajp�Q�^i˶���s�B����[|�r���T�m��e�\84������f�k�5/f�W&�rI.����>�#�3�.�ٴ�r�R��tg}B4�܅PJ�±������7�d;;W�˔$�[� !����-.���i=+��B_�P��,���`];��a��J�`��%�ll�nK���Iև٢��މ,W^�i�*]BkΫ'gO���z���.�]q5����A]��2՞�F���z�l-y��w6��\���3��:����-�`�Q��z:Ax�'�\��L�=����c��iġ'� l&;b<�y�4�{� 8���X+�!͖�\����ڎ�(�$�ZM�|�O%%�������;/i��Hx�r0&*Ǐ��طF�'��=���wP�D�C<Ȏ->�c���\Ga�Y��x=�c��wE,���RQ���%�4�ǧ��lS���,y]�r0z���<�(|�Y(����1)��́�&�Vh��Rh�Ѧ>k�5��dh���i˃R+Ե�$8e{���W�g��H�/���
����+C�M�8n:���4qh:iGX��u�c�n��Li:yӦ��&�Sjv�	�,-�\oF�d�A����7�2M�@��olBS��Gϯ�� �� ��+r^���S���d��4�Uw�B��Y�5YR�1�5�X��Wù�� .�a-�$yR۫�6K����u9Fp����r7Z��V����@�4Ş���#PS�[Pg�R��ۗ��vx4߿�
�{K�G�0�P��z"��� 2jJ�.��!��|�ϴ]��LR_TM ��J���o���-'jsQ��z���C�
�8K���}M��/��$]�u���=]\�ü�ݼ�l$!{Mp�b�(���B�����ke� �Q���Y�$`��+��j��a.�>yc)S
�7���ɫe�(fE믁6�F��.�m�,���.��N�N+�[K�ʈс*�$�ْ�[L�B�\j�>߻�>!�F���gS[)Sq�����:�����Y\��X�'��
�)����^9cC��`t�Ȯo�ݓ�;���yE���3�� ��ڍ�=���`Ux�5��G�_�Rl0�"�1�aE�3%��Rf.5r?�֠5�>9��#�	���3�����5i���TK��*����˷�r�1�U���uq�i[����������ԥ�j�pO��zpT���v�+D��{���Ŧ�	�J�L�9�U��"ȫ��ZNǮ;X��<��a�N�p�^R�ocSW�e�k�H6�t5ޗ	��y��GO��2fVqiGXήb����G�����PI�m]E�S9Fª��*��t�>i��{ ��\{Y>�`���Tb��'�0x����-*����\nP |�J����C���)�l:�U(Ьh��F�����ϋ���3kx�')jz6�WK���=}ϥ��
�G_{�=�.����x�{`������G���m����4�;0��1쓇�r��6[��#F���ڽ�pǦ�|=�"h�n���>�J��qA�D� G���� q��Wı��jq,"3�d��"/^��rC��=N�zeY��Q=����M�㞌�\R�G�m�l|�����B�V�ӄ�$M�|!OGp�A�!�陮�����xd�ڒ�ĝ���!�i�N}���ͦ�>�E���I}�`���ù�{�w���	tɸ`���Z(PFa:e$�,�+��~8�}��k�)�TSzy���<��/�:ק�/�ҫi����0p^%|��l"D��o�l�G��	�E+���|�������+�5G�u��
�jM+�3,-	���͋Ԇ�M��*�V�?r�	!�ň̈�|�C�N�v��j����m[���hM���z����z��k�);I��Ho~��H�]�^�f�PY���<2�]�q:)b�Z
������� y��c��$��t�Nr=o�S��W�� ���_�lط"3�e��^�I�<6]�J���:�#s��w|֏F�Jeş��ۀ��y�v0O�����1�5�(��,������_e���B�g�(��o�fE���-$�FhA��۬�@��0��Xlt��ޥ����R�Ʒu� �F�9\'&�j�+������� /��� ��E�":��YS!��k�P�c[��\K��z�-����"u��%	��~�b(��d��X�"tlyN��l�բE5�9�jvVI������6�O�ӧs52��m�O���B�������޼�SX���T���m��w�����Kͦ����KF&dQ�C���
ݏ���?��E�{�N�3!�O.>qȐ�B���.�����8_m�%�Y��ʬ�i�K�
tV��*z�vj��_Ia���&���_脟R8Bw��@6��K��#�_�W�|Qo����vlo;�Ge��N��@��J�:ϥD�S�`�!�4*�
�f=����{��Qmƽ�Lo�72%�8�K��埅gv�OѸ��������Ok�k|�~�m��R�����%�XUW�_�ɪ	��Ofo\R!���������&��'��b���*�-�Q���N�E%u�q���_���L�a�z{呬��a/>�F&ش��n�_����4I[t���D�$s)�U��N������D]���A�@ S���_?�Ѥ�c��z.5�N(��5áp��C%��i��Af�|�`=a�Mˉ�P�O���ߦ.���c�Fj	=ĸ<�]�r�QT�DF0��Yw��'�kC|�ܜ3����$FO@>��=��Ҭi������j�4m��-;U��)@�Z�0��7B1�k��;ix�/Δ/�V{��g���}s䦲<,~���gЌ�ӯ��TS�U�N��~�� ;N���;w���v˝6\�_?0Q�?�7�܅�"��;\71�	L���ȝ:/����t7L(�ڙ=ˍL�E�5|q��j�^��GbD����lu�}����m5��7~�2�@�6%�`Xpa��=�M���%���PD޾3�S濋����4�f����/�/�Ң�J5JT�w�c
�[ �j<.o○ jU��R��x�6K�Ag��[�v�
�jWO,�
��)���9M�a��w��l�s�6*A��Iol��|��,��Xo�����o�C1G3Ϧ�����Q�Z9�O ����j�y��=2��P��;�+�8iנ.M�^��u��Ű߇�4��O*d�F�*�v#R(�G���9�0
w��um�ъ�J�g�m%@�\�0(���������^��6��%wB���0XM-aj%+��D��j�t��{{d�o�p(T�g��$���h*�ˌ���=�' �>�E�O��HsO����½��*K�;�I�҄Ё�2�*մ���8���\�}��o�v���H�|� �\|��e),}'�i����Oē�!n�r��@�KT�ʠ��C��y�Y�������ՄN�-�.�]h���4�D;��I�ku:	�I0�q/M[�w���;?^s���(#�G�@�,���fJ�4�Ͷ�I,$��{~J
�k�$�T����)��mWZ쟗&�i�[��R�y�JW��P,�5+�(r�m�Z�ɬ
�`��(W=�z�u����
�1�e�|�����#�� M��t1�G�n�Kf��~%���6����Yv�Up�g����>6NzU�������|��sF(Tt��v����2��&$��%�Y�0������p��џ�po��K����W2���X�T��È���/����Z�ݵ/%Q�+�r��Xi,�YW���UǸ�<�7s/C�Յ�^0Gq��TrpՆQ=�<����7�CiS��+�@-J�;��VU�~d�}e��R<G���i��,\Z�J�4�
EIt�rcI�����g1�vC�|��v�R���ȚN79A�2
��*��}ǻ��H~�(�dB|S��0f��Ո�u�̅Uڢ�������`o�����'�Ӹ�~Z-�J��:b�,�_od�`�$t�D׆y���{�"�p�d��-\b���/ۇ��ψ�v�)Ov�� �"�4�e�G�֥��@�$:�U�E��s-%�Krj���g��Ȁ6�H��ox�:�D�Ww@�������-!�i�x*|�I�I���<-Qizة�em>K�9�F��k���|��xo^�T�F��A��P̾N��i+�V���O_����`��l�ʮ�K�&g^y���X fU�(�d��o�˪a���� ����e�5z$dcI1�A�נ���z�%\e��3�{ܞ��OWR�&�^_�z7�m�R��B�f�Uw�j�z�6��8:������R��Ä����(�U��v����3�wq㠈R���.�Nќ�y��Mz�'�$�����ۺ�O��ؚ\T
ɃѦf���_=�u
{4}f]{�h���>�|����A8�J��b��ﶾ0�4}]y�{f�'���U�:#�x��1?�� D<h �{�m�){��5�\,�Ԝ���i6��5��w(���`A�3s��P_���3.�v�j�J1(�� A�����1���DY��/�PJ�I�b�իW��,������� ��������>�x.�;?�4���		��E����,l<&��)��������������?w|Lǽ�G�Y~���V��X'p&L���x�D�4�.�2�|r�BR;���>ԛ���&�a��*�Y@�.�����I̕?�=��R�J���������t���N���~��RQ�Q�N�nI.�(~X��v�{F\ j͚���D��K}���o�3]j�b�t�ǿ"o���w��G�n��ﾍ�<���
��"k �l���(��U��r�&�"O��L�c���rd�oŎ�hb�u�pMϛ��H�o�~QҜB�R�Y?��2�������n:��t�#�$�q��k�o�/��s�H�煸�]4� Rn�ѤiC������W3����$�U���c�[�iI��R��~��\ࡹ�6c�AΨ��E3���:M��6SL�-�K��f��W����9�#&s����;�5GN��lT��D��B&�z[���D�8)�%�����E�0�'Ĉz���c��U��RC��a����y@��[��IC�%hi/�{R4=�H9�} �/\��;~ȁ�s�V���q��HIooAic��Gԛ(8��NX�oU�z
�^����42�K�[��O�������澼��cP~R՚�:%1����e/M�`�.�`��*�49��sVZ��BԤ�9���S@{�?_q��A�	��26w��Qψ��L�GJ��B֞Th����O@�n����������^��7�r��umLH�iY:Xm�#�^�U��(]$	7h{6/��}M'�.�&���=��]A)�������w����N2
]�jz��QN��9*2e8jQ�L<�c~Dj#�W�Z#�I9�n^q#�������'�Q\z=�oǫ{Oȅ0�7��C����N�t3�ke�� �IS�~���|��@�k�8߼�A%�,�%�&�:�Z�Q��z�:Ż�H�>ot]�+�I{���4�8����@q�= ��.c�O��C�Es��dKޜ�i0��.k�V� ������7�G��
#�{p�C��WT�����g���&�B��ZDVB���Y�#��'�{�*֪����w�e�L���~DY�{���y�B��`G�N�u�'�7Ǩ�떿��;�Mc��5Տ�h�J��.��@N��iA �A��҂�l�a��eE��j�U�]G�/�A`l6R4�IU�;����̿��2�A����}���C��-M�b�=�N��ˇV;X�OW����l�EI��t��](��㥝
���T"?
���H���S�ē�̍Xo�`�m��6>L�28��j��@�WR�!;U&�g��;|���Wpl��7Uҙ-����.�?�4C�x�j�Y2'�-c�1d�i���v'��.��֥+7�{�<��c����6��f�/�y� �Xͩ��%m���Ғ�G��7s�_�č-p.󄻭t�O�r*��_����J�)�	�:��ēw [�'OU&]i�d�� ��=H�u�s֚��Ή֝J�����v�����݈��O�\
�e���	����2�����܎��U:����a��	]r��k$��N�s�_����������Ҟ�6�1�����"L���͵u�u�A���%�<��_Ѷ}���N����e�\�w~�z>�u2��N-����ҋ�PG�mx��x�f��s���9g%��񈉄i�'����s:#-��`մ�X4��R�����07�HZ������M�	J��$�[`�`�0E����]����Ć�4�x��t@�~���%����������s"-?6V�Xx�p�N��:�.�>��)��'���C���q�F����J�+\Q��!�pW�4[���_�`���d&u��5�n(NgC3G�g�īzj��
_^г	��*�5�P��AI[Lv{u�⬉��C���l9{;h^��l�ͽ��X�>x�fK.�|x���{Z�ƛ~��XtG�G�,t��#��rrkŖwg�P��6wy�߹��Գ9-w��9��TSv��jX�ޙ@,��'�殸t�Y�F�Z�f�qk� ����>}�=h�d]�L /���u�5R^U3���@�ba���B0�Y���\*���Q��4R�#/�x�2Ҙ_�9��D^��'V%P5�u��-���ߙ^��JJ}��S27@����fc]0bh�n�X��D��x9�T�a*-C��;�R�LB��}��3w"�l�n�H�2���N�'�Zr����YTJ/ŀ���_ͽN�b�<�$J�#�[V�M��G]F�t�qs�	��$�%���&�����Q""^�=T
ǚ\�ɑqv1Q�jM"�$]xD��g��;i�[gZ_�l{�\B����b�W��z���Nil���W�����Œ�����@��pp������ 8��ԅ͂�����Kռ6ϓ��ܩ�Oۆ�l�*��Eu9-���c��d/����aA�&dxky��j`���G���tg��^�����x��b��E�e�J꓈�Y�˻c�p��ǆ����G���$y�Lr>�,�6�+f�/�{T(
�{J��t>G`��?�m�X�$��;8���"�΅yQE��w���kF4�lo�B�sߓ�XNDam�px�ڞ �K\Nj�eٵ؆pD!��ǚ��s�MG8��vz�����3.:�z0�I)b:y���O"�k,}mK���%ӫF�'��U���V���m��#u��n��A/:��e,����>�?��-�p�d/�?�,�\�'�]�M�:�mC�.�sRG�x�҇���}�H"�3�U��.� (^!�c��Ga�qъ7E��8�`�؂���/�L�Ǿ��Q�^JG�X�-!Ut�ή�ۙ�+_�G-$֮UÂ�
%��ai��7�`�䠑��q�=����	 F\[�����y�Mz�⾫���w�S3����[r+�wZD���C��AF��%�'	`DY"����J�a�b�Y8��\��#,�%� �������w;V���YlJ�hf�,z�Vߔв�}8֔\�ۢ�t���t������o"���A�=�ጦ֗�W�8�IP���+nm$��i�*>@z��JH�y��'vz���s���B��;�舧�q��x��6�s[���]����#����(� y��gq���+aȢ��w����ʻ��1�:ԁ��ȯ��`�[T!�: �38���S@D��7�����0S�YF�P��20�K�W`Ee؉��J�N���Q0��*�9�n���M�X�8T�)-���Ls��S<�ށh��O�1�ɠ��7Tf�6�w�x�]&�݊{�a-Z��|������m��`�FA��Q��iYuN��jHG�s�h�1�\m����F��!�.�!���6��!��lm��,��!�aZ02�=_Z�?�Gi-�NL:<�N���i�ʑʠ�\���2ޓ'�T��Ƣc��-8ׯ�b�`�3$[�������^r=�{1�|#�T�u�Wա�5�p��G�؛%M�L�,��q)E�Χ�s"�41�#�/O�4Jt��R0���oD� J+&0-7L�ED�R��~s�
m���'{R_k�q���P��VZ�tOt�@d"W)bxUJ� е� 6����l%V�͑�%�W�5.��i_�o�FGYi�;A1tx͎���Ad�Y�%�	y�|�;�����m�'ϼk!>��W��6�\[���<9@`c~���\�,��D��Bɾ)k�]b.�KG"�q��F|�������Ǜ%�����BAF�����ꪝ����a �p�>����A�����'���*}��^�.�;�/�C�D�M8���4�X�Q�����o,Q;g��k�O��iZo^z	�l�m�N��Y�Zb�/�]#G�������Kw7�3' RY���\�F�o�TXYou����cni'7�i��.��P[C�9�ڦ�l���K���`:\�delId�N�� Z&�t}sj��dPr�+���ɳ�r������ȯg:�ŉƝ���
\d�>�d}^=-�??RN}�M��sn��3t���I�װ;�`����ĵA�
T:9�y�,���M/F��O�����D7�=��iqa�A���05�K~��bFς�gm3e�(3��C�c�d�!�����	��-5u�����% G��e�~�gM���v֗N���2�A�뺘�/wt��O��Þ�7��Gݤ�"@B���$3��T�)6�Y�Zm)��]���7VG��
Nтxů/���Y�dmO�R9?;�'Ġ#~F�d�ҡ8+�ҩ��;(<�Ow,Ӷ��T5؎�Ы�8(g�7���m�N����W7i=���m(����M�B����!�C��I�:���)��}�k��m0ډ�@\��\�ЯN�_��j�<Rt����0�ή�� 8�K�
ް��j�ck[�)��P&lA�E��e:1rj�����%��#��Oٽ��d��`d(<��92E��f~���ss"�Ds���/��]V���(OY5�]c��bҏ'��JS�wƓ��}m��0���lH�Q��éV%�GCxz�s�1U*>6{b�J�4ƚ�*ߨ ��cd+-�l����C��7e�b~i���|��␋<Ф>d6�+D���a��л��ߚ͎��疳��r����8���*2������0&���SM�ỵ��F_�?����)Y����hߞ��r�5�d��t�R�;��֊yz��?ϕh}x�UtV�;vj�7��U�o���x�ڄH�Ɇ9Oic���)��ÏԞ�O�t��~h��H���;W�����E������YL�o7d�2�]�-��?d�_Ki��Kj�����h�\�ر>A�Ȗn]�B�)��n*�:���Q{5�0J9=�6G�;;��"i�K7��U��iƋ�p<�����$)J~�ǋ�$9Q5�4Y�g�x:
�c#@��U��"���2k]!�G��g2�8̑<���j ���8~�t�X������)�����u�DaU���% R�>||�q[q��T�3Zf4�^V�CK�C$&9�$�Ds]���G�v�O�n����k���9{�H���j�+�~HT�A���6d�ڤ���wo�4mw,�@��;��?��T��+�x򉽆B������E�UiyA��;�uQRȕ�[q3�k��q���Vg����W>���@w��q�	m�=:}��Ll�l�pt���5�0q���t����Sw�n�E|Ï[��2�t�,�骣6�n�����A�NiyI�_~�;���jk�a��	雏U�[S��Zޜ�RTe����"��5�c��c��Iy��b��˱]�+���r����"�	���Ae�����#�v5���J������q	�|�����y��>��Erw��F�� �dw�W�K�~M1��9��?$8�/��yûsWTOY�@aF��:��Mp�\�mf�\@������`h"��C��3��|y��d� ����t:��{��/� ��O;f�\������j����bp7F�
4+��y�$�,�<1���C��(�VkE�eR&TWe[��3S����N��'���>V�q9+萌 � [Z��td�Zc:_���I��K;��~�++���"ň�Q���0*��3;.{pLĔ�Æ��;p�\�2�o�?�uҰZ6r�����N,�vI��v3/E@!V�j[����+P����P��ӎ ��T�DK!��'/��4.\�Y����1�j[4�39�@�������b	ɟ9,%�Ok��i1�\���;���Pg'�V����f��J��&���t��A?k��e�5*,��L.�'�⼠gj��-%?I�a��t�\��.�90��-��3�S�^��A{��2%4z߂|� !$��P�ǅ���dLO:��M[mY�����q��Ȣ22��kU��i*��MlӁ9�MԲ\�+��7,�W!�O�Zq;>�H�hHx��R���{�@A�c9�Y?8*��4N$6u>�]K�x��&�}��xԏq���!ڰ�X�^�v�6x�q��G��	m \�,�Gp���O��8��&�F�H�m�Y�b�/���h��Q#P�E)��i�`� uVO��ꛍ��+�e��1��iЁ��!D^�đ@e�.�)��P�;��n�%��`�����ȳ�U	�%�{t.�-���`\�:?���ݫA|@��$���k�d��XJ�e�F�D6L��4�Wy��a� Z�\Wn�	���D	�
7�$l��B=}�F_s��<n5���k��l 0���M1��땂��5�5���wn�/����^�C���o{q��?q�"�v�v'�`�_�3}"�؏$��w�Gġ��(w��꡿W{�i���~
�`���V؅߻x��Ǵ �W��ȖǷ�����/�b�3]�jӓ�+T�
&�iQe�V���4�_CgE�LM}���T�Z�*h�B��*y<���_FI�lY�'�o���E@n|e�W�h/�Y�E�J�n˼��!ry��A({�K�h2=�R�K3S��VG�1�>�ZlI��zf/�qT9�w�:Ŵ�� ^��HD�2B��	UP��r)r8~���'ƠS����?rNNwHEa|�\UUn�\��=��	Z�2�Ն��-P3/fOL9���#�@���vY�6�����7ln�K����j��D�,uK��J#AG'J|h5.6�,��:��+C[��.������-C�E������7�* 
4���*�9�%�+gQeN�}�
P��&O�\FP�@�+�_�7���*V�H�1# �A�d������|{T�%�@��Ԭ�������\��%D=�^���yNd��.4$���<��pֲ8�������S(^HmoU��{��;��J��
]��䬨� �b���>���a�e�$!���<� 7��I�ǥ����]�,bWT���YN	Tl�b�T��&�����������ݞ�3���@{_�P�g<�Y�g$F�?�~]g� ��6��&žc�pĈj8��d<��b��Ǖ�9pX��eJ�Ӏ**�b��Ҕ@	6�Kѝ!�87����Ç>q�8Zff/�)�GS2:�*Y�U]ֵ��K<���a�]��Z^�ؿ���<v*��^�Y�	jS)tB�	ѫ�m2�Lko�v��L8������h����5Q�|��W�H�5k��������~ES��8����J�i2�Bs�gÃ�)p�ʛ��,N|Ä~QY���:zAQ_O����;���a�U����9BW]�*C�`:.�v7��M���z, �zE�SJu�m� %#���W/؁�e�2�_^_�ۂ��yIr���A �
(���r���x�|��h`|���Z�)oG�$����ՋR�d�Su��˜�0���y�]X�ؽcۥ7[:���~�4��v�%g�r���g,
�LG��8j>��3מ@}��bH�"��2@��:ݺ [�C���r���N�s��I>O~_�� CrD��"��=��8���I,���Xd�~{V�N8��5缜9������򋺲�����`��h�E5����)��]�!7L���,��o��OS)�#�ek����\��u���m��|�/U���,Z�4�(A]L�N3���]��b*Aj��Y�R+�y(�6�4:ٟ��#Wo=�}f�� E\j1����褕&�s���K���w	�ԥ�{��t⍈܂���=�zĦ���.�ļ���m�g��$��SszIy��4��3	�7��s2I��$�n��A^���yJϼ�mF����C�����+�iv�;i�����͠:�!�Ҫ{9���}����J�?	��ͱ��c�9D�c�ѥ����$l�P��U����w��PT7a�[P�!_5����J�rY!(��׿�S	���mE��o�j��s��j��D��a���-��MP&3V��+9��	7d�-"�Ƹ/��A�NUTM�W�
��b�/�\4w�kP*P��f�r�G�G	���͢��T���~oJ#"Y]͛���5����%�l�	�|C��F�g�0�0�ta\���WD�d�*}���hEs��Iˑ�ċ�_�pKk��k	+����{�oJ��Hs�Q&¹P��Ե��u4�\z�m��@��H�U�����s�C�F�Vz!۪21�j9
����$r�)ߓ�q�v�K�p��d-Z��^t��E�}�b |?|�{���Δ�"�� ��Y���o�$ �D	�������`��\C_c��WaL������>�w����� ���L��uhV�=����NZ�?����pj���-��XPy�;(�0�2+�k��~ףl���vr���X��|Y�Fg�T`6����)4x�)M�U���\��	%�4��0�CA�D�O���X�2�ߘ�jI�t^-+��E�,�<}�Ҟ�#_��$;qC�
�%%{��b���dr�{$�HaS�!�/�sf�c��UNB�	Wa�y;Οf��ǰ� �fk��GM#��K��8��j��h�*���j�#U����^��F�54�$7%pYsV��"�s��~����5A�AĮ�D�c��D'h�q�e��\�Q�)`��h!�v�m@-��E6~V�,C,��nc�<pC���$��Lڳ�HL���]UNJ�3<LM�B�m�5��XU3;�F]��o�@�?�L�Cr���[���XѺ)�寤������(��0?UKB4�F��1��]�����4Fh�tȪJ�6䱎*�RܭR�1�������B�Z��9y�y�/Z���'�����¤�]K��#EPGB��j�z���.=��s|%�w-R���?�$8m�/1�}�KW��^Js`'����#K]���Q��TC3���v�7��܀;Q�m�9���u�����&�r;�-��ǽ�E�[����9�[�t��ZdgGM��[c��n���].69&��lE�F�����{Th��Q�;BǮ��_��TZr�Zq���p߱Uk��
�h�y`�����V������+�j����;ۅC����о���cW�>�n�P��X�����s]����g�{1佼�:�;���/=�Vx�agh�!�Gۻl�&�h�0,�=���_n���t\���'Z�}DpƗd��驵x������e�P�]�X_�o?z&\pJo��D�c����g3�F�(~k�풔�:GP�Cʟ�3�4ǟ�C�`Um�X�N�!�n�`컃�������{��Sm��R���J�r+�i��ؾD�	b���^��!Ϡ��a-V�}M,ۺ*]�EV�<'�r�_k��`�N��$AZJ��xǵ�.齒��ɛ���*��(�FJP���pZ�f:!,��M�k8��~����ht2oT#�ƧԪZ%h��� �rH��畷���v���|j�`d�Fκ]L/d<��z���_��~؞�������L�>d_Og{>� �^�p6��2�� |n=;ϛ@�>�\�����QK� ,j���<��§����'�˷Q�6bԉ[3�<6�� 50Bvx���Pr�L� ��_fz� �>�C�w%���޼����d��Ɂ��n�ѕ�-:#���
U����3��V�����<6V�x�#�7��s��o��ͳʞ��ھ����f���yB:�ɞN��\���u�Uyt�������5ȭ�䑷��tx���G���SL�n�5o=�8�"��r����옜�|?*�n$7�H����y�"��C��"Ԓ�	Ds
�:L��hf{�k�Z��ZYN%����gc`D���sh�:��T`i�L���LM�,������1=�q�����4����$5��7Z��K��������Z)��Z�N˿5���k�-3�O%Y�8������t�V�諷%�PxF���u�A��u�z���Pd�d[��昱,W����var����&U���(.�9C�T��`��)�|���t��Ov��+��"��J����*3�BM��'��r|��j��"��"��&��Z�X(D��޻�}p۳��:���Z'������qCT�/��tv�K�K8�p@p��ò� #b%�<�D)�As�i4��yY�1B��$�cZ�F��y؎�]\l:Z�l��tK��`�h5 x�-[uM m�FcOL- ��j@VCj�M�<
;��?6��ȢXU�� >o�� 7}����}�&��<���ra8�|`�+�-7OS+a{�Z���3>L�#���7EUo_�f�U�%4펣�H��"u9���iw�o� ��e��D��G}�#�fQ�^Fz�ǳ{�H�e�����Xwo���d�-/����D�Ɉ�(��u�Ly���1���*��Z�4�IKH����3`����4_�����u�����b{(s�.O`<�II>�,�sI�]u�N잕1W��\���'dn�=_��5�����w7 �n���P��5-�����ɤ��]P�?C�?��x8ޅI*��UqC����b��C��v3o	���l�V��4�*�&vB���e �|��Q�afБm������B]}��?dú�7�)�r���̌l6�Tƀ3G��m)X�ڰ����4S�Z��&=Lj�3(�kA�iZ��=���d>= ��@\�j& M-�q��F�@�#\��.l�S���z��>�X%��F�Bh��6p���ď��0��4�uվ�!Fk�͐��ـ:��<���Yĥ���8���Vֆ	�߳o*��ɊK�KE�)4�%{j��i���e�L���&����x^[	����8m=�]�,:7��0���um_`������T\U���m8�W6� U<��%Z���d���s�8�r	�cm\���\�\z��6�ɪD�B��']�m��X��a컗��sh���Z���*��4
r����oB�n�b���'�c`{�U�uo����� �3K�ґ������q=Hp���΃���bBRO`���&�N�u*�bՆ��f�/U&��<���%��S��%��`s�	���L]\���a��@�0s�!k;c�H�o�
X�{"ↁ �:V_&��u�uq�ǥJ�.�~�9ݨ`���V/\h���jꝬ��n�=&�_8�
�K����\���>z��!������2f���A��@�yS0.��q�j^����,�o]eu�T*>)�\����؎f��k+��ܥ�9	XzB0�FW�~ٙ^�^쟴o�њƅ��Ռ�B����a3UĥIy�c�i<V��^k�>Y�C���iZ���C�)u�\�)eB�0Ig[�l9���kh���A�M� �<[�Z3b�e���'�k���>���Tt�]W?��)�
��M�h,�$�,�Mk=�SG�U[�������&���4i�#�h�!����+֙���c]B�!�[m�Rf́	�<M!��3����<���������X$��U���m������͙H�Lh�Q]Ł{��qa+)��7��#S���'��ԡr�l@�P\%��YIh�=B�u�r��QU�:Z���4�;��ڜ�U���������E�#����X�����E��t~C,'��c%�c}L&lҀ����˞�Z�)T}�H2v��\N\
�섆����Of�Q�F��e��)gQ̋%��p"»o�nX=[J{d?��@��m1W mp{��0���wG˄�;�:{m9�^�rT3���$���^4R�e�F!�*"�Z�_5�b괼gGi�1|X�����5��#��We*_`C�5yL��p&�^�`�aS�婨�a�:��[��#8`�iAX\�Hm*B��F1�N�cu�V�H���y����?S/�.��EN���S�X)�`-�_�-G���f���}��$a�<�O��㼩�eߋY�.�$�	���F��_=�6�T]+z1״Kt+������!���v�S�>?�j�]m��48J�W0�
��L�f�.�¼� ��Xg
o3��I�b}�7{pL>­t�f
R72�iM� Fn��|ԉ�C,|<(��i�_Vq�T��q�Pٯ��\�'�}7m�u���e���A�@��䑧,"��1�/hz��p��ʄ�mCJ�Z��B}��kd&2T<	0ɖ�@Ϸ�-��`��U�v���x� ���
�""c��] �]r�/�k��Ŵ%t.u��x���������/t�cf��´"a�/��7��9e;G�:ıY�Y֣)[��T�X����8��QU���?��fT����Y��ЋwOG�,{��q�h#[憺o��zb���Dgi[ ߙ�����,r�a'��.�M�y��I!��X�nq���]T�6)����[�`��O�WD����@uu����&�{tf���>�s4�u{�����U���+ΐE���7?�F�L�����ݦb����W�7[�f)�B]�]W���x+9�uE��vJS�ۭ�n�2
k�ŉ����`}3�ܔ0�B��;gN���F����FP���^>���G~CO�t$2ɾ��A`��F�7Vw�<��<���umW����9%e2���3���_�%'��aƿ�i��w�*����`��������A|`���[��F���H@Ig��z$j]Z�҈���{c}>P��
�r �Le\��`�]�U��dz!���+s�Ϙ�{��ow|[�˫���=}�k>����Y�ia��eJb��@�`\������a��7bK�sp>B �/�g��ϖ�Eqt���&W�^r�)U�>Տ+2���-W���mpB6Cd�R���5���$�⤬���Y���ڷ̟j���i�t�Kh�	3ξ}8�e��"��;	�9ة�Q��JR~���e��D�<�L]�`�����;6�?~ۿ�_O�y��#S�ɏ��7�G��2&G7Gǣ��.����62��Ql���1��T��_�L����}���K�~[�����!��l�j��"Փ�(	�u����!�~�Vwl*'d��)9Y{�!�}ni��X��4�i�~���"�i��W��x�cv�Da��ެ�d�&�1�l�W
G�>'F��wQ.�,Gb)Tc���-�O�I ��(�G׈��e���ʳ��U�6���p_Їӵ6IV�r�@ui�v����+_�8*���T=;�8��t{ߚ��/�!������:L�3��r椹�d��:�%�P�S�#��Z��zK�C/��֚yz-���?a"99�Zj��Ĥk�����\+f>F�LjT�U:��6r0��@ԃ����`�G�E������n"��άq��\H+��)%���st3_{q�7@r`�'��o�� �+]/���B��`7@��X0/m�YtD/)��U��V �dF�(�=��=�v���A���7��y��ıY�g}�1�v1*{����Ɩ��&"(�7��B��\Fn��G�Q�q+h�P��5���'��:IL���é>��ƕe��`ȸ��K�pp�%P��AO������2E����VW�~��_6XT�~I*
��p�Y�b���Ҿ^w��$�8�,R&Tݘ����u�7�:$a$pJ�R������r����%��MZ.N�����$i��-��<�g�)��������Sz��6�Bt��i�����\u�-��IY}��7��)a�~��2-/t�E-�}е;|��;v��u��N��}l�}�_��{5S8~r%��N
7���4ə\�f���x�Y4`��}vy?����$���r���~*���	{��%]uIj4P�V�<2�zTuÂ��d���ȋ�t��Y��͞��l��!��������)�������ƹ$��	O>�.{�F�`�sH��]p�#D�ڼ�v��h��ı��r�ok;�cɄ�Uj��l~i>=3����8U%�fC������#��B�í�m�f��T+������������źD���,�i,��!u��oxi��h�<���p�,�uͭ���7Z����T_��?O��r����� �c��x�1�(��E�}D�>�bωf�e	t�E�������<1iԚ<p���<�"�*�UNW����_���n��#��qM'���>��4]���%554�R���<`�c�0J>ڦ���go$5$�`&�Z���Ӛ;�{)��5!�E�,��"�n�Z�+�x�lc	�P�'R1�V�)C%������!�����~��7m��2������U�w�n�=�ʊ�	�r�<+�ϴإ�����do����8�"1~W���T@_T)�l��e
��������Q�Ľ��+��s�|Ķ��L��5��IK���w�����]0�M�_��9��ё�&/,��>�|*T\kK�ވ���T���x#U6gxYo����[GH�4�Զ�%��A
�nf����(�Rf̐+-a�X����3x�jC���3Xh�TN!����u��?�F����+	�La�)�
���9�.���NS\�t��39~u�a�Y�(Q�32!�ڍ�Gg���Np� S�Hcd�bG��ͩu\2��G��Xo��î2��V�:*��J^�Lfk�Hf�)���-kUs�yL��nE�u�-���"+����J�����������g��Ѷ$�PW� 
�t�C�����<H�dO��;\�t=�mF�	�����PXh/��Zdp|���6鶵�pA������B����	Hƹ��i��s�lM̌94	i\ͳ��2~�	�:.@����͍#nX��t�^]��6,�d�8�OJ�mg�K,���V�T�.��;6��\�.D�1F�|��C,���쪇�VuA�|ߘG��_x�͹Y r*M�O8�a�%U0`�7�}51�b�)���1�HA�Q�Up�8��Щ���)���˥��ؽg;��q��SＮ��Ē"v�ro�c�fQ�x�����3���[*��y+ ��D[E�+�f��/;���H+�x^Қ6���v� ��!FrT�auhQ���|9��:�e�
�$�GAP�74`�Sp-Uw�O�/҂��P9�u��wbn���A
!y��KjD�,��Ɉ��o������h�e���F���Y��C��n �^�E~B�P���$Ru��{���q*L��OƘ���<���R�J�HrO�4��=����ռ �`i�h!+^�Xz_�<6� �13�1�C��C���^ە�ʬ��2M��A�~�QhL�ˡv��;���U7��v<�we����~BF]�B$�'��3�KJ8~��PD�����,&�ی�`��d����4.��2�0gm��瞳�H��S���5�v:an[�&�?b��B.h+	 ^�t`ʽ�=�^ڭF�yJu��Ep��"�#�Ao�)�BbE�l�Z~�/����^��~nȖ��uOڴ�o�J�?�XГ3�͘?ث}Š��XBN���,���ᩲ���b�pmb&\�Fp���Zo�I�Ζ⾩��|�RBF����R�Uا��R�>�<��N�S�ż�f��=Ěx�fY=rDu�����JA�Q%�(�WE8��z�XD�L����q��9A���D��qj6�e����pG����wo�=�����{!p-��-���R7x�V�W�4ͯ*�)>o� E*�qG	�1U$����h������N�4d�v�n�[�&������J4���KtO�x����y�?�X��A���Q��9gj�j���4��c��"�*3`��3�zI����n��D�GDp[1�	PRKt,߆Ug���|��U�)�q�_��$
@����]F'�!��#���U9d�E��V����Q��F�wB|y�/wl�K\=��F�G�o�4�c��qn��M�N��7e��t�m��	k>4\��R2�)���@�����t�i�jW&�cv���`#��c��E��)CU2��ǂ3"�+�j(��,����o6�O�0!�^���lB`^L�����s�߃�^_���J092O�k���Y�f�&�G�K�)4�I"��Q�!�����C����>1�,+��_�d�_7e���&��#F��ﬄ�_t��$Q��V�sΦ��M�A� 
hhЩ�`��V~�rA>���]���O:Q�1M�
�����y��bл�pucO�&;kR2��#�����*E�\Ng"%+9�:�F�}��U��8��)GAZk������H´�!U�d��r�D��?M��08��r�E^��Tb֓�5��F!������N�7Z%[B甅 6��<�bf"�M����$� HD��kY��T���"����E��p�%��믣�=J��e�{5����m���H�F�@�TV��&����H��a�*MsPW�Q/���'=�̶�_~,
�A�=��5ʬ��z0�!�xA��c��*�$$�^c��;�ܛX�J�H��T��_(_f'������`:���A[�hϹ`�^k(�!gM=�g�����Ӿ�\�1��^��P.;�
�΋T}���-�d���7�ٮꡚz�d�T��1#<x�N��6��^s�iD����XP�$(��<���;���u�MO(��7��{]O�}u�)G��΀�֪<�A�L�#��B�ԏ�uO{�#[��hʚq.��XjC�9���/�z{���n�g���hE�J��=�U���ɨU_0�xbtJpD-�b~�M�@�4�1Q/�N��G��@>�N��UƼn0�9���j����Z�ѻ����/�j�)$.7 2��ÿ�1OWT�2� �-k���OP��;p�+N��i7Jo��/[g��＠���v@��9��ձ�WD��k ����&x˾�;�%|�ґ��]�O"�D3���(ঁ#�)j��vSG:-��;ha�œ�!E53pL��H��ϴz�F�G3
Ik�3�3�k�rB�׻������93>l�\Q'KYWV���i]�&S�0��,��z�t��{�>I���\h"�0�	}?�'vҎ�G���7��n}������Ku��9��=��"&V�|�T�/)��;,�܇ϰ�}�ïO��x假΄�����ĹgW�/?�F�YAy�?�����䣏�H3�W�0R����*yab_ �����S@���YS%&ݟ�J����R6�����o��b�CN�p��������d�Z��Qi~���b�U ��)eP�L�:�S߷z�\>�䋘ݕG5A���V�߇�S��n��u3����)O�o�c��i��q�%�;�y#;���C����V,��t?9x)P�`8"��v��/[�`����i���ӎr���������`<�X�?���C��ch�o]|8�?�W�Rm�|d��,f�s���v�5����*e���BqrEɴ�v��JK����
��
�8�#���ߵ���y������������R�)�^��#7�0j���J����Fk�X��%^����VM�/���`�B��e��w5/r�3!�e\*"���1�g������@��.O�AyӈV���Ǥ�L�����M`�0qi�S���o��w)�Ȑf�/��c��m�2���MlW<P2>P�uH�8�N�#*�_� ��Հ�[ZL�ӌ7��d���B�>��9��e�A'F&@4^�D�g3y����!G��Za�;�l��1�_�>��U�LkL@z,�63;����E��6f�M?K�)( ���}h�D��e{s��[<��@h����m��Q�}^Xlp����0âSe�K�S0$��>�$�E-���>�xÇ��)�{�i�G���U���5��ͼx�?L̋���M�ā����-D����y9��"j�[F���X���*h�����5)h���(Bぜ��/+r�m ����ˤ VY܆�ل}��P�����Ñ��O�ZLs�;���,ٍ��G�����Fk5AWA<~��%����`K8B�z�Y.X|�*��]``�s��aX�Pe�,ubO[R~����Su*�r>�
�H�����*34�b=�y�Y�6*1��N���_;|u�vE��c�6�<3cO}�y��&M6h:�(u�]���"|����@���B~���ae;Hz�#�@��<Y�*q�y��m�6k^?���~:��\�L�����'�\��p������s�m�����e��r��B��s��C���~ﮀ�|�:F�o-��:�	��r,�`%Qܞc���bĶM�@��z>x���&�nʠ���ٜF�?��th���vt��2���1gW#w<�M8g}����?t�5%���R�Ư�.�t�7�p�j�J���cI��2�����7vF��&8�Q,���'jf�=<�������Z��>����(lb��~�G�z䲈rL�v�`$�,Lj�I�`.=\�8�M&��jM"�?{ăv�/I78�pm���pbҕ�嗼���PL;hm����-�f�%+j!�>��ݖ�&�~l7vF�C{��W��#��${�b�]'ip��������}���0�F\�r-^�-�vZ���XlU�1k�T{�aU�9]"n��O�F]���A��V*z�e�r�[��5�S]N��L�V�i�&iϪ��]��GWbi3y�N���N���c^�
�����h=ӌ�ҋ����w+��OI���3���+0I���~�r��/k�p}ra�����?<ɝ�}���ץZ��G��	eeB�����y9��G�]���b3��RIi��d��=zo��+{=?��(͸�V�xg�SFv�{X˳�$œ���W�R����Uq��`��e�-�Ì�:����M���v��BGՋ{�4v��r7q������<�m�N�grЧ�ͮn��^8:KQqD?��1&���[��3�!�ާfCz����4�(	NB��s�2��+��5MH��1NF�ցb2�&���>�'��S� N�J�xŧ�WF?#@k��f�L3��f�3ڣ}���0���ou�}v��0uV��35�L���(�ЦO�Ĝ5����Ā@㽋 �Vf��Ql�	(�PRN7�Çm�.F;��3U��w�dT����6��O͉ �6~�nV�OT�,؏+�'ɵ�Ӱ'T��K͛�=�@ ?]��u��Pku½4���'o����w+��}�Kg�(l`3p������kZ2���O[��n�}��[�I����1֜>"Kec�:�������^��H.:*0�f���ބn��ġ��ڔw���%�e�=CO�;;��
i�A�c���H I{J5��A�nx�J��:�r�R���<�:��d�n�g�kMd�9���B��Vp��3��< I�Od ��Uy�����.��7�n35��b~��^C���t?�8��*hQ��r�=-7�Z�� ���-��5mQ��<��(Q��+洄E��Y����3ۧM�����(#�C������V�zaa�P@��E���J���)4�:�ZO�2\�J~�]�l��sM6����Q�;:�~\V?R\pdO�J��=OR:0,��;�EIh�T�字�G���w����읣��f��RwB*�2�{����7��Y��OB� l���`Î��d�,�ڥk�^�p�	N�o��������q�ހqZ���v�Y�<l��^r�=%��u>��#&K���Q�nH�{/������l�Qd�S.kr�&�v:�!B����2S������u)E��DA�6�N��fיh�E0I\���u��vqohIjc�.!i6��]�$�����cs�{3��*=?��;&�%R\sBPc�͔�u�h��4���6��4j����p%�.�,���-h����"�b{�e��ܘX�UZ\���IF�k�}�����ޕD�uy����5l�� p\(�\zvp�`�ݼ���3��%.|�K��f��!�H�s�dY�# ��n�M�δ�,�뾗���&Q���>����Z2�F.�a�ޢ�AC���pX��}x>	��=|c��t�d�Z�SJ@N�׉����d��C��A�S�����8���4���&B۴$+�M �J����CS�D�}J�!	����[n����HH�����zGw-YGv�����w$������)����%�.#φ�T!��>���(��`��AL����ygl/�t"��>dXL����_�J���8�]��yI`�G�LH���DH,=��4�U.?���bԶ���[ޥܷ����=b�>�Ė�w��o�|pax��l���9��a���[�}��H.1i̲� ��S�,�Φ�_�?/�6��6K
���n��=]�YѲ5��3|�d�А��DQj�;734E��@k�G�|�ďkv��v�(�z�߃��o��-���+�"�#��c�j�í��/9PV�!�+��῁��Q^9:�h����3�es�q�t����ɐ� {�z���j�4=ǖh���C���is��]��cM~r��y��ѐN0��ʾ�ˉ�rdx���d�����
H�؈5~��Fk����ȋ�I�EO|5(b+�8(�-��?�-]�2�)�#H؎rs�M]�j�]מ�|1
����ϛ6����B?�~,(���Ʒ�C��R©�<�Tӹ8��;|�og�����`��m�!q�$��⩼tz�~I�ZFRlln�k��3FH��Ca�&"�!���;�Xh�

W���3%K�#In'r�OV��J���X1�.��8��!ً.�Q������G�Tq�b���<&�7_R��������!��M9M����:���L�<G�' ���WP:iȤ�u�N;�	��˵˧����n�jD�|��Y.4�f�Y���J
4��vdu��|�UᥩgY�2����U�"e*�dFG�����p&v�,٣N��jHp��R����*S�	��'�����Zf�9��I8�B���	�U��c�B�(�d�1�qx��gn�Yy�����Y+:J�&�.!��y�O���*��D�q���WȌ*��F7Q�hF/��㛯�l;o����g�1���d?R}���D������4vQ�g̨�KX�#����	�q����w�o��נ�VjhҶn�s�*�_�K���!d����r��Z2�qՏ�!�����U�`%�9�Ð��J���D�Q���?^�o˓T��gx��}�I:�O�)�X���������i_8)?���Vu�6�����X���_�B���r ^j탈�?f��}%��!��\nEV`a�ec��C�f�_��D���܃���ir��caya��9�Aŗ��� ⺋9�r��Rң9�m&�\U�Ǎ'�u����U6;��^���/�R�ф�px�?��~f2�Y�H�H,)�q��Ҙ����a�OEW֦Hd(.gX<��Պ[_Y�?�<��J�� �ƫ�"���:��+!a$��3��8��9�*3�}d�{��ņ] ���p����/��=�s���4������;�jr�	�{��仃8DH(����v]���yoKB\���hE��y��������ʗ8F 7q��L��U���Lm���م��͹��r���>F�u�< U2�( ��w�m�^����ڭ�/w"0�M�K��=���O�����6�(o�T�1 �F7t_p�;R�F��bxh}������)��Y���!Q?�*ƕ���w��'K��� �n��Q���rO)١����X ��P�_����!�=&�UI����k�3���
�T�����hKp�Ķ�d�QQ-��ׂ)���3��	�)�p#Q�$Բ����9�,��K�"���udͽ�P��d}���4�:��{d+�(�RF��ź��w��N E�=B
�q�\�v�_��;�r
1�ާ���p�����t�yxU�f�!i���8t I��񠔊/���d�.#k^[5sF�m��ҁJ�fK�}Z�/�N�(^������m�(ؓm�_�h����
Ưz)D.Ng@�Tc^���2�Pӯ�RTt�`�E���� ��3�q�~񻇲����yn�s�G�\���0����O��������LV7�N����\��S�ڮU��v?���5��}&2U�1�`�F���]c+]=�O�5`���k���o2�g�
;o&t�I����A��)V�+���`T$~�#	i��6e��fv�d�-�[J�K3����-���س�ץ�����PUD�&%����}J�$ "�.���-#V�1YHMc$��U������Noĵ���k�l�:�<OIxS0� 	[G���r�⺵-����q����k�4���m:;�X;�X�R�&�YYn�g\�gm?C?9ě��Fk�G_Kt�T��ɉ��\Π�c�q�()���VWI)/T1`n:�iU�A��.#;�(��2���l�n�;8S�v��/������S�+�rK�v��k�p�2�d�m�)8�rw_�s�0D�3��z���vi��x��z}Y���̻� V��4�_�wS2v��+))(�q����-�kPE�Z�q���x��_�L�f�ռ~��.x�]�}����_�o��EW�nVb~����=ˡ�m�\��g�\3�_W�
��Ƕ��},e/�Q�r�m�:�B�m�K�l����kt�%��l��?��GZ�۹����&�p�(�c�ެR���'�n�љ�=��)F9�w	�Cyn+B[`Q�|�ݭ����O���E��kT�+�`2U�3�Ƌ�l�'<��Q�T_�R��N	O����g�7ڃ�s,xO`n�2�	ɳ1��H95laU��n RlN�����#�h��0.�d��y$Ӧ������j1�d��@<<��6��τ�V�Meە��]���o��W.�q ce�����S��]�w�C���`�#�M���%Ϻ�+�b�KL@�>��Z�ϓf�����2����)�Zx�h�n?�A��`�n}�kl�}�[�Ͽ���\��}�a�1�WT�Z���v{lv�js�����X��m��m�b J���ƟX�F`9�C���OG��	���o&�L�O$���A�[��Ø�6��ˠ!��Mh� �Q��z%��w���!�#݈	����Z��}�	��&Af$�oK=���9��w�`3]�:pM���u�[ �d��ɮ�������Bz�~#�/a�Fh�����2~��`���<P���3���T����ʢ�����!5Ό�U�ۯV��^::fZ�9�n)b!ʎW�-�j,��{�� l�e�M�瞀5�5x��=�<���?�5n�����	��G	-g��u�8sN��mU�Q ���( �hY=8�c�t��`��ifpk��w񛡬���vg�4�+�JEꄋD���<)YAj0|��[��C9�S�����p� 	{F#N�`q[j{Ӣyx��%�I7H��Af�ԁ�O$���/����U�Y��L*��	!d�X�x]A��h7/┨tK�h9����\b�9YPu�����@�.>�/A���)SF�Ki�M�VF���'��+uI=�b:����К�=@��/1u�1Ef/��}"G1o���-�I����6wԻj�T����<�LT��k��D@�_P��v��1��k�~N�P]y����Ɩ2��&�ɏ���⨄5Ӗ�K�X_`�u�y�_ˁE'ټ9���fU�K9�p�[�c�jl�3=U^'������)�M5��K� �x�Z��|!�'(�>�� ��s�go�b;���:>�K�4�pl�+d<룅��r'����X������-cH=�|e��G���;mđ��yG����IrGD��O�f����W��}3�vU``B!�]�? ��p�@�[��*��ģ�_��X`�v�<���9~���3��(3���&R���MqY~͂W*jw�����~r��{���v�O��B�#y�ɶ��;���k���1�.Fh&�R�҃"�s�%'S�ו��v���>���00خ���s~=t���#��o��,*n������
���Y�)��m&Y�M�u�u���/����+�^�Yt�g"�Ճ0��@u�	F�HtcZD����0�Y:��c��4�G2��H�8�E	q��2�K#Do�̌kԥ!8�N�xb�����5n0�6@+�)�Q��`� ?������2�%��ڢ$i�`C��`�{���c��Pk鲙�G,S������v-_�LF:�n�5*q�i%��3�,� b�m&ZccJ��~r���3��i�܁�w!��$������t�j�/�Sx�i��J�e3`+��j���$��5u���7�3�n�Gu���vTf����	����?aݦ��Rs�+�q\U�g�Tlg������'H:��V! ��ބ��.���@���k�u�ꆖyw������ѩc���y�UK}1������,�������i�%�'�p���čGp�Ij���c�rQ��T�g���d����^����^.�C���c������SP�Lǚ���k�'#��"�C:�+j�!�� `�`�K]F���k�CƸ�Ճ�qa�O%p�%؜�tю
�l���~�e{�;X)�%�7i��h�OU�W��m�$ �	��ʪR��<�Iш��)�A�������8��)��L�����H'��|�)g�
�sUI�+�r��""�?ٗ=fG�r��m�1.,���SQ�\��姲p��h�D��	���UV��pwgs���%���H�ޅ8�&��$�@d�����0���5��0WY���7��mhɪ�y�����¯!R�(I��{�_���7�"?�Jf�?�Y�)<=k^�y���U�<e�!f��绤�_��,Ğ�lbk�����Y a�̒.-%@	���GB. Q��_�b�&(��&ƶ:P<b��GC���	*q��łh�,��\7I�AD���������_���B��V��X�)j�=��x� �ގF�2o`���D��A �eXO5N"��n�k�_5�|��h}Kے�jT��^�k��4�Ȏm\���{&��{lq�Aiu����?�>@���κ�Z^�P��
)��ĸQ�4o	3�����\\�(4�A��*��o���ɿɹ�7f)N�6�XC6�35XI��9�%������RXs:��LZ���'�Gk��I1��ŭ:51�d��S��a��P�:[�\�ŭ��)O��heu��1�t_�f���_B �X�X����=��Nw|�k��@,�U��b�`AA� "l@���6GV���ؑ����x��+��O���*�օ���m"���
� �Yǖ՟%�)��e�lV�ڀ� W��U|��y�@��'s0�!"}���{iį��`�ҫuk�z�,�}�+Sɽ%z/�����������<d����-����Ю��D	G�Ԫ���\�p-44�1���Z}�XT���?k f��,���lGIɔ�=�0&�SW����mq�#�+��nva�ļ��ӽ�)<:� t��D����ym�D([(�Ҿt�E�2��.9>�j�⍆	�V��z4��F����0TD)
����5��h��{�W�pQ(��T|�S����=9��G'g��0]3�ӓ��iE�ܺ�w���<eX��UwJ���B'-�MƝA���&~<)
�v��q@8�i62[A���Y��"
+��
�Jd����r�0X�N��n��X�9J�r'hWo �u�7|��6v��r0*V���f��G��F�,�턽�}vX�$��9��E`2w"���e�W�ѭ�m;Al(
��x%�a5ɚ��ȕ�{���K- \]����)B�S����羿p&�.i^T��+o��lG���
g�������}�0*�"�WJ@���~��R!��
Q�ַۥش�U�ت�ɏ�hz��;򙅐8�F�-x��O�G�����y�Qrvѭ;E����k��&��vZB<��Xs�5t��y3����X��`A����!�G+�׸O��OU���4��B�w�O�!��ܰ�>���L��3��FW���0���[x�}�k���%vC'H8w�מ|�t�+֏-�/ld��4Sa^�M�̔%��9��@\���`<�:ͽL(���cՈ��e8I��Cp{�H7���%PO�-
�C��_mdP �5�MGkB��u�լ'j;p���e����<������tUc�(V7��ʿs������j��-|\4q?�b��<�ěĕٷ�p�0�C��K7]������#��Ahk@�7����T�!Mk��A,�f34��\�k�v!*r�3���D;3ū'��⋙���kӫ,Aw�N�������:PG����s�;A��'
��-4Ͷ��I���F�.��^JFV��U�1��
�A.3���0��#"�����@%�J���;��]�AVկX��P�ա?i�f�����H�i�����O�~��Qŋx9/9� �f�;���f<�7���X�Z�R�>�u�J:;��S��ل����w׺6��X�������������;��Һ.q|S��uoƥN���(m���ke�����<S7w��pS�(�L�d>c��n��W����+��L�7s���XGX�&�+�官��VO��:x����yp�����iE���_�tx�_I~����j���Z�QR�M�d�.2��$����y#E9E�WJݏ+�G*,�N� ���6L�Г����ܡ��3��cZp�����Sʻ ��ܝ��De�������8�U�ꛧ��"��v��ک���  2������q������߫#[4�AʅeN�����i��Eh��ᆦ�E��ٚw&��3�F#�|-�	�.�ٱ�bуr�ݤ������w��»L4�Fގ�u.itFd�
���VϺ"�����%�=�Ö\�-&��ۭZ4���8����X4�/pL��oT��L�Pj�|K?��M�Fx�w�BWgi�ݓ�h�D�H���j�|����B�z��dȱ�]��T.��J���S��%�ŵ�՜��{T��ȯ~u5��7�sˎl~��pƁ��HJ�1w�V҆ �մac�B����wQ*�'A��I���;����~������k��ʛ.����� �ۊ�c����b�=Y�|\���ڊvk(�E�RX�AVn�4W3i%�����zJ�i�6���Ǥ���%d���6иrx��G�Bi�o��z!��Ͷ�)�]��L��n���ݫ�x:�71X�dۯ�˂'U�L�qS�،5���D�s��Q�\��g!�.�-S�b���u>/������w,�8���d��_��A7TMO�d��'>�#*�I}/���5nI��H�Ռ%"�+��#X��W��Lb���뾪`.���Pg$� ��<`���ϲ5��\���n}����z8S��7��T�cؐ��tR5RP������j��;'Tt��� O�usr&��j��:�m��C��`6&}=mQu�}�;@M��S�W
;����am:L����o�9���P���<2-i�@|�w�̺�:����f^`<�T!�7��3x᮹7X�ـv�'sq]麆�qf���FkW��9p����w���_&��7��'���B@��k�}+N�S��C�O؏I�I`ŭ��/S.���$�� |��h�^�֙�</gǦGc���6!�s;�N�~��,�d���>%3�K.*(�y�w�3~Z(���>�S���-1�a��@Iu;���kz��l�2��\`2���`��!�����")�W�������6��[��MP�����ܫ��z+0���&ϭ�%πFi�"b OO�1�����Y�ZGڕ��-s[��6ϊׂ@9��a����geA�z4\0�e/�u�6��dL;�����Wx\=���LڄM{QI�i�3#�Y�_k}Ro���>c֛E�L����x���66F:�9R@��(h�#L@t�A����f0�����|6DK���������2�_,����"�Mc��a�@O�d&u���2*�X&.�'9�K�U��N���>��r���Z�
�W�A��|�Ur�21ջ&�E4>��2�K���(�(qU�����i;1*�B4�^ �p�ʕ�y��������wN;>6{�>��1y�d�����o�J<��L"���u3&t���.���T�fX	%�ؠ��I�r��h4m3��K������׶�I�)]���s>�y�1tٹ���%I���9o�Ә�nF�T�62��v<�|��0"��V��4�q����θw�H�5Z:
���ǅ_��g�DqM��Bɩ~�<���`����ϒ�6�e�R���;%��!k3�vOOC�+�n�?��R����KQ��
�ҿ=x�P���F߰�sXuڊ�&2-<�����2�m���	�>��]���'j:'�Z�Q��$r�?B��qnFμj44�Y�^����������0ӷI4Y�{��A[;{l4f<ele	�q3ӱ��)ܪ�ن�o��1�ey5�nX�������y?Y�U��/�a�$H��ʔO�w�2M������"C�i�j%��q�_��:Ė��6:e��rw����ɰ��I�7|=T�,���a_�( h)۱��1��}(OT�-#c�q]�&ȱ�˵(��.�9$�Ie�-|�f{ʻ��m�ީ�>��L�	���K�u����z��#�R�3�sL�S�T`��_��;u5�~zZ�ܮ% 5$'��S�TAY��!|��t>M��nE���xB�r&{�n�~ơ"C�Y�)/����;��xXJ�C��p���6h�.
_�c�T&qr_�DozWJ�U/ �!�d.��ܣgvxc�!�Xb0t�:0;��r�i/.���UД5WrIz���|~�y�=ٱ�r��[�`3�,�}��(��kH.A����W�&)�j<k'����:#�S������B�b\�ͤ9�H�����.���Y����HQ����2�8�ゼ���zM|R�ߞ��[���06m�vƌ����>�x�����9!�1�2`��_�gUr'N#��o��O�	��[|5�k>_yBqk�/~m=]Z���X ˂kD��s��7����t�s ϐ��,�_}�l���e������ѱ�Yw�^ҪĊ�=R�Ҥ˘�	|wi��oL��	�b�l,��e�S!�<:gqQ��U�GN����H���3T��?t���R��s��=�CA�!�O��\K�*��^�Ĝ�G��x,eœN��D�[�\�Q���~\Q��$�C5��+�!k���`ɝ���i�FJ��~wx�: �"y�G�a�l��&7���¨{/��O�;�Ql��^D�:�g��8W�����X/]Sd��av���p ��ãD7N��U
j���6�"�{�k���u��?)`��n�$n�O���B\9c�4X*,��P�=���q�n#@�Mf�6nY�����
��-��řj�D<��������M5pA�B��Tr� x���#��ك�0���.�]]��Qv��xm��ӗ"*e�(_[� �
k_J,d!�6�3��")��&O3�ein�ʩК�Gq;�8��(<>²�wbK���,c��(�W5/J����*.��}q-L[�+�_�K�'/�P�OMs�I}W�y��/:�e��&ASo��SIL6��{;�gf�!Y�܁ں�q�$5���`֥@J�9]���R_|HG���K%nY�)�;��'w�f��ҳ���\�u	5��zX(�gG�'H�h7��{����-NRI���=8p��ld,���:]�A����1/����L�ZW
���^���,9i��J���b\�" �_�J�����2���<
��6�_ܑ<z�Me��S�@QU��(�$����^�'��������J�ڸ�߰U�\q���t=�&\9�7�KcSnzr|	�&Q��ĝ%���4��M?���xx�j�d��G��	�_�ض�Ք��W�|����	c*ԥ
|½������
l	��/��x����tǼ�m@C�
N�d�S8!�7;yo�L,��-8�ϩD��=�J�nP.��6f�󶏡�(�#wi._���O1B�>��9N��H�<B݄��$�p��v���@||�J����eӭ�� ���}�~�c�su��n&	��\; ���M����+k��'�h�]t1d�W#_�!�!�0M#{���y�^��&�]����>k����BԽ+mZ��|H�op ��@e��>�^ C�U1����Ȭ��&�4�@�|�}�u��-y�U	~Bt��#_@	!9�\B���<y�3�y���{�x/�#g�uA�`������+Q�(ޟ��+�6YA�J������Ƒ/�I��A9���56���vh��GS�����m�n8���,���n���V=��t�T �]�?���Pr/��VU��U�/�#�C�'r�=�����
ἫgXqX��[V);���xWt��֯E��XY;���U�{ȋ��*vs�,=�e�ǩ��>`}ZNȄ���m����88�wz�`fB\T͕�n��Q��G�� ��/%�5��^֢���.pf��ؿ�x%Az�&��W(s�щW,�<8�X�h�]߈������-9L�����N�D��}�b�#-����L^Y��1d�]����E��g^�u��B�έɸo��Z�I�0r����u����ۤ��*��T��K�=�'��w�u�a��n���rC�����r�!,� ��|�WS�?��z��̕C;�x
�sӝ���TB�4�
�t�ǰ L��ax"��{����!=g�$C�! �|2@B��#���B��Qb�f��v;�J���ͫb�đJ����מ�ey�X�6���0��s��V:;�+^ibd��W���~?*��A�<��T�.���3��v�n^R���H�m�-?�ж��T~P�o�.�i63�����S~�\��f"�?�Ѱ�N�8�c�+��P�i��q=s\h�XTG�B�@��i��:%�<��pU=d~�*?�K���Ӥ����e����U�e����{���-Y=��;y�w�u�J��DVRq�V�A��R�'a�Z/�G���=�3;l.{��b�� T���r�4A���'V\' �&�i0�Q��K��Q�3�ӣ�u�qg��m�^���y�aq�+0�����q:� ���+~}G�I,Lȵ�â��7<�P���!2N��_����p�۞�H�&����P�h�9l�[C�&ѵ�*ɬ_|_�;���G&�Ez�!�@�i�ո�&_/�V��Z�o6��ם�C�p�Pv����ώ�U��ޒ#�&D��߄u68Z(1
{��
����^6��Ά�V��(�YJ���w�9�	���ni��<�Hn_k�B���MF�6yB�8�o��P�Ix1�iǎ�ko!h˘�t���8�@�@��4LK��$p�5�GQ��hǬ�QD�B�@Z,�w��c�� �7�L��'�������@�8I���`�'Ay�G�իX�a��R�s���鼮�Q	_%&����wSc��P�e�
����x�H��W;c 픪��Zl�2L8X�2�J8�2h>��핂$�t��D�\��ވg��s��4]�_�JXd�������n��,N�yR��MoU�Z�*m���P� -�8��/	r��)p��s��Œ2����G�X��ȧ^��w�b�&E2�,�,m|��M(���kY�O�0Ci�(��\�t�R������D.�L�y�&D},��$�f.pi<>ᇤ�-���e|[�z���ǯ�-�����q\����&84�u)Upu�Ey	����T������`x&�υ�2��٠�(�흲`�.jcr�J˦��F?j4C��K�\(ciӖ�	���?�K_;���Ik@���xv����?~���+i-%}~�qh����U�O�0�b�ߑ�؅ҡC�ѐD$���"Q:���R֧:boc,��v���o)��w���ї�~A�YP+�(��_M^U=~�����#�	��3a�Ͷc��؅W�4��:>k�qw7�I����Q!<�^��*��_���5��hXo�us{.��]��YG�&8,!���鞧F�d�t��N��T||�!E���!�)�Ӛ]'�gQ�6N0�����]�6��
������=�[�/�_4���8��<]t���㴧q���-(�ݱ����ZϪ���'�-������?�5����s]���h�������x�u(�v*0q�"����ܻ_�Pd�s��������5Z���U��2�k`����?G~�����Ñ���qN���2��$I�,	���}f,L졚[�\�fLB,X���i����s���F �]���A�w���Y��W tʧ0��Wh����f�Y�ZyU��#R��0�0W1I��Kb� Z� �h�'�P9�S�`:*���(0fӅ�Z6n��e:� 3��tjJj�V]�Ӈ�m�k�ʍ}h$�"�� 훵���G錭v<���BVظ��9e���#b}����ꗶT^	c�h{=�QSɶ�κ����`��v���˖6IKʯ�Z;3�/���=�D4�xm2c[~�rP0xdcA ��D a~�G;�Gd�E�U?��|_=������Q��|�y]`��}�Uמ���j<kG�xln�'��d�Y}(w�����D2l����ȴ�dW���6���g+�G��XkQ>E�w�Q���܄�<Q�\��K�2\0�!�WjO�k߬(;����0kЭ?d��U��r�(��p_" �}E\��jf� �"��I�v���8Q�dI�,;~07��r�z�7;\�x�Z#��%�f/�g�J�t	���32q�H%�$�b�'����|�\S?0��o��{dH�7����O�H8u�%����f�<�A�땛f�C%�0���+�d�бb�����fR3 ��
��ɋ,@�΂˶����-*��1�k��
�ad����"�z�Q�к�,��D?L$��0&Ր�.��[������*Q��],�Z	�{P �;d����P%T~ѵ+�����
F�J��1�p5awh�Y���@�r���np���A��4�����h�9�P���� 1���v~�<::�f��k�F�11����G(���ҿI����fYV��*�P 92���k��#�ͣ�N�sZ)��#�wM��'�&6Y61�]��5������l��׉����n��y�X7Nrj�,/E���Ka�(.���R�p:.�J\��Mt��h�����?�OtM�.′��g9QLϳ&9ޟf��i��������=вW��6pX�J�1�.w_�:�=#X�������n�te`w^J'�M%�$���G'"���Y�F�z�j���$b�;�6�\�T:�H���lz��s�x6T��	�'�D�,*fr����3��4"$��"U�g*��J�ޥ�K}UD/��G�S��w����އV��|�*��+��h�F�J� j�����#J����#[�p�)7UJ�|dWw�a;���8� �X�x�*�0)�7:gu��E���LB69�7D�iz�Y0@�r�C�5l�n<��#���P�.<�zQ����4��z�44EQZ@'"�D}.y�p��}�����7���5�橘���޲+�k���T�R�nh����7�:���{���Ԁ�s����)_�3���*t�g�	�*���w��p�m�dH��T�5�~�0�~�F?�ߪ�u�s\<!�M����b�'����+uf��3	c�r�Ѣ;� ˞Ryu�-���Ĝ ��=�Z\K�^�� ]���׹��X�/���B�~X�[�2C���n��N�,_in�._��x���c�luZ����F�ĺ5��ֆ�f�C���!B�ˇ����$?`�s3�:�i ��զh\-l�Ü/���(�ۢb�]/ۡ�g˦�Zm�c��$���݌�,�^Q��t%\>O�c��l��/G>�2���$����u��'
��S��W/���O* (�)��PT�\3؁L�d%�0e
ꗀ\b�|Q\SwCh�]���s��V~�ݏ��i��8����Bz�=�k��3���|xW[�K�x���+�8k�xW����'u��]��Z�՛#>��N�{�\�N��Y�v����9�ͫ-���7����o�q
�r
,/��Ҏ`$R�Ȧ�K+>(_e���d�"Bm{H^�k� �4_���J���O��e_�<�F�Hq�ShG�`�R��(B�*���.��6�ދ�1h��G���л]��ͻ��$� ����/3ԫ~o�9����Wj��Dޤ+!44O��Dez��>(�j�)-`�u	c�m�b	��4�ގ�X4�>�6��T�N�f+��I�������Y��$�%�{�ΐe�I�5(PP���ġH��EP\���0��+��zW��H2��#?����:�	��=�i(#v�*�c�qX�����y�#��=��hA��������Ni�Bh d��n��Ʈ�zP�
�(���w"Z�s�$sO2o��z�ݺ��X��v��f��D��l}�?'���� �����0�ߔ&4J��'���(}��@���&�|��R�����擽0��HԂv����H�7�B,�KБ�S��q���N�P��E,���a�]����[?�X�^v�Q�|�#���K�C�h���f��iX������Ѡ}��{4zX�ݩ�)ʠz��,_�޾��7i�}�k�W��-�T�w����`hm/
bH$��IkI����VLIcW�8>1ł`CT�q�h� �X&�YFc[��산
)؝C�E�q
ؐ�/2���]�����FP�t+�K��q"Jُ�n���ց9R�/�x���DVm�ڧ�Fc��//z�$XiE�>�z�"�α�'X$0_e��X�iOQ�o��Bk��0�"��?�[٤�*d�������'[�掹�c䩌t���W�m��kaf� 
{l济�7��#G���� �[&S��8��Z+z	� j�G0�5l�w������tS\�l�!�>o��$�9Ŀ�W@[�����82��~�~�GK[uz!�]� ��^[��ՐN�V'���]�}<�#���+����{:��kW�ǩT�62�K��{#ӑ���{'�h+̟p��Z��J�\	E�������)�<{}H+�1n�����Vٻ�9�:�KY]C]8J����7�4ÿk��-2��t��U�uO�U���EA�����κ�0�.h�e*
'�ya�L!�Ui�A/ٷ�'�p/��o�HFiN��kf)����n�V�a� 8����e��Tc�;���El�t����h�')�C�����7�`������x���&=3N�6��{���t3�2�I��:{�P��-x[�3�dNR/n��	�RK�%L�̅nO;6W�������N�x��Cj��1x��[�،i�=t�:��HG�6�d�ur�޳LVջQ�0erw� 䈗$P֒�{-t�`#[��EE`r9"��fWx�D)�F�n�"}�j�#&���s��9u���f���*^�������{���J�����c�g����{O�����%ʂ�qk"o���F���(�������w���:*ηح;3G�@_K�(zǃM�;0}�У���þ#kk�g�@��u��
�ݰbkY`�be6��\�)� PT���W~��Ʀ*�=�M�i�Њ�_�:�R����$��4����/���i��]�j2���9�	{A�h<72h�:G�k\�*(z�p��[����7�B�69t ՜�4("j�����k�ts��\�ED#��'B|:d�l(�ä27Y��>q���\��c_��6$�J��>���Wig���:>�sG0��޵^G�q�ΰQY綽'&���c���O�~yB@� q��IP��D��|��|C����7��� �����w�`"��M
;�M�V	>�+�A��Z0G�� �Ĕi��ī[!��*?��F�u�F�3ȃ��4a��l�w4�_V麑�py�*��F�����:�(�϶��:����pox�2��
�_,��Yą��E�����"���$��{{*��d�s��Zv�F�y;۵�����f�]�+)ՙ:���6��+�AQ�l�[I�^5�1�+����тd��٥+�Cb��0�g#��Y��� �-0h�	����T|"�AB�6J��ܬ�UA)
u�kg�:������%��_�sIڌ����~�u�{����̙� ����x~	�|�����Ʋ���ʬ�~q*�_����/��M@�2�몋�K�6��п�:�ye���o��\�l<��N�v����"�n��?�	�R�	�T�K�a���ſ��mse�]�H������wN`)Q�^ц4� ��/au�?h#�W� e����?-&�S���z�m��끎�~�:o=��O���M�k`�UX�V��R����
O��)������������dȲZbV�y����4$��o&^9��4�m�.�&��W���%g��E�pA������y]�����/j'����o��cG豘g�Q2R_�"}����U�c�@�-~[g��$g�q���Ӿ/lj*�����>r@x�2�D���rt_b�4�eZe��H���sT:�S[��i���ŪDKN�j�\-�2t���|���D9��1�0FH��?S;~ )UFUF�p2�D
���xo����׫����ǎwJ"gyM��Fڱ_k;zK#��ZL�>�XJ8�~�o���'��f�/�#Ó����ك5ݒ��#�VGこկ��l?�_�Q��������q����	RP�x�J#���8��Y�ԕn���BF�<#	N�Ʊ�o��ZR�s��<�a���~�M(5 #����*�t`u$��B��pԘ��F�a���~�*��>��w.,'1$߯�Y�̱ʴu��2�Lc��y9���!�\撏R�|�[;���� �{���G�ʫY���v�b=��#>.p�_:4/Tڔ���J�k��ˇ���FY�r C�Z���q��3�k]����&V��a���m�>�4�ߣ�!R�wS1�����R�L�{��s�H�y����H�E��lNU�PQ�Q����KgT=h5��&�5�A ��q.�<ˀN�صc�i��]��}&����&���N�Q�Z��<�}�s�����%lۏ������ޡ���WA�+���pyw���Hp0�Ҡ+q��"�f��L3wٜ(^4�'���u1�U�J MM�%�}�u{S�BhjE�?t�lm>��r���Uΰjꌿ����`��G;JP�s��t/��������f'9J�B\�n]	� )�lM�Y7Vk�.�U��5���$�P hC<f��g�5����(k�+�1c�%k� N��\DiG���:謗s:�^�rJ��E������
���|GU�&Л.����"�ቺ�p<���J.�IO<nzEb�K(��F���^�z\�H� �xp�$ԛ0t��i�l�H�$
5�D�d�^$r�h���b�e0Q6��#8g�7�L󅨔��ĕ;e2t�d�<����v�su�u�bG>��ZAT���^'�⢮���Ф���4SX50���b���a����ʢ�u8")�c���m��F���J�? P�l���?0'pO>�e���w�r< �E����&������t�>/�S�,o0��Qm�Pې>;[�ݙ��W�`B�17�T���g]��g��Pr��������{ ����c��X�G����*>�R}�MG�:%��$��R	 h�F�q�W@�Y�I�U����u���^�lȡ�#j�j�#:Ś���љ���I%������m�����r����	�v�ȼ*ٟ�!R��[�%�ӷ�d��y�g�>��������A�W�E���P���ba�)��\���4��.Bav���4������Q�'��`m#�	���!�oE�����z�'�9���yj%|~#���
�Ԙ#�mԴ� ��7/�eV�_���D��:��*�T�IC��W�����d�hpD�|�ܾ�1�Iy�����i��{���äa���CjlX�B�;!�Z���ʃ����G�Ab.�d��O�+ �b]%l,m撙�2ȣ�N7����gi��o�$�Y��GC�9QcȖ�Q\�xa�<��3���vj*�^_HA_���������(�G�i�hgU�O��-����e;��Ur�yҌD���B�sJ����3��욎I%j�z��$��v�dL�A�=K���o�:{�2"H�I.�s�m*ϛ0=ކ.[�S��uutDޱ�{��n��wsN��RBQl�iZ�j����:�*�����V��đ�6���VXuJb�����2�+8�t\3c�	����Ce&b�'E��ڄ�!#i
0�X>�ڲ��"1w	R0X��x	�҄�]+7>
s�����`���_�Y��)�g~���7=����U8F�}ԵF|������\gp yDT�����4!��.|���r)W[I�s�e���@�pG @ w�d��Y���X}�\x1z-b5֗�BvЎ� A�΢%%+�����;��k��c�I�m(U-��Ў�j���0#�گ4%������;:x�T�u�x������p�n�_����F`�c4�N���#B'f����1Ҋ�5����Д>��v���]���YA�
�U�������J�d�yb���a�V����>���6���ұ!VE�w�n/�q�ߕSiRF��.���Ŀ�7>Ʈ��E|b����K��_�7��t*FK�����Ҭ��R�]��'z4�I���-=�d�">ܣ�5�n�L{������(���6��J�,�2�{��pf��R,$��.J7��v�Ҳ�k	E=��+ �6����Bл29"� P���q�����G�W�F�4*� E��?�y����!tV}cq����j#,<p�D��Ai�[H\W���B2��®�Yp6iwQ$-F^�y*.�)�׷%Jh�� W5��P�rMD������u0bV���L����Se�9(.q���q���`�_���P�(��^�o����ʍ�&��F5��z(6Wt,�����@������W$�p����c	�e������Ûҿ��Z�
7��/�B���l5�1��Z9"{�?��:�s{��Ji��x,�8��Ê!;\+��;��}^�� U����8'��u�����Y<���Y���o���"��cי��������s�X,,(��W]�����de����/Ӛ'�SY�8mt���Ռj-��B�Zؤ9jl�fy�m�3��;�W�Fu���G���L��N�,
�QwX���|�;�E-F��C����I������`^��q�Az�������Rw~5i�*���r�x^x�f��׍H\��٨6��z��NP(��ކ��߰k�e%x�cO����[�zJfUЫ�z'?�v+U��9^I"��jۮ��'����İw@�>��U�Ƀ�?�z���p��O�2	0��a&��f�"X[�a�����#������1p>m`���p�<����-��.���J�o�pҽ�}��ON�U��z'��""~`wno\(��D��#;�μ�<��N�R���+�'�tNl�p�����J:U3�4�Щk���Z�>�#�'rQN�c@0pͭ��<ŗ��6O6�d*O�]�ENVe+]��\��S���~�v;7���X��Z>�ȼ���a����H�T�q���#�ڹ��
:���]���M���5/	ib<�TmG���*tb�W�ִ�t��s�Sw1zL�c1 ��h����fI��g�)�jR��-�#d>��f��w���&��k���J3~d��6�>R|�m����ѣDPyv������8�$U��Vd7q�>
L>��ㅿ��[� �|+��&�_]r=�xjj�M��S���}|�)� 
A����)��̓�M>�o����w��������a���{8�ut{ '�U�"#�C�R�����ǫ�]^� ��xԦ�ي�^����0hM2�IR�Kz^&���a�='�YtIY��icY>h���/s��`q��H0ɑP*����y�%z6ܤ��ʢE�ŭ��]�B�%��n$neQ����*��q���˂�����c((z�H��!�B�T�
 �S����'������D	y���p�p��