��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞���Q���F"�O`e=݊�+��x��en�D5��<��S�� �P2�{H,jcA%"���Mq������ge�Z@׸�"�SKQ���ڷl�u��;E���%���E^�/�&���(�#,J,L^��ľa#�������E�w7��>)��p����#��u�\����i�=�,�2��X7�\e1u<����Y�6|�m�2L�����c9�rb1�Y�	��\X��n��87;E��/c�O؝�cnd©���V�Z��m���<�g�CG�Re��ga��l�;÷�L��=b�e�1@3��0�{��t�Ca���!�t2��g�M8�5�K�>l�5�vNF�V��ҁ�JI1�/��d2W�;^��nn�c#����p.�Xp�Ø_[�?.� �|֋� ����ww��#���jU�	�n++��6��E9?�)Sܱ%�]����^��R`��%�%$U~o�쟪X%�+3����4�$<D�ry�_O�d�I3Z��5���r�&Y��Uco0��i2m�bʗR�AȊidu6�%�2fU�l}���TMP����~)�"��f�D�@�u� =K��n����o��#�o��<\�h������TM��H|(W�P� �3z�ZY�X�p	Z$*�tC��>�����H����}�Ğ�	�g�I�e��le���d46�~�l������WD��R��KwM�.6��m�<��u�k��$�s���d�y�^
�D`� �#w���m��"�Xy�/rr�ϭ�)6Fzn��a`����h��XI��4����q�<vb�]��%K��h수����{�k��k�v6ܣto�p��E+=�_fMx0YO� ������
���ed���{+�$�"w�s�P^*�n��(��Fb
� �T�Fa6�1^�t9Ԧk���h��䌛;�ݠ���w%	��-՗�:P��Z]y!:��A������=�2@c�fKG `­��k��#�wkȂ�zP��U��N�m�PУ�Ϙ~�ܯoR���>h=��p����"�vE�J�
tI�$�N�.�`w�m���A�P�]�l�N��l|һP'��*�8��W%���[t����A~��벛V��d��K_���.촨���&���dSP�E�<�m��h�3v7˿�ݑ߉�:� g�$��Z�S��7��v�p�c@L�B)ȔM�*������r�#)�p�d>Ċ���A�[l��wwD=������sC^�hdU~�F�݉n�Òxl+��H_ARM���\����X��k=����̓��X�T�3��˱&9���g���������[�L����� ~c'm�
���^8,P��S����3�Ke��0&e#�0�`|�9�jb����F�=�\�h�TUf�U_M�L>��F#17
޿�mQ�����4=�p���y��A�{��.e�����T�#p��F.��I�P��Ķ��� Հ�bX��_ �*�?]�ya�uG���>��0��*b���/�@���� roM{�Pມ|8���("��j4ҿp7�I|���eu�w-��5����^C��W(���R?I�ԏ ������ݷŬ�z�W�T���Y�{�ň{�,���1��"���СCc��ړpvIY����I{��d���E�7���;��_/�f�:�T��6qU3R�!�O�MY���Yʱ#G}��<��Βz�|�pbu�P���m����x�ʷЦK�in-dܺ-���vH���]gU@�ROL�%�+�K�"āL��{��zw��tL��ԣ��-�-c�~2}��G�t�K���
ND�ܚ�M�&ty�6-K���;�g�j���m������geܼ���I+и��g,n˸���j�zk��M�J��vU��]�E�1�۬)��ҝ�$1�����G���g��Ajת�پ�����x8�S�!��Hj���&ӐB��W��i�ve�th.�S}�-����=��itp�	��Z�5W�ȑ�'��{�&]`�$Y�O3p_��RF��t�F���8X������$����N��d	�,8�^Y��a�Xqca;8,�F�y���.P���5�i0�Y���b<� �Y.v�I��N'���׮�R>�h�[��ޒA����X�<�Ou�
y^4�,m�����m����\�b��K�W���IDiau���J^��o���\]}�(����,������F����´�0�cN$��L�� ����k�޺J�R9�Is�4��{`E��a	?z�Hz��Un/�ω�B���9F��c�w��!f*�)����>EK>�};��g@�lڏ%�h���Z1�ѻ��֨[1[�������!�E~�٩��$3�S�_!a48p
P�JXa⦝!x����0��v�'n�\���%o���F*���_b����z#�&��lԒ#Y�ȯrq�g/��2N��|��pce�r|&Q�ËK��ǐ�S�igE��afIV�5��z��%r��;_����I���.���.&�5��&�fq��5y;H��GTĲW�:BeZtwPB��ڢ&�V1T�3��9�Ȃ�i^�,>��mM,t���v� �׿��d6MN�Z�:G����$���+0R-r?������璍�
��B1�qӏ`V�in�MU�;ؒZ�-&s�Lj�ߍ�4_���;p�x�'S���'����H�L���w~#j���O�ްV�!�\�'G��DK2�Et(��z�{S�JmA4����@����*�XS:��X����H[/�S����f�Q�o]�Zw�����G��5�m���J���?x�5"���tʞ�ڱ5��M�(N�Dܚ>� dN@M)����2�q[����������5k'���?���
�A7�a�t�K�υ�P��0��!N�%~��q�u[�$��ǂj#{�ZI�4�+��$�
k��z��ݻI�N�Bd����cF�]!�j���;�����XOk��2t�K�}<��\mRQ�0%�I�K�*���`+[��'�
�?<�[�ݬȉ���D�I�w�U7�QEל�߀z��&��e�l�'m� ���EY.��6ӗtԦX~Ta)��%��5_�3�vX)�FA����ب�t��F��"��dDa��9��� 9�x�fW�Zߛ׆X��o��s��a�����Y
E9-�Zf��fx�:<6y=� k6���MD�_V{�5G�;�f�E�[и�F���@���P����Y�K����+D3G���^�.l!тh�O툪p-V����=�+���]
K��!���󨈡ԌIv}�`A�@���Ow����~�����G���ҝ��ub�k��=DK:���΀Epd�	)�3�Ul^�*P��	]���kO��<�v/�_���$�$2�Su[T1�Y�d����B0�0���uඨiyJ��q�	��y?fv�d9
�]
☙���Y]�,p�5� $�ݩ��D@�����A,��f�/�0�f<epď��O����q�$'�jc,R�X
�T₃��A��o��N���5��Z����Xp�T��$�i�M��]$��v@[���zy�]�:4I�,�k�����c�4��T,���8&20�����E&�qV\�Xs� 
~^�K�,� #�F$�U�����L]͓�;C(�8����?)��n�Pq�2{��{7(qZ��-M��>�̩b�"�.�Hp7�N<�1�*CM-����Ta��2(�5�-���o]kx60��(��q�a�+�c�^?7��R��˧���zK�M�} 4�F�Ǉ���1C2�w��p篺a�r//�^\�h���򌸜��l�L���]"��sd=�w�qU�$�W�R��ށ���	��o�a� �<�.�&ebc�1���Ҟi�37:��l�6h ����x2��D�[c�/b\f��`���rP����`���Ǫ��!ls
����B�ȑ�И�	�2�%A;~��O��^�r�����:��֞�2]+zDx�0^(Xb��Ȑ[�n�^d���-K�u�,�¶V��	�:�&���A�o=i��~�6�U����zs��b�f�!ٺ{R)���تtę��s�c1��)�.��@B�;1�bw Y�t��</���"����XAqB9x&qJ\��ʡp;s�|��Ei[����K��\��>,�Kg(f�������%��߀hW���9ڍ!�R���2�JY�MC$r�K�I�_����9.��lc�+	��U����\���d��:S����Qr�w�Qm�����M!}�tGh�Z,u]>{N�c_:bDܽ��7nɯǩ����v�[ Lo�O�~���eo��2%)���f�?��;�_1R:�� q����k����p0Ge�(�Sld�tt�Q<3q��P����Mg�@�XH�wh�Le����wC�-�:ނYͻ��T׸0���_��#��k�(�L(�A���^*:���;_C���[;ʗ�����9��YL�'�8�G��:Jo�x�yW�{�p��8٦��v�(T��#�#��B�%ʖr\^�ͽi�T����5� �j�	�h$��<A qJt���3�Υ�KQ8ӵXV w=OB�Ƕ���uc�
/֒���O�TFIِ���:��Z5��{��]���^++�a�PӠ��uc�Pɞ�,_e~�7�b�cotm���<��`#5eo���=0�2E��:�t��o��"����I�c74�h�� 
���NYdO�$c�[}H~5�B4�hV/��<Yb
���P�l�W�T�s�M��Z��Ӥ���񱄬��L��'��d�#=�f�hJ�� ����f�h�i��*���YOz�]��hq�k��Y)<�-��K�*L�xsfUˌ?2ئ��Bx�����җ`�;�c�{�Hl�j4�ھ�ez�����9������~zx<;��%����Xe�;ܵ�D�te�Q�ޞ�`�z	.���&=�jK3m��3�A|үgV���][�����wK�U��F�sԡ�9��=�|�l�%��Yf�ayr4H0�[]\W7dT
]4�`T�N���oJ��fNn~��39)k�����	�k���4��Ѥ����?ᆐ��u�5=*DZ�	T�^E`�U��W�t��<��=�e�$O�<�<�a!^k��R��H�)���RWK*�^s�룓����}DRD�Hm��Ȇ�$Y\1��Y>h��Fߣ��J%�0�6���#��jT�I���S5!r�}LI�>�Kp��娑`��=f��0���z�N*�9��n���:�Ȧ�'T�F�:�P���"{�l$�Y77�B�1]�'��s:�M��*87w݋�k:}����FH�q�ؓ�Va&92�R��ϦK�hc�=�ǎ�ا����Ҙb4� �<1�.�\s2�%r���C�zG1b,wn)�8�Ɓ�զ6vӉ&�#�jC��������.~��|G�Eڳ�l<p�N�'�3�O��C�4PO�?�tw"w��j�q�`��5]�f�jro���Q�N
��B��R`���) �m�R6�a=�7�:&��̴g#�<��ԇ6��5��A`���4]�k��_�N�'wm���َ{p Z��2�+��
=O�z�Ny?��ٌO��z��,26���_��o���6��ɝ�N=�-4�o�	��X�%��EwP�C������Q��Hw�-�vhT�}=���5����h�h���r;5��\[w�d���U7�T�1Z�)�����B^��0�b|�K=%�u��9�'C������Z�viEIs����cb�뎀=�v����4t(:�ܾ��-;*�������C���q���$�D�`Z�v`�k)i�8�os.��s�Qi�
�
s�T������Vx�an��P����Ϻ!t�k��x<넯"�kGn̮It���@Ý��	ŋ��E����)T �e	�Jä,�Mi�Z�|�n�rT�k��X삥 )�K�O+�ئ|��uA�@D���! 7`a������;�U�&�+V��-�p��Z`�b�F�W��_IoE��*��׿�w�2���k�ʇ�l"q���.Y�x�Ŭ!)|x���=�{*�4˶�l�.��+��� F֧m/���s�G���W8h6���$B�ɨ>`]�;S���֌��_��k^k�ۻ$ѱ"?�u V?M�\�=�qC$X�'E
(nqL����\��^w!:!ܖ�+Y�)V��_d��O)k���i۶��ɗ��p����;��
��0;��I� &x�� HY3͕T��q�#�8��./\��Ǥfn�&���zB�
�H�	��Rb�)9�r9�͹�G�HtXe�=��}�q=��=_�Cd,�Qߌ�$�N��Wx�2�ÿ�c�<:�_;X[�
\p���=����#P��*���8)���e\х��ۼm>��}��LX�\=c�%?SI@"d@{w%��U�B���j��ٽ�O5X�#B?C���=�\�~V.'l�Ճ&��v��o���R���X�d���n�������Z�2�q�gGn!�z}����G��e��b��xc�U�h]/SD;k�gjk�݈*_� ���ɷA�ŜN�|��h�w��ePij�e���)c�pSp���k9�m���8�3�*r�H�@%!��;V��~ Q��9�_���D�h�$�E��4<����@�����Be�n��%ǣ��0��`��냽q�L�k�s047:=e��)�ح����I��;y���ѽt ���X�C��$����J$�74mt&��9�����U�>�/����pq
�FPޔ	��ʕa|�)ucS=�MX�,t�����90}�t�'�hw؛Z�8�f
Œ�6�i� ���S֦���m��"��	�7#��1H�~\h���-���c�Q�2i�[�w$[��݊gXN���p���Fb���7 �s��I'�xtf��{���P�ӝȡ�\��k�H~���i�U�Y$T�<VwT�l�,H.��Q����w�+����)m�O�ti5ĕ@�
4�!t���{�˼�s�a�O�#���I˾b�B�Eѥ�N
mz�ݢ�z��3V�pA�(�ȨV�x�HF
-o���|�6��;�a$�<����~7=%��E�:p�:����y�W����~r��A�V�=�������(&��Y?�=k��!l�>����*mA��?��բz�����xC�"{��j������<Ф� E3����)!�[������m[D���S���(�V�3&�O`�N>�>}L(�Y�^Uү뙯MI
�!՛�xF)>�~Ԅ��Xux����&8��8۞�Ѡ�m�w�7ڳ3�,�J���z,c��Sɠ���cX�S�D�7�>�~&�ڣ2���t�hf`
�pdh��W̃�3�����W`�!��[����j��.�� b���S���؞f�F�6�[q�g����?�6v��K���k�|�۪o�d2�����Y�B�Ò�B���<����\�:���� L��РM+�7˳,pR#��Y��>
A���Ǟ�o�u�c������p¿��uT�ف0�sap��"�yd? ����$XC�=����.I'`O���TU%��`k����#W~�E�L�YX�lߒ�&���K��/�2�6�c�|�Z�^�i����)�oDf���S����h���p�z;��`;�����P�������߅[<[�n�iD���I�����<j���^VF�Xe�,'�$�t9�|���\@�#+�D�+�4!��śUy���ʔ��}�
QBM�9=��k�����`M�����\���!ΤK�����ɩB�(x������; h� @�z0�FP�w�2�j���rCD;��W�wN��,��'/�Cd8~�Aɖ`�)4��#�H7W��fUT�砖R���8���;�"�%$�������'��%�!q�	i�1�D`�'�av~�P���i�,O�ø��zw��x��0:�ʹ��_�ZP�a�fNK�o�݄�+�i�ji�]�ŷ�"�$�(��X��~umѕl�PWVդ�b �0��S�o7 4����Cr\�{c�2-���8����H�e�����=��}}w.��
��~�o�Ae���m]V
�X>�S9hv~�����B�*����e���odGd�����'ڿb��һb��p��m����t��u�����C+��=i�s�s��w��eMPs���_.~s�Y�~M��_�g��z-Ǽ☬�&������D�ь�� ,f�jy��CH�L�V�?h�Χ���0���(ܝ)���8]я��!8ץRkT���a�-��Q��x|�@W�"����Cܶ�S,/��L�=n��r0
��V�{�:�ڄIgh"�h�G�e�D܋��V^���.P=����W��YӅ׉u^���~��c/ġ�{]��b* zkz~,����G4���4Eox�|=`ɳEn�8��G�1'":��KDc�::қ�T��G|��@��1r�����ȸ���r>�
/���t�/�~#��nh� ˺�,��6-	ch���[MD`P�5�%�	
�s�(�z>�u9����(n��TY��ָ�M���>�2C	>Ap�Z�4�֮Q�1y���O���F%.���<��џŗ�Y�8��$�{S�[��f��x0^Ԝ�y!n[G��+Y�Ұ����(0wW�s�FpQ�7
�� ��NRY|�[�i�ǖ��.�?%.���.)����n�Ӛ�*�O%�҆��V?�q�l��k�!�r9��Ғ)�A���$��!u�ڂ�'Y.�?h���W�D����%N��B�(��}a��=�Ο�pڈ�����d�q��@�����g�C������H(��o�Nq�h��%��h'�]q?�6�_�����W<,S{<��X�L�w��i�- ~�'|�;��,fB��ei��~j����>�AR�C�9���,�y���Lwi��0�jJ6�H�Fz7��v�uH��â�*��c�����5�R����QOB�,�1ggĪ3��D��d���g�x�R.5m�� ��H�"���j�(�I�%��6��ڑAe��)k��t����l��5�_gy�0ԩQ-�j�������mj�Ӂ���^1 k�K��fh�4<��6�̐q%�w��_��S��I>��u��AE�4|��7R�+�ـ"C�?�痥�T���r��618�� ���,�!��?���5�^��������;r^��&A���x��3j]*:���i����Q�-���F��O~�MC��������J�1���Y�{͌���N]v��Ē9x/�Pj���W�~m� ̘d�v���CpA`�j��y)�o>��<2d7O2<�_�����z�~l����:�fT������[bk�礭}d�D��6y�Ђt��ų-���VTT��5ߎ��?1�}��zD��m�^GӖP�����J���_5s>r!����ǐC�Uŏ�0�$T��������-��W��}r��l����Wj��C$���-#%p�xʎn�|�Ŝmm�	���m8^��A0��	,۪� �r�+ٴh�i��M��z<�Y�ŕ�}��/��&T�b@��3�.�4�a�t��`�a��`D^+\Uk�6��8m����c��d�K"�V$����OÍ�J��CQ�0jߘ��u� ��io�tϦ����x!��Z�[QG^4��X��|e�J���t�T�^�~�^���g����o��wإ�����ʙȷO�q�N�2�	�C=噆&�(��Upy�xvg��'3�:��/�.��r�ߔR?5 ���|r��ȡ>��7E��QU=�|�1�C3�%>FZ�?�]y��*lɑ��P�|/N����x�J�"���L�c4��o�в���"�@�ve:�V��B ��� � J_�]�B�l|�	�>��xXW`�ieO�H�H�k>>���x�<����_X�;���ϊZ��d��4c�6w����0mb�h��+4��YdF���ôN��p�k5a$;��j��σ��������1�16�y8�'3�-4_?d{���wLI�!�[u�� l�c���?A�GG�d����FX��P�ը���v�p������F��5r���<�@.��m3+�aYxS04�"�2�X�
����Z*��?�ְ��C����A���[4ͳ$�|������*����˂r�P>5[L�I�إ�{Xi�6(d�!'�����J2�F�$�J���zvX��8�)�2��0��f�I�udk��h���n��.uA�j��ν�=E�И�dK�L-�_��������tB�˥������Kݽ}`���Ƌ�(�����U���Azb2����GG�b���s�$�[� ����Ƌ�D��?��Z����@5��0�B�Q.�>l#s��&�)�5�<� ~�I0�s�ΐEp^Ɲq��*��(�D&:����\�8rX���6���߉^���Y�=]��L���n������*�G����o��٤'6S��f/��@��M�Y�$Xo�UᘆR�����I�Vx��H����K��e�ς�����9	��c��Yp.�zk����W���W�n1���G�%��f'�Ƀ,��g�Mv��~�4;,�4c}Q+�	_�p�����(`m9�
u`<e �(�����'���@������A���PĄ/X�Iy��8�-"]{���S(�`���3�e��c�u�_�>�>BU/�kBt!����i�4k!P��Fe�F����S?��;�(�V6A7n�ۇ�LA���n\�IPFٹ/(�_����:���-�E���H�_���Ɉb���M���K���	�p��;N�U�͋��0�~P,q��Q~��h�C@��c�;l"�V>ʿ���d��Se�\����6Rڲ�
v�%F� ���=���C~�)J�O�t��rp�֮�ͭ?�<�D�d��C�:6�v��+��V�~"�LqC�bX�� F�,�}&C)ÂJ�ǘ�k�hu�GI%�Z,�E_/(�Ok�a�P����kSn�y]�Uv(�ȡL�)՘��ņ,0\9\�J�2�yw_�^p����u����U���Ͷ�4��,O-���j���}�2_+&e�in��Z�������=���=S	�6M3p�zJ,C���p] �Y��o�}�]�@�l�K��_~_Sw��K�ǋ�o�qL��&�UB��#{=0�E=|!��I�yc���&���`Krc����Kqd��Z�K|#�-4�9�0aQ��J�`ze���Z�L�y��c��A��u���S3ELr��ifR2>jxh{��΃a�������sv������n�KOi��	;���_����l�ܐb��3D��s�?�<~�F�l_<Y���Z�P7�<i������zϴ)��&��a~h[��P�6�%8H����07U{͋M�x�W��?e�,]t�8�t>Լ.�%��T��$	a;��nf�u��:�[�+�ZB�fP
��*%�o�d�\G3	>q��Н�s���)�3�)��X#��){I�t�ދ��V!�P�@ë�>��l���� @E�rXa�x�m?�'���[�
Jât�HC@Z♑ϟ��ΉUS�or7}Ŀ��}�dA�����Bz#�|-dJiB5��Jz�+ʆ�OtT�̸ۛ��.�Ե��p�Kj���Z
��5t�9HO`�l�̠]j5�g�L�LJD_'��>��L�0�)T�Ż>Km)��&\�b%�k�{'M	�*Q&��SЅ�Y��n��<(|��茕-�t ��F�������;�۝���@r��>/Ù�[ �X����0���+����n�.s�:��Nz?���@.>wB6�z�_6ᯏ�����?�C6�|}����~�^�=v��ݘ��!(G�E��w��xNvJ��9tGTH��D��E�UUpQ�����Җ& �ZQ�a \±���)?׼: )�l��&@F�l�P�H����������B�VȢ�)�DsmN �-�#r*b�ǈ�iB�7a�x�ɋ���tF
e{�+��E���#3��Y�jhB;�-\G��*lj�(������DtDZn��=�`

��9�%��?�EYg���S��$s"���ƞ���H�r�Org����UK�H��v�{��p�m!������g���0�Qh_Y�*Dɳ;�Ij�9NI�քK�����Wͣn�k:�D+��;�o��~q��"��5��z����ִ�'(ƻ�O��Jz�tܱ�����}3������5��@(�� >��*J��v(+�����ts�5��Œ߼��a���x��*��5���?��uӆ
��FYz��K��()R�{�k Q�x����b돩j�#~�M;�g���e��>s�=�Np�J�u�l�ᐪA
�q:�A�����λE3��/��ǫ�t5�<5(N��kA'��y������������+3Lq����!zNw�W��%܄~9��+�Cm�2I��>��
Z�I8�1�Im#3e�L�Sex�N�#�����$c��v⼛���9�e�k�06W��������h\�'��Z1�1�<t���*��68	n��rY�v��K���QoG3qv����=�^������؟��b��|���xn!L�	��e��&�X�H�l��VuV��m3#�k���~��2/��ڣy�$N�Σ���M^�x�/
�t�;��v<� ��G�<�tU���� �i*b�^�������a%���\Kz}z(��駰��s�i��$hA����W��S��a��9	����!��˝��Ve9 hm����VI�XƛE�����jJ!4�W�?�T�u�K[�c<2��ѱ-]k�Q!�%T�7��^�dAX��Q�5�|��2ㅸ����[w�31{E�j��;yՍ�<h�q����xI-�[��2���ޢ._�)�'s���h/����YR���<�O������\��e�F'������Bct��:����8��'����f$�yqNC.���ߋΚ���o�Ƽ�×��Õ�x����L�ڣ�ޜ��$�[f��5���Z��'�x܈_g�����L٘%T�|��}�Ů�+�/�M{k�-�I���Au)ѾF��� >?�K��^������Q�,Y�)sm?U��	,�T���S1}k�eH|0x�{��o�1�wE�B�lg'�0�>pL^y� $d�fX�zkpn�^�)�h�عUrt��Vh(�`蟟!�~���Y��"�=!$��g�n_�#A��:^p�����aU��
va�-T+���~$dbԗ��9�ڧ�ݞ/������0�B`b��aKC��1��<�#�\�m6�9A�ڗ�\�۹�v-#u>��� 8[_?�b`Q�
$��r ����g��|��7�n���� �B(p�� "Ĺ�>�9���qI˕+��vR�`�kG��)9�X�^�dȘ�;��ʄ�yKܑ���l	y��(�F�KG�GU�G&K�U�(�g�<��VE;A0�V�$��h羀_�l5���*P(�.q����%��S�	����d���Lt\N�D1.��}���F�����/1���\��%v�ܷ�>�����R�媑ܩml��/��E�I��[��!��u�����dCpS�r���^�,��n��EV�%��e�c��<���B�4~A��MĽ��8Zx���>��~���q6�  N�@�T�G�������-3�����3�y/3a� ��MS��h$^!&����W�Y=�X~��Z%A�?�~�xI�����������)�l�$�ݺ�OiJ��g ٍ!\���E������7�9��@���\x���Ζ#�4��2�i	��<��6̥�;�:0�C*�	'��;�i<M&���n����<��.���"��V�j�羘U�`��D��I�E��㢂��hQF��)})�����=��f��xc�a9B�˜k��5��(B.���p��U�!�f2��ıi��xp�n=�� ���uE�{�*	�$��Vs��}��=P%���3����V��W�w��Wۃ�,�e�O��v�z�l[֕Pxp�:���^]��,>b�s-q/����L=�O�#X�q���s���Z��qţ�`��$^�.y�q4ߵ�8'�"�՝��\z���

�� �ܔe��Ƨ�����ӽ6j��ߌ�tDҫ�������TB�Z}#�^c
r��٦�+���'W��DB����R�������ڮ�v�b�����L��.,���V��ղ��N���v1fX�Ax�,�􃗘���?�P�=�SM)ݭ˭�A�D:|	���q�A���Y�Ow3^X��vH��=�1|)s������v�׾W�[��#d`jx�s����AV�lY٩�휮U'��_XNߊ/Y�7��GT}���V?����>Fq��{����XO�U����+7c�UjNOg@�Ny�me%';�d��9�.���M�!�#���b#������	�X7�U�/����m�s�s�0����c����=�����9�R$YI�W��E��a�&-j��m�Z@�xYZ�b{6{���,��c����(Y��XK�Pٌ/)�.&P���4�ϵ�z݊��]���F�����1z����+ 4j2I^P��{�HW���6��OI>d��	�̘p$ ت�S��{�璝�S/�?�\��f��C#����Zz�oۻ����D6H`?Lt-��'G��Y	�v�O\������vq��L��z!��\/��3�k��� �/�MYhSD��԰ED)�[��QQ1��hc����Ƥ�*��8Q��+ii��n��a�_�t�;:5�D�\p.[�� ��WcU�5Ba�+d2�mA�x��R7��kз�wWŬ��s�}{F���85 ~�B�0��� �~��)��øK+6U�j�!�t�#����7.���/B�~_��Z:����	���g�Ch���9�4	��7���ϛ
j�!Vq�a���.���!@���_�ʙ���1A:�f��꺆SdW�E��
<��pq~�m7K�R�P�O�f�|(��F�(B[~=���
p�PtX�|w:C� n!��t.8����TH�/6n��C��?29�ga��o��`��\����*(��J�+1u��Xxot�qɜ	�#3ȲPW	v��"�|n.����lң���,Xӌp�S;*O�١����Ѩ-`"��F~e�Y+��1��HnzF�^��\P�+�;�
%���C^��>x����� h��
���.�z9��y�oF����iv����C���[S��O�Z����l܇$%1�r,��dl��S�t.�G���S�u�C1�r!�{�I�(epE��8z[�X���������Tc�ț� s��m����@�l`�^?4n��Us���u����U�~��/'�����8&���b�"�a󤷼�lǓ�����R����y��z��~�Y��eD�o��}F���5n
J�⦵��l�4_�� �A��tJN�6��ĳ�Z��ɨ
Nop[gtuh�F�0�V�܍��3����nW���@��4kM�!x-���%��ݥ<�E?PjV���3���^c8*���gy�ychd4��=k	�H��>�����7V"�g*��ۨQ��5ΡĀ����X�p��eO�b-}(�5ح.=35=���IK��b��*�foZv�^�c��%>\P�la��;��x�D�7�:(-`?���[;��v�f�ĕK�H�?�He\����@l��,�ª�KF�nͫ���N"�nSѝTq���) *1�'��1QnFL|�Yt!��>:��)i����!,V�g0)+������xR~��r�lA����ݘ	j�PЮ1\�Y&��J�wJ�u�=�[(��Ԝ�gspٗ\XO����>އ���gs��o�v���N���_�m� ���W�<do�Ve� Ƕ�>H�%ׅ#)i�>�,O����v�;hx�gM�D��ms�|z��`�~r�yk~�W�d���y
�qs՗kI�,�7H��8Xq�:V(ǝ�ZRӦ<yc�^�˯��vԡt[���I$�j��R��f�{�W�U� ��Η�y�">��j���ur8���C
\9����*ȡ���ӣ�I�߯Y���Xϖ�$��N0^p�k���|�-.B�r�R��m�)CW3��u������u���F�F�Q�u�Yϣ��x�Y��+������2A6�?YU�*�<׹�(�:��/��.�R�ID��'�x��w7�	��0��رA��5�S��9"�w�%�����Ҥ��z^M�h�Te�E��`�[s����E��)�#V�����|�1��LQk�0�i��J��Rt��i�@�26�}UO��(F�M:��G�7'�a��� T�g�b���5�x�
S\L�s�m][�be�ar]��)�
�H�@��G�=��}	o&4��QUނ����v��F�C���y�C�=6�;�˟��^����=�c��;&w�i����b��Zl��*�^�WkSF��t�X�m�3]���o_����'p���>=�O��ݢT�4�Upll&�(��h&�Z�>��J>����mx��Z���CaU�O5�Ԍ�1)��Мt�ܟײ9��F1�V����O�8<���#�~�� ���\Y���x2��	�4�����V��a��28Hm�Sr��ѕ#房bY�)⼮����ՈJKp�>����ieC��X�ģhl�X�s��(�j�Z�����+��� 2���;���Ta�5v�|�q�������P4T�F�ud?����b�[T3�6r�����f����޴�8�FO���14=%��w#�7K=�$��bc`1IQ��l��sC=I^��U�\�t9F�9<� �{�iqG9F�c�����i�Dȅ�s�8.�N=��U��Mģ���A��rAǰl��Hy�%�+���Vz}M̆�J^�T���f6z&C)��&�({�<�o���ȯ	�sߨ8��~����B���ջ҅0� :6�6��!�p�1�4�����}��O�B���Fa�H���V8j-��]l�B�v��Z��Ơ)�Ezgr#r�/����l�N��)���_V6���v��dhu�xw��Ƽ9d?�|�E�T����"���h� �ܳ�7Vz�|�1�tT�9�;g���|�]��%r�4��g�F��WA&*(���@y��s犃)y����|MS�T�+���'6���k�WLn�
C�i�e����rP��̚���4�/&���j��h�Cuh�ºT�%�0+P�_�@Q�E`v+�yb���NH��Bb���b��%�Z熊\0s%Ŭ	Mw�>�G�ۗ�)�B!��lm2�R��t,tf茖*d�.�')��_8]�J���.).��Deƽ�&+h_L��f$A�J5�3�=�b�}�9�">�:}?٬��EL�.����6���>t,��e�[仈k���bZ��:	����e����\Uר��-le!�m?'p����Y��WΝ�`vQJ��ϰ��Z�"IP�~�����PRD١u>$uUx�ed��L��5��Di|�513�8� v
�9��Z)a�D�$7�g(q��P��)50���
#
�N�Hb@�h�E���Ь�ʿzM
.iSG���a�W�I!�u=r޹ �!ޡ�jw�u�gSv�Vw��뱫�L3�5��}/3i����X>�f#���k��6�	�덕�qӑ@��ٱ��-.][@���N��
NGJ]u/Iz�	��EUyKQGS�"!�e��*�eu"�H�a�S� @�O�n���Y�4*�S��v����1�|Ga�x�(T�������@yW\�m��M�P���p;qFrظ��Z;v"���`Х~:Lփ?���[�������G�U���� �Si!�ŧE��n��+�Pђ1r�x�Y�H��lj��Z��:u#^�c�YRt���O��ϫ�O�u
������i�xcB��slN���&)鮆��h�x���=�
Л�XZ�2��=�3޸�H��w����0��Q�k�R�"ox�R����/�,Ks��8�;��Ñ��W+ȥJ��&�</�_�Kd-��p�%���q���g�����͉^~3���X�M�4e1�s\���=t�cO��LJR�?-3Zd��!ͦS��[d'5��8Y��?������C&�N��De�;7�Վ�W<�h}2���x���T	�.3E����˚B������Cy���P�pk:}��}�
���Ӽ��M}gka�ڬ�Xِ���1��R�Z���T��iD��qe|_2��b&�$������N��.�0�ј��ة��-�	[�p��.�X!�GnFi�mN�Q���Ą���t(Ckn����`H?)�{X�����rF�i��԰�[�$�Tj����U�g9EJ���b��%T���z9�(��{��/�CWZ�"Ŋۻ\��Pް���e@�m���{���W���=|�K���Wί�5��B!�h�-��ށ1�8;@�nۅt�)�zcŦ��҈nN[�ݥ�"���G�%�K����+$(D���OٖBA����ey�Z���M��9�Z�����|�Q�j�L��-��PH��ϥ�_H��.�GM�:O8�$f������^aDN�W}j�0��xy�SB��S��ص���(�3+�b���D�@�IƐ�3�|B9Ujt�0�7np_n��캔D�AM��.n�*v��,�mR�	���
��`�1]F �h�ѫ��q��3��"�-����Ьd
Sz�����5��"8R�����f�1��`�(L�;)��T��I�K�h������s.��p��Q��Q��D*���KP?�v�������
�ā(䌞��m��{	˶�� �����/��m��4���1�	Q�4���$��]�$��mC���Nݥ�J�2�bT��#&�_�\`@�lKl��C�A:|%���2̝K���e|+4����.���X��e��b�I��:�콡��{�%`��:t�]D��ۗӪ��̥sD.�;����Tܖ(�x�.[@y�th�x�9��USbvfa�FIԆ�����F�8=v��p�p�ַ8?�)�+1M�H��%�k�(0�����J�7���V����l\��?+�.Y�ޮ_A�Dk��8N��,��r-B$�Hrb4�� `�+�1��֊8�&��,"���Ej ��B�Zr�-�ه�1-N��_�I���"T���҇��J�,��зb���}N�>��K� $%`��ԯ�N�Y�NХ}�k�lę�6�(�o/C�	)��U��܏�Z�I`�9�fOG<���� �Q����ƚP['#tNsMzz,=�H�V����vD���|Hn�	Qc=��ʋ.L t��$�d	��r����!�9�Lp�8#�,�i������D� _�c ��+�j��`�2B��Q;��%���a�� 7��&���Y��n�(�7z���ȝ6$�;�I�����UW(�H��ie�W�kQ?uZ�	����MHa!�ӔZ-����>ۢ�8�A՟;92~C�&Q;���������˗ay,TM��.|�f���E�3D�.��458�e�|�,����9��7�M7x�k)V�� ��.�n#�,�$-��	z̉v�1�w��)�PB^|(Ac����k�����(U��B's��_
*��&�O!�e\�\��G����p�5O�ϑ�eO�2`��^2muӃ��Xk���v@�{�$��5!W�~��>��L�"50/ō�~��;���{�( ׋���yZW�����̞�\8���^�#ʣ��@n��@��yV��f��N���7�FG=w�e���s�p�d+G�ݩ��4�;��h���M�����g�LX�!�_�q�{V�����d�\�i}�~)�h��9V㡄��$�R�n��N��-	��0�-���ؙ�j�O H��"�ܰs�� 2+}��2h��V�A�bq�r~5��	����2��!�l���d�1 ��jj d�!�txA9n�����U�&�f+��!}\�[���׾����+?_��dy�N��ͪK��'��o���v
�'xzcb����]`�!�D���x���[�����$.dH�=����KiE!g��.Z��{�*�@XMV'���S�/ZD�:K�9(w-N���b����#0>�d�v� c�;�;��
�\V)!B\�~���9kr̅f_�i7��]�1G!^��+5����֍�_�ZD$Hͺ��M��b��C���E˿�.��9x���,�?s��ҸL~y��@1�vA�=ϥ���/��?���� ��C16�]��}�0�hO�Ct�0�Ǟ1�=��86�y������.
9����"�ɻU��{[�ǩJ�+n<�(�C��m1��	�lnuag�o�5�[B=bA�B� ���]�Mt(���{�~��jg����G���#�H���q	v����lo����+��<����fن�YJ&�+�5O���G%�q�C�j.0�xe����tZf���PV�/,9�av����4��6wẹ=���XQsS�gu���I�+ }�27t[3��Hz��<2kvrbtvf��c����<4�1w{���2�+I+Z)�2/,TB�6�}��1��%q*�&��+���]�+@�jڵ�U�iub5�t�[��P딲��R�g��\�C��k�wH1� ք�%�~��J�y���01JOlEM4?���J��$)g�������ᗝ�����C�{r6�9�W7���a=��!�h�w��6�)�v7�/�ym�3�,�'�x:ϒW��V /�%e�=ntW�m��8��n�BT��$$z';��Q�P�3	d����٣I>?��b�?X��Y�f#6O�{_������Y��܌Q4}j��ݾe�� x���g����k�O�+L$�X�	!v{�����$M�w��4:\Q��i��3��lKA�5��6N��Ց���2�#���KB/��D{'�-i���X�7��^�͜{��8��¬� �Cuԫ�RL?��Ph�7IF>Qm�w{��;=Q�M�1ј�E�Xae�-��FD�lF9ÿ�S�	�m�a�L��D.K{�I���Ք��B<��BR!�������gT05d���g�%u��=�]C���ŭ݋���:c�/��6r)��[ZN��b�^{���E��_�ۀ�X-�RK\��@�0vˤY��\����:	p8@ |P�y�g�|�)�������v��
�8��k��D������(U���Q��2$
�NuB;�
+������Uٔ���E���'Y$%V9��	�P-g�+!;At�qC�L��OF5Æ��)V�	����,d���U�Z�n:��Z�M��_��Fσ�8S���T�����Y'��*���_���j�����ȅ�I��\�R�E%^����z_.3L�^x���<�l��ǖJ��#���O��d��-�$a@w/YQ��d��
_�_΃G�b0�>b%%ڐ��듛��ȣ�����Ã㘷�A��o0ă�s��IНq*���#��6K��$��ES
j�Ϗ������K��|�f?�%]��G�cՔz�ߪ6 �qlbX�`F���g��ۤ�x*/Cێ)�QP6wb�
!�g�Cc.8���&N�S �@V�������>
dۯ������b��&��^���¡K���s��r8h��ٶ�X��9;d�A�n��񀰿i*#a`	�2�?�u�����N�b?�6�u���yZ��k��d)aep�N(����V�(�s�״���R��^���5=�wB��{P9�$��C{�u�g�z�j�S��<k����=e0dU����pX���G�3PGw�6�Tj��-�nh�m��A�>���kSgT�B� �����g��f���y(��W���b�
�����|����l�Kb���9U�����)Ҏ<�/G���t-��;�SC�*>%����Yo�,� �{(���a7$L�ia�&؃xhan0�#���6b/\��p�F�7���$w��w���4�k>���m����ٕ���d�f�^��
���_�5�rV�N��N�r�H�c�fM�'Z�|s~�W/-]1��Y�$���W����y�D��p0�\�P`�ft�w#�nFHA߰���GM�ҌAw��T�
J<{Y:ڧ"x��>�M��|���զ��_f2}U=�W�&=�_����R���U�Y�@A�����Pli��'up��F�M $�hm�!����(柘 '�b����)]��B-�g���5�I��
����-$L�W���F��̠����/��[9�[I�	��AÊn]�Qi.j���P0�IgX0�:1��e�ĞX�v�����A
���A�8!O��&Ho�R��n.��M.�Ѻ�F�z�x����I��S� �F�g\p8�9��z�����w����L���O��M��z�_JVK攵�	�&��f���?7���v���שvXfe�E�����$�q��}`��G%	� �L��v �K�?KB�C@�9� �yԉ�L}!3#�Ѽ�A�5BD�?]���Q�2���i��~�QR�g�Z�MJ�q���ID�Hr�!��.��!c9�(E�=���X41����=T4�8FI!�@�9������A0���i���EoشS̄x��T�i�"5z����R�F��P�5`:�o"�7��� �M��.hp��P(	w�������Z'�T�Q4�U�Egp3>�X���Aê���
��WΖnmC9?��.��)3���K�	�V�=��F�x	`o�b#�l����N�K�$:�O������X��{�\ѓu�ޮ�3��P���Y0�����uG�I��W����g5�7��Z�r`��Mh` i�L��>'��G���ׯ�qG?��*��!�=���h��]���	َ?�sDaoS����jڑ]�=��G�d��R��Mb1)Bؒ~�B�	��X��fr�r<hzP��Zxg*e�{����t9�\�v�E��䜴��7N�ȥ��������y)-��2E%�[���#sk�C�>��׊lt��m�)����?��8L��ߴ󦦂�{qe8���}z�zH��fi@(�ࢵ��	_�E~�4
z����{� T����B�l�<�i����^�|�� �̳1u:�/^�Q�R=���+eoj��A�ɾ/W@�oI�c��cg�?�?��͸D�@>�\e䴗��R�mB��2��~�w��/�l`��2j��'���{���dUCl����|�X�z���Z��g�fO���g�1���nļdv%Fӂ2�>8�]a��N,`���u\�1�Z��j�5Ma�p��@�zZ.ļ� H��'�5p���F�tz#`�����i���eV�?`�q���� ����abfN!5�gN�-�"��b���v��δ�.�%�� �"�P���\/D�n�#>�7�P{��L�B5�rVt�Op�{�#�݇U�>Fn �;�d��9�Ema! �} ˔�*�f�^=$������.6/���- (d0쓀=J\������5k'�0y�Wq\�uH>S��^P� Dr�:v�f�����O0���g�%��&�3��`��E��v�e� ��l�T��*̻ܜ�u�a�B��B.���np��	�A_/���{r��b �ގ�56�]泱�?D4���]cN.����px��!��S�RC�m�tn�%��͐]��N�6���l.tw��@x��ǣ;�pεN�T�a�ͮ��F�����-8������-��\3x�bmm���C��,������r)x�ՙb�i��SFCXHy	[_���6���V���i��ۧ�+�9�E-��`_��5-��,~�����B)������zUx�>.|���2�� q7�RX�Jha`^nj��%@W�]�*˧6}K_D\)'䅸
���#�½�Rx�?�rMZh�M#�6����� �br�\ ?|���k�y�Ր��3�^A���ada���7Z+n�5�m�W�F�}��c��.=Kc@�-�i/��~'�X�~����T���<n����X�޷�@���3J�Q	�}���gѹ������a^��M�0�'��|�))ˬ��BB�����C'�����B����1�%�n~.z�s�Q��~J]�<|ߞ�'�ĈߪM.2�GK1d�2�)�����͸Q�}�n~T�A�����oO^�� �)�����bv��[�5�P� ��}���a��BU�$=P>|�����PkdOvJ�=���D�1�̞��I�(�z����?��Y<�Cw��!��M��X02N�y���tڅ��y�����M�B�t���ZH�p{����"kc�p�����)�[��n�!�di��K��X���u�u]-iT�u{���_U�����h�a�9��A�|0����8�)����{"o�U/�-V-�?׏�gߢCq����5���,/��[���?Hf�b�"l[�N�~��N2f"��*�Է���&�b]�!^\MzdԷ.T����a��.M|��P%�3_�<�D���9C��7av�e���������O_�l��c�c��iv�ҋ6�~����9�yt��;؆mB9�u>�j����i}��+�
=�#g�-�� M6�"��g�H)�fj����7�t0�Z���"������cLnE7���ai�8g�4�l����[~e�Q̳O�|�������χ)���{��
.ϲn�O�Zk��R�����r&���/��q5��{�ZW=ٗ_v�;�A��ҔM3ӂ?�dp�_l4�(<쫫�rn�h�~�m���(���&̏6�Ci=�_I\�K.w�OK�=$v#m4;,;����2�N��E�_�|�x�w�^��>��l���h)b�{kL?��>��k�u	�E�l���[���v��a�$���˽YB?�%g�QŬ{L�S�v���&�h��]U�$�2jD�Q���J4�Q��.?B����U�\T;�J���'ߧ�9��)���]�j+>�g��ͫ^7A�^�����K&��
����[�:a~�@클�K��,��s9{�B��A��3Q�H�)���n�{f��c�H�� Q7�ʙr���4�#����~k"�K�x�u�Ro�8����p`9��m)����y3���1Ŏٰ�7]�}��[�V���������U��?�V�N�&���D0�>s��|X���~4��a+6�Vj�s���+�'nmzC/j[N�ׇ$�#��4U���[�	s�Q��P�V�w�O����?~���L݁�$��;���1��
,�H�K4��J = pm�fn�*v�XKs�PFZ�:I�-4�7�I)�	� ��<oi�>�F�����_�y��U#� �jV�i�P����J\J���Q{�As�C��<�5��a`ݧ�c�	��Ils�m9��m,��g�@�T����b��eN�{V�18�U�}�4Q_5�7���:^�ئ*��$'�x�r��`flt]��ߤ�yPp��7�ɻ��c��8Y���ʿ��=���CN�R�5��&���df�)���I
��H���ms����>���7���q����b�^��f��m�=����w��A���J����	�-��a����RQ��<j�KP#�yc��n� ��f*�<1)�k�-�|kP�-B� ���:�Ch��%e�	�Y.�b�[C67gP��C���3>4�dIw��}�� �^r����58-ՋT��n�
"B�F#���Z��xIA-]�$��x�ї)v��[{���N=��B8�<�H|}$)�%��)�\e�z�t�˱<M�i��rY��k���x�7��y�ؚF����%o��2k���_�[2R6�b:\���ϐ�����o�� m$����ߦx�!"[�/�vCN�H��8V㗘��s!�-$��A��"U���
~��0�\��0h�ʌ�Չ�}k���,���{�_�y `W�N���}�ۇ>�}T*t&�ȸ�4]�u��}���� �N���+ʭ�^��^�j�8�g�t�^���8���\G��+b��WG����+���f�? ML��:�Z�e3��a)kgT��m�}�0
8J�m	��O �NdCm���u���':o��=��
���@zҷ@���)��*t��(�"T�����Z�A�Q��"T�M���NLTA���U�⤧f�\d
1�vӫ�j�9�I�AX?�srYL�;ZnQ1C��)4z�̖V�I���}:���>�'ͥ�",�����Œ�B�e#�ZҲ��K������S��迣M
'W|����4�����n]��{�f �6�}��Ct���R��`�H��[��!���(aq]#��\s�ϙ�p�9ᣩ��Z�;$�V�mҢ_P/�	p���hI����Ϝ*u�Gq��-�9��`�� ۜ�ߜLh�z��km�%��Y;.��M�t[k��.Φ좨"�γ~vw%s\F�ϯ�wg�j&��RRL���-*b0�n������|�2� T}��x�f<tZ#��n����w"'^���u����������Ӊi����ˇ_��F�&ZA�὞тVW��eϡ�@ư�[l	�X�zG�a�#�~���0�L�he���k����S�hI�֘�a+�V�_�Q;��U�8��ܴ��5�+�f��&iS�.F������f�S�S$ �k&�;Z��lO��ٍ%ɰ�ac�։�n�$�Y����QieP:;'��p����70�&a8��-W��\^�}Ҥ1&��	e���������%:3�Ӱ�]y̦�S�"<
χ@	�P%�'̔���,)Ɋ
��r�P�J�Vs��h1O��^�7[3�+��>�H�1[7�h�[`iٍ�eǿ=��3Ԓ�c�Ly�S��ts�8>ҳ�o1S� >��
s!�ϛ�>�Vv�Y,��@�����?��uM�� +�y�i���Z�� 5�5i�~���՘^˫6]&�uO~�l?5$��a��˾{y�&���pZy���W���5����K
�"�W��������LW�n���J�#��M.9隫���@՜�;��$RA�Z�Sw�d\qń^�����`l��>�kcKE�Ə�	1�w�t���BW�f�

d��4Fs�?���	Xj"��/�;g���i?�h-�B�>��ź�&��Z164�Hkq/`��b��ߖꛉ�'aCe��m�H��ԧ\�7��a2jq8Uą�`|3i�m\�ui��=^�����s`.OH����%�������t�!Tt�������G��	}���&["u}*`�xG����2?Ǽ�꣊��c�*)	��#sʥ=��t��]W��׮;q�?cn�~���H�H�B��+;���߽W��sM�����,��%�L��h�gl��嫞{�3`�M�ָ�}LN�zx�1�Hgj���so�|4QN����2���l9��������Ҭ�;��}�J&��Ů:����[���=�����ث�W�M�v-�W�.�5��'���<�C;ϓݶ���=F�	X��P��ā �(p��#��Љ_�e�rP�&����,�լ<�*ش`���J��լ�o:U���'�^k߄ìf�q��?!+�L�<pv(:>]0����)�%��E�r�?�iS"U�|eqP �)�o�U����s�TY�R����4�����>�$��7^�����)�_̙2���x�[0�wF���պ�U��	���Č����.I�S��,|��4��?ҋ9��t1
�cD�|�hd@���ZD���@��6�8�w ���Q�yE������?�}{�<�������cq�p���F�T���2�A���u]0 � ��r���{�8�|���/���츓*��0�hž6�K�#�c2�	�J�U�񫱿$E�j�B$��&���������@��g��lz3�9�Z��ۡ�� �8ݾ����}aZR�H[�(R_�͍��l���-z��ܟ�5O�J!+�RڊMȫ���y`q/?��1[ k��Rq<(�<8]�҆<������h��tt�z)3%K�$��t�#��\ђi񓗜���9��dz!���>��w��ơ/��Ǽ�#p�2n�LA䂐f$/8%JN�N�*�YF
&��vƀT�\��QE�[�f�*M�އ�`��C�
���ʘw}������ 8��%H?��}BEa���S��X�*N��S6=x�.p%�����9�Ƥz?��\��~zHx�<�M��'��K���r�߳ǁ�uJ��R���2�澋M�Kw����\`��4)��Д��jX�q0�j^�l��$���Z���׀�v2�jW��=� 0�gv/T� :�5)��"j9��qh��TV��#��{��'��a�+�-�Nb�ٷ?[]W�hGk����<�v��f|��������cp�]4Jv0�{�j�h����٫n��Y '�n8@*d�V�m��X�#��zky��4�\�̥Df&��ͭ���!�ˬ#��(���w�������.��ۈJ�e��7 `�	n0<�*�V�{d]�_���P���^{��;5��iD�tT�B��ꍠ\�$A�}j<�T��s�̿�J���P�쐬o�T{��4�$1�������u�A0�`+ݘ�q];Ei��]�J�U��]����gU�-��2y�j �3u�_n�!��q�7��$��@~�h;������rz`�F}��o�����|��O�N��㿓���!��4s��:��f.CʪI�/��շf-i_��˵�ll�/A��_�m�K�a���N]'�C1b�_&��o`t[�Y�Tbl��#\8���ז�o��=�H���_����6/A�t�q��1ȇ0�o����,G�P���h0�֋���������F�~�v���A,�
��}��tk�,[����y���OH8e'|����ۗ�"�P|a-�F�R�i�Ϟ�RI�Z@21���W�x�W�s]r�����Y��Ɓ{C�Ҋ}�7��HY���R�ĝv��*��
�Z��<�R0x�t�G-p`���Hg�ۢ����,����A��0�軕L%�hѧ��A�?:�&�4V{|�Z�xYU7�5������R�E14��v�ĸ�E���*t��@��鉗 @P])U��P?:F��?5��_>��$tz}!����D�y�M���@4$�t��֐^X��R)=�9�ZN|�ߤQ��i��Q�M��1dx�HX�.�#�9��׸=:K�8C����G�3�[�s���t��Ͱ���O��e>��u���p�����O��iP�g�Ѭ��Ȑ�/�v>��������R;�A��a��&~N���t������# ����<n��#��]?Hk�r)8���{ז��zn�b�]�o�J��N\�j��������i$��"���K.��<ɗw�[�P�P)�t^�.���h%���-�?��h�q�b�j���z��/&9���j�N�E�	Uf�H3Ġ5�e��&&�+�u�<�3OU9��׳8�L�( s�К��ͷgoZ�i�U���S78��)�_9��X�G�:̬p�OE�>��UP=�0��S'%.]��eh�p��g��܍z�YTt��ٍ9�n��'Ӆ��w<h� Tv�X'5�ٛۙG7����!�2�ό��巑�,�T�%S^�ґ���B$���{:L_�jٕ�h4��Ɏ/�3�-��6M�-=.&�w{���=ޓ�r�k�I*����_���|������ 5��̙��}:	&/�R/� �.+�*�g�`a5o%IL�jU䓎 �����?�^�U�8�/7Ӑ&<7�8�9��� �e������~�A*��o&Zr�Q_����QOKk}!�����7�d%a5���ɴ�Z��ތ��=W��!L�z�x��\�B�$����Z'u�}O�mŐ�!E��)B��VO@ӏ�f�؁����s���\����Y�e���+)�7��_,�cukϊ�oý�J���NT����ne	�R����:�y�A��)Һ���d���v$��l���M\f� ��{�fO���7�~,̋-����وdg79�z������	f'�b��s@��}mbh���F�}� M)i�eD�r}>|�5�P���&� s*"�[!��O���J�N[�� �V��.i���)��<����N�x`߼"�D'#A�E�YMJ�ZV������0�r(��l����#���6����x�{Cޢ[P�3��%��O��n��2�		��32Oc�A��?��'�6��@ɥ�C˧���"Q"���1@-�#WMY��?�{^����j'^uQZ��*r�ݲ�&��/��i��_[V;�{p>j>�џ�vTD1+���5�tsQ�����PM��6��:�����r���i�����z���r��iQ�'K�����d�˧��+��]ك#.q�b�c���I�ޟ�������s#��R|�"`��ܸ��z&`�C��`>������i��96�����ǈ~�̲�j?F����ĬUn�T-���TB�91�ʫv�sT��:��۰�:{�ٛz7���� �GD�qg�q[�SY艓<#I�uՙ
��rbW.�1E!M���rͲ^��Ol1K
BX��䆕.֏��ө /x��S5-m-yB�@�`���X��d��A��nb�����ϑ	 �XD�j��toM)����9-�pRy���;����/����'�Y)Df;�_��aw����<�\sʾO�aL��>��o��oKk�V�7h�K�I���q��!DL������'�]�/ףJC@Dv��IF��r�a�� ^����h��z>���y�0-���W�<�*p"�i��{��a����2��߸&�~x��_���2(|�ӼJ�w7�Ѿ�Rs9:�������g5��o�MQ�A0h���
k�|��B��`��d��.������|V$��/'2�6�륑B����%\ MFb��_�aۿۢ�aO���jQZ��P���%u�W?I��Aob��
wGa��F�$������YD��({�B����i�@;f^+���X��ʧZ���Q3����v<%�M�"ժd\�o,���+��*��;���w���ħ *U�4���$a�񅋭eG/�W�F�9�t)u����"�m��j�vq��KA�M��u���錴�#���jS�PC�A�Ὺ���B�:�T6��髏��ݎ����x	͑�O^�P^i�<�0���u��NRi�Od��f
��d6����u>ҭ���7mDw�:���Y�;�Ș�+J%���s�=��rg�~���9c��� ���d2:�4�D��)��{&�쌂�����Ϛ�.����vSu,T���׽�`#�����n<�7C��*�3̗��\�͹��t[�Ǡ0Z=S�5j\YG3���{��,uW$�U:�QaZ͑�Q��E�{TҬ���j�cс�cȀ��3��xyZ�s�m��Dܘв+.eF���?��`��*ڝ'$]��������_��	��r�U읳A���K�-n����(�蝟�SD3�_� y�~>�Ue�/��H�N
�y�Z�)&P-�"Dz���}�R�2B
��bj��X�E��� ��ό��ǂ�{�2�g�,���K�ˁ�ʅA�|hF �����
 PշU��v%̵�x)��y���Xٙ|Ee��E�	�H��`���׮g���^[�Me��r%[�V��x�EN�خI֢eEZ�K��4��c&�lߎ6��BE7���g��h�A��� is6�)�>}�wpe6Ι�����Cn�/�e�ZkkE	��X>��]��C nӬ6�T�r�g� 8��� Wu4�	/G-h%�['�$p�h�j��ƿ� �of���Kx�-,�w����K�X����6t�\��\�P7�a���8�㏮b=��K����x�C��P�Tnu�|�0�u���i��y�B:�����[��%U�N5������+�z�=�D?-�5��s<+ץG��ަ±K����k|��eW��*J��>�2A�-ʭ�h�^g홅��x/����tդd�A��_?q��E�&�q,Ӎ@�}#g���@Ɏ�:��gg�v� *�'_��?��D6;�3�<G��p9~'$�I
?��ҏ�)=��ߧ�g4���^����m5WH?g�gYm��������!l�봧5鲫?j�z���8L�F�B����ª^�ς�R�Li��J�׶	��f���{����B`{r�V'��O��@U
N+��`;�$�(!�c�|B(�m�-��P���;���m�Rn���R��D	1�%�Sy��۽��V��d���=r��}���^n���>��� fR��qz_�{����B�3��2�DNJ��Ʒ��bcY���S���薫dg^1E�[���8����q�e��,_�������~��[Q}6?�m����YfP8 �۲} �i�9/�DhF�u@+��}� �6J�HD�:�� _D�4d��P�7N���\�U�2j�����/�����.}+�G8���f`>"�ΐ6���/�?�
�L��Z����y�����|�Z�!X�V���eN����w��i"%��'OE�RR$NS�4p$�wi����	^7x�|���L~����+v�f�L�NǙ�5YJIdT�
��-g�:��w��[��A9�g�x��`&{%N�W����)��*2���@��L��W1=������4�g��=j�G��G�xA�!s�i�ٱ�8��l�7��-1�+R�ڜ�y[_��!&SF� `%���0{'�mo<� BPbw�j�-��a�~�T17�>#)#�������-��m�4��@���N���;� ��S�u��\�D�Ć��/������P#W.2S?~��a8���lK���PF���;u/F6qC��~��u�� �v=��&���f�_tGHj��tv���AG�K�� ��`�s���7g6�n���`į��`��ݤن$?B_Ѧo��z�Jc���z�<Ma����x��em�6� Z;�Y���ޗ���֓^�����h0ڻ\��9�c�i�N��J��P�L=O��|����|ȗ^�[��?������_��y�yyUE�r�zB
< Arr�x�1�+�rO�����i��T��T�R�u�S���u|��A)f�xv��b6	���j���^⸷�no�NO�g��4�v����V��ң���I*�)��2���eD¸%$=G�\���� t?,�X�HJ�n�nU��aF����7@}@��l�&��o��l4��K�K Uo.P��]��_�=��#:gd��Pch�l�3�m/ϡp2�ʨT6l����W� :�qێ��T�����=�L$c�ŝ��r�����ٓ��ݺiTk�)�������N��>{�GJBW ��Ĭ��2�g�֤����@��������*�ە���
B�����/��Q,�S���/�u:���r|+r���m���;���� :��+gwLK&��&e]�^�K���aj�`~����B�C��1$����\����th[��q>�����K9vW���U�qk2�qd�����
�>�_�>:�F#i��_���j�`������U����!2��{y�%�$�%E�dŠ��l��-���i~ڹOp&j5k \g������UF����Ji�9Fy�\ْ葲��ew�Y����Wbw�yV�~�T=���A�����3iV=v��2Fi�^f�i��H�&�1\�c���)��n��
�J�{���gM M�9��M ��Q��3<Z8R��BVt���*�����/��xTN��W���(j����+�I�q��S`�C1fi0(��� ��N�g�T&��yWź��U��՜Z�;�|>8rT����֝	�����ڔ+1z�s�Z�z�j0pߦ��s��k��-���ƞ�;,�y����d���8b�.$y��&�+Z*<:V���ޏG�/�[!��}$O��_�y���H�%ظb�CT��Ԋ^a���q�Ź	M	�>�ur��7��?b��uX%G��qw���_@�q��M�`Q8�]dn�\�
��V��f҈7u�]���:ա�\��!w�}�Q]�_ ����	u���v�\����%�>Ӯ�D*��y��X�_َ��IJ��<_+|PsNI����S��Yr	�=�l(�ī<��������cӯ\�RӦ�� P5��Rͦ#0�}o��)�&+DQ�NǌxZu�|,([��m��UlnF�������sٹ-N��C�U�ԙ	~]��
�WS|"~i���֟��cY}ƳLn��(��e�t&zW_|"�3��^Tyٛ?L$�A���/���_Q�l�M��-���RA:]���=�
�!�Ow�1�C5��hQ���,L��H�'3�Q�A��ɸZ�R�%%� �ܙ�=���
 �=���v��uF36��b�E��R��q�����1d)�Zm1a.����W�KR�h�p%�:���%�M�֏t
��-Cv���y"�D h���n�|�+��C0gJQ\��2��O����Z��.~_0�� +�瓐�p�J��5��q$��S ��d�J�ǅ�s�	DzY�:.����1K�ȽQ��>=d����p�,�� I?�d_G
z���pc�m]����J�l�g$�*)���������_f�a�2�����{���Nnы�~i���؝�8���
u�ݓf��-YV��0@{��.���{���cF�q�}x��s[��wy�H��2>Oߺj�{�Z[���>�c<6���6�JKL�)�js,��������ђ��1n.�!o(#-�K%9�8�w��� 8�ʗ�wy��~vpҔU�,���u���0���+N��І�R�Y�@�U� ƾ�">�	 �Q����V�cp"H�65��*���p�P��I��Ob=@1:}�.�����ʘ��!�B�9�U?xYm���ѩ��i?��D���8r��Rw�6Q�uiR�݁���~�	'vC���ȇ���o���O�p�Ut�"��d�����ICw�*Vˇy�Ȥ)�"eQ{�mR>y��� ���?D��b	n�"�v�
���:d��θ`��Rt|�$e��v|� B�ikY	
(�_�)�}]̦a�Gs���s(�h�Q�<��w"��I:rU�a��tyw�U?���t&ɁaŅ :�f��ɼQ��e�=��>}Qw=AbI-mpCF���'�����G�����5�}���..�?��9��2��M��.�Ԃ������!���|C�[�AŁPA������fl���>�#Q&�}��,�@/Nͦ��a����A,67f3�iiA �͋}Gp��k�r@z@�g*Ņl�E���������m?+�¬'���D�^��B{�B��z����ey4�\6iА��fT�Bl:+���0 K^�߫2�EU���V��ұ�b�tτn'i���*���&Bgk�Vi���2�z�2t��P�'ٰ�O�j�N<G�b��G$@�t�<k���R�����b<��߁���(�A V��k�y���5J�XN�#L>��3x��G1����0v��#�j��Fܕ���H�¿[���bC6%��ƂѼd1{�$wA(�`�g�֏3Pȱs.��l��{4{ֆr�|Q�Q� �R�jYI��d�ʈ��ڏ]��yv;X�s������O����>��x�rg��zZlaS�1YZ����"L&DB͝�厖��C����7pi��.���n�3t4�N���!�cYn`��ve]��O���F�tJ�'�@+�}��"�;�Q�E�����}꺦���nm� #�#.pv1w}�j@GJ=q��Hqv
k\84��D�5���4��`�	����j��byڻ��'R�GB���D%���-�`ck��E :(����H�;�o	͝J��6iW��V�c��"�$�L����yĞ߱뙝��5�oR_���iF�o�~��ḑ���g�^�
��d;O)5���4���}9(.J|��^s��(��r�jrhP���R &J�p���=U�t8b������-0���a������p�ɒ-p,h����:^�k��w����T"�$���W�CU[i@���Ʊ�d)��M.0��R�y�%��2�x�]^4�-��)��(��xV
��n���U���?aя��&P��_@�����Fʷ=E}�a�7���[���֒B��8�g$��]t!�俧t�1*�c(�=N�X�4���bMt�]Y����?� ׉R�E��;%��IQ�(h$,�R=����0�(��;��ƻ8�-x��� d�p�8s�Hƥ�)�f��ѷϷ�PR|�Z��[�t(�;��@����|u%��>piz9D߭�1Ǽ �sV�����khOO��7���@��4=�xs6 �?��w�����S1����������s�[b��^�$��l�;cJ��A/��x���K.j:S7hq����zI�c'��a����]ZO�gq��]�19�o�D|@~�n{��0��L�r�Ư Su�6��f�X���qU���/;hS����S��e��.O.}�x�;Z���2G��f�K��X�1��U$(�?���&�1t��5/��n^������H"|ٮ�L�hؐ��4i4����n:�#yQo��f7{
��?���x�)1�5LA���z�� pe_��fm��IU>�2��������kR�n�}��@�#�����A%�)>�?d�]>:��g��}M&gEG��	���(���o��G�]��@�¡.5r�����������zٜ�`�OYD�=���˷�Q/[����=�Y��
��^���l:�-ݧ���� ��TO�~T:@|$��/�iD�Fcg�y����K3	M�R�Y6h�@�*�熪<���l�i��D�s��X����H���M�*��Ԁ`�$��g�5:�`-9yZ('�pk�č��a^g�2=]BL}:32�/ ��P��.����k�]'��&���=����U�f[/������Jt����I�)�������,�X��K��o�n��ێ����QATOu����A)O�b8�c���1cW���yMv|�/�qs�)BiJ�f q�$M�q���|A�w\o:��O�Ak>ݸ�@9@���$J-�*���<��6��P����k.U)�cA��jh�=e�3� $���j�on�z�,گh	 ��}S��Cq��	*Eq�Ss��隖����<:{�L���4.5�%lt`fT��}��	�~>��2p�� Ѿ)�r6-inm���S���	�������h�1�'���{�;�o���h/ k�MWqM���4�fui?�����
֠��c�eD��X�o�7��Cn�'��}�J�@N��ӍR	�� ��h���Q�c�^�G��*%%V>Ɣ�h4����VG
l��#�:޵z����+�>+zY��E7Б�$�WskX�c�����I�A��ϵ�7�� >��S(pj��71���]6b�Q�K���$��UE�<U��\KŶj�aAk��W9����cq{����F{���X\@J�3B]!U!��͸�G@pLK�Oټ���O�Z��,�F4�Z�&|wA��.����;�f$�d8���~Y���V���C�a���u�
?��d�)�$�m�|[�[Ͱbo ����}Yd�U�w2;�[��I��]o���SI��A�����CP���K����&{�@)��d$/j���v�-��@Ӈg!�� �-��Cy���'|�k^�$��ؠ��dF�L|v����:T�ح}����T���B��Ϧ��[:������|�%\4����$p�˳i��^5j� _���%��}�g:�vc�5n���Թk�al�!Y���	`=nY�Z��ji�h.��t�r�4��fT�/]��p�-��Zd&��v��x��;���hWx�����~��w����t�e*!�T_����n�'����d�����za��$Wۅ�(`#p ��0�(�m��$c��_�p��V�U�4��]h����G��r�f�����#!����A-�C���*��l���6[=]���$��[!����7>�<�[�p+|4�*�X�+)&:���es|"��Mr4��B�B����ԒA��~��H���c��0E	�X�5-�'��~F�n��9�h��(�fg�6��=�2#�'e��]ܗ��EX/��I[/����y����_��o�E�E��;�l�ݚC��>�Q��9�%Қj��m��q��؉�Eo�E��gx��	
�u�P���r��%����SҐ�_�o�kp�FV��kȁ��cW�c/��뙰�����>j�)J���>�R,��q�-" V��Ar�+X��~���_��Zg�	Ob$A��MFWk�sWa�2T���[G�O
E�=�ְwu?�O��V�g�L�g$2���"���G:�t5�Ǩ���cԨO�2�s;ބ�����VKK��s��a!�$�#��_��^G,J�M�����7 K΂d�iF,Ԭt$�g}�X��d,�P��aɹ�_��#ޓ�G��% s�!_B�i�Ӹ�������1��uv���c2"FH��̣F�D�aoU3yq�0�u�[u�	�X�pm�!�5r�����j�ɕ���,g����,*��	À��{�����PB�g�E�e���^w��S�`�?�XTt���(�V����rn���R�T3`��S7'��'��n>���h���-�ix������*XF0���o%�ص�l���WGz�O�A��˱A(��D"6�oxiD<&�������
��1��-:���r~r+��A@B���k5;ݯ��/,�WVl�}u��dH_$s�/31�!�;�]��6"���	�y迕�z^��Z�������V��9�.���/�ϴ�چ�}��_�7&�,"l����V�o+~(pw��Z��t�S�;�W�����[����K�����˖X�&{�|�]U4���ڡ�e����G�5yI�Q�ca���rP�ĽM'��DK>�[q�B�ZtuXA�w��.3��>�Z�Y���iɮn�K�$�������6-�o��l��	�ַ�x���U$��;�a�0M<�W�@[���I�I��������R-a�cG����}5�Q�N��#�	��ț��2��ѮԒ���#�S]hJNf]e��?�[-D�4�����T�7!T��4xY�|z2�&���ۏaB�}�X��7m
~V��vc�4�J��h�p���سfy;6�5�'t{��l4���ϩ��.���gꉃ�� Ѻ.�]�
�Y;�����D�D.4��A�'"��h�/�.W�~��c�+T}��eFB�
h�
��2�W6����*t����3b`����e��C��iK��a��1v����?�RH�lZX^����I�~��V��$�ʢzS^c��g��Xd�e�9�T��z`k���J���H�Es�{f��J�����]��]�껨IC>�F.���m�FN��ԩyS!�a~%�N|^�R�Ul�;�1��gX_n�Or����+�G��Oglo%t"�9����gm�*p���C8��8���V���I�I��$�ς��S����Z��,��z�u�Kvh�Q��ʓ�V��"[&[y�`UX�_=�^��i.��6ӹ���w�	�<�N��ꐮ�T ��A-�q�	w�(�36{����%'u���l�[L�5p�\NI��2a���x����ì�>#�1H�F�!N���*l&���f���G�W��T�Pr2�a	bR�4\��V�����8�Ͱ������F��=��No�j�F@5q;S����4�ؚ���M+��@<7�j������(P�H:�/�1��T�x�5��'+}֔�@@N�v��m�k2`�L`�F�b
�d��1�ĸ�Ԍs�n-:{�w;�fsp tM8��}Y���~��� Ցo�(��I[Q��	�ɵ�p���)dk�a�O�����5��"	��W��C��aұxs��
��`k(���Us��7��l���.�ڙ�@:�)��ӄ�D�~bz�VG�5����܊o�2�s����-'#�Ԇy�(��I�Ϳ�Z1��A$�}��d'��B8�<>�����<���5E�v[&�\�E�2G\�rT�12�j��V�Yk�kÛm�nG��
��7�.��{7���J$U�Gcq�Fx���R!)��MD�3��%�J���F4�=�[0	��S,t�/�&hL~��R�d,�V��`[��	Ě����!볞װ˞aV�o���&�@$��?�b���EUp���D�4�Y�NX`[d���CPo١I�!_�
T��{�[�m-�ֲ�Q��9����HJFg�|��u���T�<h�7��8n�W=7ޭ�r�2 #=̶���畛G�ᱮT����{219D��ݙ*��H�
T��_&z[���{�=	�˶|���Pnל��i�=�ĳ��i���Q:�I�]��]*3�����'��V�%���&B�{�A���1�g�4%��o>�����) m<��s/z��ޥ���إ��K�����+�j���4tN��us`K_r�.X{T%�}�]ǟõ�_Ά�oOW�||�K�)��v��C�2��a��/��}I��
7�<V	���j�m]�rC����B���b�77�y]y0\�_�a=��Z��o����R1)�V�p��K��%�-.��e�PW:�CI��5�G�c�zU�u�H�.�y�˴�|:��C�r�渫����"����Jõ�C;�����\(GvM ��)6G0Բv7��y�~����g���ә��<� Ǳ�����18�Y����x���ʗJ�<4w�Q�i��l�Kx�X@�$�>�z{��M��dt5�&�j���"��Þ�`�!�F�����]?
���!�b�N�d�
1Al���\�����vg���!���8��C!�1i�wМ���F��:?�v�K��3;�%w�U�!TP�	|�S	0!^��������cd^�%���0�{U��I�.�uD2i�_�>HI-!�jG�؍�;R#��C݂�3�kڌh�t�k����3{[�\^�͏�����=� ��R��.+��8�˰i��0Vӥ�f�C�Ky��vl(������Q6d���~���8p��q.��*X�α�V��e�*���4�Ԗ�v���v{P�V�]��!�$}��M4,�:��M2���ٶK`���}I��h?୷^�R�$"�;������|�ma���Z�t�9bϲ���H��S�� ��n6G�C�\�]Iί���Y3��0�,�||c��~���1� )�]U������ �f+\��?�Y��S�S�ݴ��m��n�z��)��	��<�7��}�G�ۤ[�a$O�=?���j�g`�#9mV�Kk����&ZK&��h��=�ADN��
֔�'r	ok
����k�$p�ޮ|�)7ͬ1��$��[�ud)e3��!Y�#!�WĚ���b�v�3)��OjN�E��=ݛn�$�8���Ir}�������4�R��=�ƙIV���[x���1�y�jgY�����4.ppJgn�cuj"����.�ر���U�b�hO+�֥n�/�e�P��7hu�Ku�)����4�`���%f��Lk��������o��x�2���@�S�bh�š�r�V�t8a �Y? hǏw��0����"��(���l��E����g��v|�1�1E{q0'41�Cq!����J��e�5�a����Ϙ�|6\�����q7�+��@�N��b��<�������m���yR
ء~�j6��p���vI���5�(6i� �w{6��gآ�aO�N&np���lp6Y���6�*��&�{���k��47���K-��"�Px�3�=�}�}�t1)򴃧INn�m��+J�<���M���Z�}�)e!�ۈ׳�o��o�}�jpQ�\�#� �.C|5�".%����5�v=�L��9�"#_	�I�sϹb4�{�$��� ��^���~��LgT"B�)����Nx��B@��\�{��xa���OR=� �N���2���ŮV=�w�D�I�Y��
��i�	b��Yь��M��Q�^�5�ד�jȂ,�����mt-*���v�,�P�陋������n�[�9�����e�L������Vgz�p�[z��r�
��z�(��f�`Į��)��~�������eQN7����V�W�I�G"{q$�^�#��{J�ҳ�X;NN���al��H���7e���р5�ț�+h�������U�� z�K��{�>Zw��O��&b(&Ȇ�(��k,� ;���|D�e��r"��S���T_z�b�:�I0W�2��
Nu�-3w�M��/Q!�u�/O�eii�}��̷$�.����8e�L����_|��*ԩ�I����o4i��k�<O�_�6/�ގ����rۊѽ�v+ƱP�!��;�VY������O���B��8�p�8����A�j��5�"�̤�X-�^ �U��$�rhȦtS��T���.a�3�ޙ��u�l�7�s��dT%�;j��\����Q��cR3��t�x,�U*.*$ļ!�m��b���������	�^-C��M�"�j�xY�`�}af����O�g �6o�`���Z!34���� u���n���zI0P���Q]�bX�|�Ɗ����TYF����<N�}Т:�O䲄w�A���V#8���*�Hd�賂#�R�#����의�z���?s^�H�E�$:�2�b��.i�M�ܩV�ixĮ�G�K]�\'R���f0ޭ�ī�-�*�n���/���=�֩�5";*0��Ǖ��2�I�Bh�F-����d���GF(��[H1��6}�2"3\]��E��D}{n�[��ٓ�}���qFC��dU1�g>��FtQ\*<Q��/���B���5�rp\���HT�/�)Ѹ�k0����]o���q٦�޷�_
���Gpz��\T���e�H����87�p�4�#j �J���$���&��p\����O+?7��3�g�Ѧ��%D�Xr��6[ I���`O8f7���Y���m�Wǧ?��`��u�1�Eٕ_Q�Dz#c�:.���y�����޳�n\����Ѳ�f�y|Xg48M|!sXX�ئ��7�樖���
g�D6B��������Ǻa��)l"��0�Lg�}S.d�(�g@FVV�)�NBڛ��xc*K�|���@��w��}j͜O�����A�} (��pW��
��w��:�r�C�N��k����z��
Cr���Ğ��g��$�%���UBF�_s �Q�y�V���,�Y��MO���ușӡ�n}F=6�z{jv��5�c�ZY�~Y���D��v����Kh$�P�([.7�b�=�:��K��|0}�+)U���7�V>����k��4����ݗ�]����wa5���כ����ϝ}LZ\"�6W�h�[��O�O9Âp�=����K����e�L:K)@�ǣ����{�)�n?�����z�ف縙^�X/_Ί�+ػE���tGz���s~J��.�]��	���0YO6���W���J1E��n�j�!��^(���ˏ;>��>��.$iCr,�`Tj�	h����L�����|�t8�e�0�W��Ű�
B�*7*�!�/��n��ġ�-6B
��Ig �$ �t��x�1��~�`�?���ȍ����@3_��M���K�nA��A�Xæ��/�7���
�ۢ�� .��魑'�J��&�����Ylģ�%!�y�ү7���$�1'/�=^�(��a�$j2D�q��T_��Tg�Z�l:���O���,���n�{�Ȫ�ϲ�VWB��׀V�b�]��g7�������(kg���8褰���#R�.?�o����Yj *X�X&x���j��:�2'u�!��zi_$aVaQ={����~ޛ*+��-�ix���yʅ;.��XN�l�r�'e趱HA�q�p�O;r/Ia�ѽ��/���]+{��%L�xA�X��������+�2o̓��ů�S��d�����r{���\��8�8�2�:�����W����O{�%�
��B�ۻ������[�ĭ`6 �3|m$�G_�9�|[����aD�0+�dNl�p��e�����A$�Ԉ�K�-ǰA�ך���jQ5��{Av��������9x�K�Lt"y�Px���yz�w�M'��i���{�_��l6�$2�<��E���/��FJ�荴R��7n.���>�Րmk����X'i�u*]��S7�6|�n��0�s�*��R�$b��9E=E��R��r���f �ʾ����癡�!��PI�(`�n;��� d�^���5�s&LH��"Z(�`I.����/��	��r�c'�
I�M���x����ѿ/�(�$�ku� F��5�����Rt��M��ܖ��O2���~�_p��"��Q� ��,N��k1���r�]
/����_���3��5ۺ�ٙ�� ���p�Q�@�I��g�.F�Nvp�֘sУ��8�D�Ӏ��Cx�8#���.a��K
I,�T�3�}HҢyS��"���]��Bz5�&z3!�������%P*w�Ob��.�������J��_5鼡��TKQR�-�K�L�O�"�s�>( �r��F�߀[#�B���@�Ϯ�:�������r�T�� /B�C�+�[�,�����=%��6-l���s�\+<���PS��X��h.#.��F��g����g�ލ)(�|eHȰ�T~�:�2�P���e��� e�-�߆0xnǦ/��j�q���͖e�!o�rɞ�p���Q��m��������s!Q�ϐg �~r|46�f�gx^~�x񺫯�g�vJK'��k�A8r���e��2\��8'71���)�A�3�Cb��H%t���N�F݂���|pV{�w�u�7l�/{����0�����EY<N�V�Vw[����F!v?�tpU鑞z�;��$��i����E�9����h�N�U��x�H�Aj��=.&��8�����4c�`@�i���4�x�>%����X��׮iV��ZOA�J߄O���]+Yae&�b��Cb �`x�#(�Rr[�ǻ�X��A +.���`U%�*���W����r�KL��7Ezun<a�!a��A�ĆW���슩�q+�Q�۾����i���ʅ2=PG������@���f�臌�<�v0�?�$��I(�@���F��g|2�\�B�2�Mt��c"��FO㢼+����E#���!���:�D��4�)���.�o,]k�����|H�DQf>�d�5�QΛ�E�R�����|�~��ߖߚ4(�݉��Y � ��>���Y@�j�N�����ުz�r}�_������EtE�����ܡڵ�?SB'��l��>+�{h�.�N���&?����*��``�������X�q��g"9��28���NMO�s샳����"����ʂ�~$���2���Y6f��۝	K��HB J���X�'x���p	�S�@�ܢԓ��M]�OB`6�S*<|��gI�HZ�i�S7�1lt�����]�Ad���_���VNg7
M4��Q#=�l�&�պ,� �-�g$���bh����E=�����iC�7Z3_�d�����">��D+9̔�C&�ә������X3,�z]��zt���[ԝ����9n�޼��u2�Tk�?aA������-ٷha����c�zБ�s��"|�ٚGdSK���B���:,	X*ˤ���,�$���;��nn���� /f�G��g���Zj_t�W܌>�+;۩��1E���K3U�j���8;��I���qh���lխ��}�.�h9fř$�C/����I���D�H",�6�+�+�D�Zxe�+[�6�N�!��o��c�\J�Q��C�G!���d�d�G�o����Ld
��{T�R{��K7a-������%��Kņȝ��W.v@�Rwv]"�-��������B���>��yy,���^��_ D�,~��1�}ap�N߿�Ы��n��Ւ��1��L�:����f4�,���#�o���)��V�Z:t�B���b�` �Ed�G�|$�0|�Zt�\�� �B_�p��8���K6�����^��17�V�)'�P�E;�dU��㕢)�4���x�q���7�@��27Q%)����.�j��֤U0��!2��q�DF��Ӈj ����k�3a�ZtN����
�mR/�A���GT�h3�$~lv�#���嫵�P�:��+��Dq�A��f����Nྭ��,���}K��6ρ���A<����1^�b=N�e�d��j��'�Y])�,�"Y�^��Ȗ)�z�O��5�_:�y�M�Y��끐�������>�bY��4�{���k���������{�YS����}bP�f�%�����+y�s!3@t +o��T�����s�R/&�d->W��ƉF���+��Z~��4�H���q[_N*�i��C%Ĉ'a6���@�g���F4���7��X@o��B��͖r��Ŕ-��'k�1��@dc[�.��[��	�X6��?kyIG�.�� >+��l����=���o ��M�D�^`H���HlB��ܿ��&ko.��)��KמEb��� $^���s�/��(NwPj+�c˲�Ɇ6�V��Z�A�i�!v9U�~������"~��N	�f�d`UnPhM&w�;��|�U����M3l��Ȇyo9ކ�c9˯�ftU��(JD{��[}�"���E��ܦ�j�L�݁��?�z�<�"Q�F=M.�yP��e�Q�Kr6�_Jo�A=��z�
���ХN�[�g}��ϼЕ�
zêN�Ȭb�>-�-�Ύ ����������mtH;w�=ÜRظ��%;��!Ԅ��Ncl[N).ǉ�5��b:9��ۍ�D������`�glXxS���p'7Z�4�W.d�M5��p�|��NČ��iCWk!D"�~�S�;��XO���I����S2�������K��#j�ڈT�%��310�����]�>�CZ@|%���\��TA	��熞�Z+������k��3�W
r���"Q:R�Y�]\{�:��n$��u6k��Tg1qq��D�{oV{X����d�������b���z)\'L��j�	.�o�ss]�c�x�վ}�S��UP���T�错mܿ:���+��`���UGqC�oK�6���,��� �Fn���r/�C�q;_�<HԬ�P蘙>� �$�9&��+�Z���məX�u�(��a������ݰ�6
礑# +N �i-�d����Y��� Js����u�%Wly3+_� �;.P�����\G�}z%��9�s.+cE7�O�B��!����"CFՠ�V���J.�ݢuY�:��g/�Q|��!\�q	�O��j����4$���,����Dm��ɺɚ/	��9q3���)�����$���w��q�cq�Y�"?�0�O܋�U��C ?�z��˄�<!`6��4����|՟7�颁�H�wI�� Y(�~Tm��M7�;�P��)NH�M��HmMÿ!�zr|��g�-9�D�}$�	[���.��� �N$I&	�����>�1�/;�4�v�)6�j��6.�.3�2l�f��G8�I�:h|�fƯ��D�A��4w���jv��W6�V�z���Y�t�M�zOGt�c�h�zE�������0�i�)�;R���m�]��`�~�����	��UT�c#e�(
���⊤�O�@�>�qx1"l��)MO�X�l�rG��v����5���Mc��6e	t]�V��"���L�_�Gb�Xt������vsE�E�d�n0	�e���^��{%�{^ؘ�U��#!˪W,K���>��:X{ٿ���v��mO,�Z���M�]Xyt�uYd�J[��k�OB7��&]@�/���{!���eGR� p��� zpm�7L���,�W���/nZ�M�aat��#��!�� �xێ:@~E:e��+�p��!u��n�-c��ٸY$R���6cCC#�+�J��W^��X;1S�wUX����\0P�*��`�HH�S�b���L�Կ\�I�B0�������P�HOB����p���V��`$g�vg�@#ELr��� ��K1����h��Աΰ�����1x|����.[�X���e�^刴�r4�)b���H$��I�왶X���,-���H�X���AL7���E�ݾ�U�-���\��G�SG��pg����.�Og0�C>�%=�ـ+���N�%G����N�A� �O|(�(C������'{�,�1��0�Po����\X/W�;���<0��	/��5�LjNa�,�|/����*��V����!Y�����?H����[�Ϊ�0}��*���-�X��[{И̞F��`2����%�Xk��؃��W�11���_�?h:Z���G�<���*���)�PS#I/���Ac2��A�'�#f�iO/����*�n�I0g'%��_� ^2� ��*���[�f�u!&�[��U� ��/wq�3ױ�p���4i�ej�j�
��:8蘒B5�K�4������1l��p�xpz2�6dsQXh��OИ���P��Wo�Ѵs��j��:�T��"�׋�Ő/y���,B�S�
����,��(ܷ�n��i���w�o�o����P��C��gD$�`F��j%Yg�?>�389��"v�5*�����Mi^ꐫd�:�p�,����t�i���嶻J�� 3� Ӑ����f��f"����VB {�������B5b��ME�I�nɗ)�a��Y�jUv�}�a!��T$v!"�^��.-o�n\�V�AD_�бY{��R4-�߬�Ie��nZ�ar���.\C١�wS{h��G�Y���2/���:jߦ�������N�MA~y��`[k#�@�����_�v\Q~�z��uN%lҳN��	6�m�������<K/�h��#b������bʪ�+�%^^=��tv
�r\��C��KZW��v�q?�>��X;�Z%�Ip�>|D�&�P5d�N��v���N]?�߹qt%-�,��mZ$�/��Ti�y��e��9�L�u���([q��^��o���57]"��疰����C�j�?�rQ3�yErZ����PVC��hx}R֨�D�ci����&}⤜̮"�]N��y�dy߂�)�Uy�%�m��z04�:O�I�<T/X����yI�oۛV��8��+�C|t�ȷ%����b���jy^I��P�`�#B�%_3S���0N{v�i�f!��_*�Ɠ�}w���E������/���(�t�{�KZo�<e�ȷD��
;�t9��Ӗ�ڮ�5�-6��}�pF��� Yd���Ӵio������Vo�%�}�Re.
���s�|c���%gA�pE�;��L��=����|kRv�����S~ǺS�~d3�IL@+,��5���қE�jfYN�g?��{-�k���#P�21j�ٰ��B���t�!=q�D�\�|9^�E�$)Q��T\�+3�<�GvY�y7�X������.b҇�eǷ^���2m.G�K��#&�F�|uJ��}�^
�q���{[-qѵ섓U����B��On���\a����*߅P3ū�'�2��A��E�V>����Rj�1���I1=�˯hS�8�oD~�W�;G��1K��aW�U܈!1e�fo�,?��P������y�gͧ���;g�VU�k���2ߊ�$�#�;쌙�%j&���/�����E,�xvdBΣ���ɇ� ������c�c�"�O^Ǩ[�����&N�eo؟��w)��t[��%�C��4g��=�{a�Ц(�1�{�v�R"��:���Y�X��K�.��p��=p^	�����.�f��U��6A�x%�Sc.-�Q�g4%���Y���`;��SZB����5�U�/�Az�xiҍ�9���R"طZ�u��o��f���cD����ԐY��%w�N�0��b]y?�2�gGe
@`�H3~^Z�^�>~�ܕ�k=q+v`�v�;�w*��qq�<<�9� �Q�1��=�Υލ�?0Q	m�O@�e�W[�L�HA�`�XPm�"��}��ש��@�t��Q����ǡwC�G˓$��\��^Մ�ŵQ�L��bl������2@��J�k8%�M*WӒ($�0
��4UW��d�����z���E5�|5�\&2��͢���5q�-�?�6�˻�hv���L�x0�D���fp�j�!��n��]���)L���$O���H��G�8�V�iг����V䮠,濛�����_�r?���C؊A��c%1?�7��8�F��_s��וW���G�IUO�w��Ն�ɉ����1!N^���g���d7���e���h'�7i���JU���06��C��	��0�B\J��#*�k���)���M�y�T������<��*�Ps�8s��&87����Ǔ*�<N�t�� g���1w=��>Ή��8y��Mmނ�:0�ׯ�{���#��
`U�����#c_�K�3�.S�8��,h�z˱^=d*]���ŝ�����Zm�I�c��X4�zn���;�4���"�M�"��9��͙T��ʹ�l�rx@j.�|?�,7�l���7LC�/ى�x�w�&	뢶99k�]de�^u]띣U>�3cu�{a^���b�x�������>d_$�^G�R��o�"�'L
r!+R��9��Q�O6&�ia�P�
9Y�����l��6��X�L�kf�$�B�����wa<�m��#�q<��=y�b�e���]�o��HsQ�t>�{<�F��Q�~#�#�7 �=�=�I�%�`�~Vx3.G�$li��-��2C!�P�ُst+�[o����*�F(��{$H;��&��~巻=���D��h ���4���,b�Vd���o�6>b<v�?5ӕ$)� "mhA�*L���d��錠[E�� �Wb��+xn�/lWRfX��G��_ށ�4��D�	�Ο�
&�x��˷��c]���O�F߱��4	����*��� gu��)�$q�rb1��V�pA�w'3Ѫ@팦(t�첝n�}s�|DZ�ewj�j��[�OY�>��up�u������"�.�(!��@a.b��X�tQ�Q�8/GE���SA��5��J��2%&�0�G���MO�D�]�r���D�9��)������Oh7�B�bK
D�:6�'�9�:�Ɇ����{?H��R_ l��u�R�BQ!8�q"�0*�;�0��`�q�˿��<�u4��-��}j���9r�U�k�J���V~q�}
�R؜`��>?_Dџ��%To����Vg�Xtd7��|������GA�ʪ�&}G�ڕ���z�%�۷c7��)Hؾuz��ѯ�Q���Ɗ�<�ǔg��΀Lr�.�tGl�}��;R^F�o�#�F.^f������c�a���9��~�Φ��\C,~,�̥��C���.�fa���@i�����k>q�q�Kf�xD0����e��Z��r�Whڠ �:�h�R�J�[�Wd��K�IF���9���ԁ�}z�QO����y�B݆�57�P�o�m��a��[ �v���q�hz�yz�r��۝�۝TA��{�@I�X�k`Y�w��Չ��z�O	�����ceT>��i*�� �9#��h�Y��Q�v�Ԉ����뽇ޚ���
��i����W����ȓ�N�J�bnl�ji��O.���E�fk�*D�@��Ã*�>�����X�� �?��w��{����=�_9~,�%,&����;��r	�+�9���;� >��|�]c�M*z����sq�o��D����
斏>�	�x>&���<�Q�G���p ��;Z[M�L]i�Rt������[�k���2az�\�P�oQޑ2։8l���t�KV7U�P�a�Б~�;�A*�z��B�ʎ�pWUA�>�,��1<�@	�g��oC�8�-貈m�zP��$a���s�G���
�p�s��d�Ð}��I���mJ]������
e�$Y�lb���(O#E_�o�Ƒ���%vZ�iPrC�HϿ����n��5���6�<� I���E�����|5S=�/�˞:�p��B�-wLN��`��q"�g��{ia�Չ�^�5B�]V�'�KGwx�GQ/��o�uOC�>!�yNq�đ�q��~3r���k/ؗvf�*(�]��3������&��'K���N�c�2� �ۺLQq��6��WQm����0V��4���O� '���C���P7�M�V��G�q��E��C=<Ʉ����V����:	q}L�,�UA�9�m�`(2_��l2���5�ڐ��\��rȢ����g)u{����7���DA��q������mg��T*��{���İ��,���>(��Տ#^p��v�dS�c�X�����qy�DT�5��3�B� �g�4w�jH�2Ƭ�K��
e{,R����ֱ9^�1�^͹�Wc�I:��]���g%%Ŋry�S�^~mi"�D9���b⚶�*=m����֧�T��m̀@�{у9WZB��&ܜ��PVQ���Ρ����"c�u6�tw�8�d��O)<���tݔ<�;0��G;�iq�UA+~Է�ih�����^x57?j;cBc5EO	�`�^��:��~o!o��^�z<�����+�Kܢ3?K���L4<�.�L��h�7u2@����*u�5�����C����vX
:nG�[�\?��v�w*�a�n|GO��4��HJ��!��Oӎ�������WA���1@粧���&�l��V�Kw-����Yk�@�O��ƽ;�b+"a/B���T��]Bhd�Q\Ѡ�����j�a-3L��Ќcd���{�E����a@p3�ΒP���h���S{��]Xlf�a�e_�3��rLL� �,�z���v��I;,e��ZD����ss��Z�ڥ��bgo�Ј�(�p�o��G�>O���1�����2#s�}�����:�=F,}cd�	l�*��y���-�"�Z���˔���"$o.�:wZLu���bX_(-@����3��p�����;�c������F��t]�=���
�wG��;�L�jޭn����b�x�(�t��Q��x[��x�t�!��#�k�5�	)�eFVO����z��!�.<N��b���*	�W*a�Q�Ԅ��������������rxf%۟T�	x���#���]�:��h���ѧB4q����8�>�z|��&�{�N���p���M�e��G�/�������I���4g�x��t�խ�U�e^[]h��Z���(��Fӈ[�MO�d��7�0�[�#d ~BɔL]0z]�F�0R�a������+O��n�nOR��ʉ�GANm��Y��媴3J�����Rt��91v�.g�F۶m{QSS�Y�2�
f�79�~�PV�95�[�"�Х�#^��Ö�ln�Hh�#�"�?�xr<F�µT�LZ��IMRse�6e�4P�E��rI����svt��{��i����v�q Ȑ��ޓ�i��	���܀*'���|�(ô[7�Pq`�*&m|7���x6Ը5�.k�Ů�dXF��G�q. N����:L5�ԍA8��(9���P�)iJ:�������'t��<���X��.�郎��O#�^g��c%N��p�Ϻ����Ra�^�U��5b�B(�W��n��,�,�����#��m�u�q����ۨ��g�66��XU�ߦ���ƀ�ZH��3@β��M�O,�dZ��^N�� �{mNL�O�`(�?>K�^y�?o�<����:����]�®̸y0@a��<��|��%@�� $lś�j]�R>�s�%fގKg��������g�n(Co��TM�Aq{�sP�ƪ
<�OO�zH�?�=mW���H�۬?}�y��(zn�`e+lÉ�p��&q�	�^�a�YE�H�]�T���Gֱ�N��,D�V��<����]� �(���Y!ut88>�=�2��E�~�i�C�a����t�p�D'��}��M��&��U��)�B/��<������ck낶;5��2��o�#D��N?����ڣL۠��<�C�x����%��܌0��g��)
l~�a\��������TV��Dr���I/U� ��ψl��lS��1E����<�FWǃayՁ
nP�-`z��ҧ�[. >�g�+nXX[�4nFѦ�h}/E��a�ި�<���c4����������9"�E��ٻ��bJܼKx��A&�5n����p
�8���^K;�Z�d��	���a��6o�LZ�y7��h��{$��򷯑�"��xX�8��(ݟ ρ  H;Ү������X��b�%�	]�Qؖ�~{��F0V���0�3k'<`��o��3�(q�cF���x0�$z1Œ�ա�Aɮ�Ú(�QL�t���O#AMR���g.�� ��bSΖcd�=e��F���A��ܣUH�ɮVz0'�iQ�Ӈ��&��D�\fS&o�yɈ�&����#x�w��;�I�c�O�η�p�J4 ;>+���\Uz�=��l��8;�X����Z��e�c�'��<��B~]_i_.��`�[Q)�~vj���
2J��:�1�Nt,���hGX�@0,ت�l��SA\