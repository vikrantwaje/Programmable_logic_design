��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞���Q����90�mUe���-���W�������]�~,�ð�r��>�������$S..�~sƩ׫���\}����ճ7x5�1�V]���V1�!ym;U��[�����7�*oS���yώ��l�k�ů��m��$T�!�<�B�����2�4�8 Z�?+��fUb��6�4�2�x���T�-4�B�N��k�l��[9a�akf���
f*4,L��O|حY�\��W�+*^rK%�Pٔ;N6��޷��qnݢ 4V��Y����� ���E�GK��޺�u��ܽ��5�H���[sM3oy����k����_$���C�w���|h�^�6�|��Bq[��Z��ER�$�?	Ж�u�)-W�>�G�* �h��f�1۶�~�e���Bj�{!m-:�����H�3����x?rH�rg`6�-ʼ�-��1��NqגO�h_$a��':D���d��%8���\�zM�"8���P��	�e5��:6��Y��~��GH�C\��q'5�W,�g�pn�-
q�q�GF�G{����'���z	����
�+��R�m���yY��x�b垵���=Rh;�Zl��W��t^���(��s�(�jJ%n'����׸�9�$v)���t�{�W�Q��iX��#PQ�y�n�/=j�j��A(�4�J��-Ӣ<�iE��Tš#h�/N�c���`��6�"a��� M����
H<.��Ѣ�v��M�r�.N����
��@c�o(�u��,�X�ad5Ҧ�(��|6�9�t��{��\Ph����.gfv�k�Oo��%]�̻F�Ս��¯gN%�0twO�BVģ�ٿ�I�̮-�?kk�B�QC0�^����
��;�޺�g�4��u�㛰t�M�e�f[k'����6�u�G�� ������_��w7F�U�����e2&[G�����	�ly� A����g8A�� ��t����//�ϣ��	��U�H!8����Н��i� a��a��@��x��]^.=��F��C��/�7`�\-�I?Z�!Q����	�)�A��s���V�����G	:��l�%N���x�6���M���3���d�Lw\E��\˂"�}d]�qj@�듭��2P�q���B�o�%���B��b%��������ԅ��&�ÛI��}�?����*��Y�u�k< Q�(He�}��}�	�]8���C@P�X��r�]�A8���*>��,�ۃ,!:�oY�#�?E?����XF}���	R�Rh;�Q���ꏤ`-�P4d9v>���\S�i�؟	�����Za�q��֬pY�U�1�D8�4e8��dsWq�/M8�U�i�G�,P:j�%�Q24�<hn�^l!��ځ�>݌f�g~�P:��צ9�r\�ʈsi�N��G6�+��yb��^m����t3\9�qv@�
�K�.����g���|�:�n^�2D���f�_��fJ5��9	 �$��j��U�+A����{�g�p��1x$�!��%e�?�u �d�{�<&X��[�s�S�3A �	4}J��(�W�	�(�P��π��/�RKz��ݱ�\�s�	/��Ns�a�جJ�]с��N+��s@jK+�D�*˂Nq�
ɠ�oOJ��<���Vۇv�������q��{�pX,�؂ ����4��x��d���y%��&�?�m�`c׈"r�4���h�&����o�,�x�E���T�fh9��H�ą�m���CT�=�	�A�D��"��`�qe8]*O�O��ZR��ǈ�^�V����\ئD]l�᝔q8�ώ u���d��X2�,���Tɣ�C�'Q�D71u�J�'�GIˤ�'5#�m"���W��a���~,�����"duu[�ڟЦ��xbQ�~9z�F�����^O�z[m�}0������l��u�_��u-���%2"�k����5�P�Ѡ����C:a�������W�?�P�O�]������KY.�~��h��1g��xG��5�L�:�
���4ep�?��2R��T³�d4n6��S,�v�W�N�����>�_�Lfq��`~�b�`ލE�Ǝ��_���i�� �w!;(|��ukw�5$�p�Y*�T>�h:Y��j�z�!��[�S�nF2����߫���N ���$�u!.6z�rr;,�棟�Ʀ���h܄�ܼڕ��q���w#��LʶDb�G`÷O*�͠�s^�[셯��$2�jbMj��^K�5qL\��ŪF~�B��N:�B9�Jk���$^�(�N����#Jq=����$�ō�Q^�
w���w�����5�zϟ�>��֒	�u�i�2qta��j�E�2��̇\i _Z-ȿ�VyU$�r�Y�փ՟�ɺR����4Ql�K#K��ֲ�kT2n�ʘ�����阭�������ks�@0Ja�h�z�x:�z�A�b��Q���֮у�b��*��D�h��;A,oK}�^�A4�k� S�O�K7��ѓ���0�����<���Ę*�����.��u��{�2�o�"3���?�do6jP���{"S��/送.7z3Ŏ��L�vm�R�b�f��x˸6Zb9���(���1ۺt��gF���&�z���d�q�bXq���A߂��H�S(�����!� ����� &w�O�5�S���Gee�[�V ���,���7$��=[*#���PmL�9tW-/�b���C��l�2͚\�S|���gW7IP~5J~R��s
�t��9W݄c�˰D.(G
��?UUI��jB�"i��զ���7�n�Y��9Yl�o��o��J*��� ��#��C�� v��1rIa��'��0/I��!�kQx��un��w���N�����F�Bw\��N�������댊�3?R�����wq��| Ǫ9I2n��,�/��6?�b|ƒ�Xa�@�v����V�����1؉��62����VZL��@N�'�D�J'�qQ�|�Q��"?pL�ؼ�g�o�������O�-�lB4����]7��0���w ��jo�yvϹ���mM��!�63M
�ߖu�ƞ|Rm���[�������er��]����X�@I�G���|3��FrE8���-XI�58�k�$��u�vr'���Iwx���}��>�t��$�^���g9I>{3�lC�=�.��&��	R'���z����vh��<�\^I�'��.09M
&l6.i*��1m���w�2�5�)�y�������pFNո�FtmO2�e{%�c���@	l\��`PD)�u�A��%��NV��}�� �ГcI\I����Oq��t��tx�u�Y��L{_Δӵʸ���
���]{�@
"wư �ܗ�&��&�oRݘ:��"�h@.�4P�dz�W/Y7&O2�е��F�F��c72�"6%l$I�e+�L���N@�Oָm~RQ��;���5x�U���|�I����n��$%���4��d��Y8C7����5	����_煌<���ma|�/M��ʼ�*N��i��+=�g�_�eD���ic|8�Q[NƅmO���G{�^B��/��0��v3vyv�.��aU�!+
XCv�u�:M�W�>����Sa�����o��pg����R��7��ӿc�t��Z��|T��G	��< ���M� s�r����.ɠ[�ہ��9O�&�{<\���Kt����iF=��/����pA�+����l�C�J�}�b{���g�c�.b8�T�	��uѩ�^����8�q\\W�?YSHx���/�Ǭ�%Φ��XΕN_䪨�OG-=D&��:Z9bjl�q��K7�i�ɰj]�`�730]]���a�<Z���&�Q�v��'c�ֵu5N��s���f�6w����T�˅ ����Es*�����2��_R��+�=Z�Ei�(����1Y4~� ؎WaL���N�K#�g}J�K[�Mu�j[L� ͸�W�W�tk��V�h2���n� ���|�	���|.WH;��c�f6=)��!��X`��H�`�i�B�5a����v��F�%f�2�a���Uo�`X1iw�gZ�K��L��p�'��Y{p��6�2�z/�X�ǻ��Q4Iv��a�/�p=�@��kn�m���+C-���h]:�t�fMI"\��L�Y�V���,�GC�g�G&|K�R�o��]\��%p�cdSV@���� �rLYay��ڐ���&tk������:\NE�a~:�Ą�>|;5��E����fX"b�i�A��YK�K����3�P��`�@���z��^/���=��u�;����n=N��?�{l=����&c.Q�Lc�B&f��L�,��w��S����$a<�f��k�0����S{AA���F.%�����}�h�ףpq��,j@�� ���]s�ٶ`�ɉ�@��q���Rh�>_�o��Ô�ӏ'rF�֖aㅩ)��E~)C/O��$��]����@m\� �O�r����f��ۦ�Њ��;߁�.��-�X�M����{=�咑5Z	zs���i8/,��3�zn��_�����9'%�m;;l0�O�dH���^�ԺB�%&=Z"��I�W�>��{ �+��XZ�9&D�L^n`����Vt	fF��]�7/�<�g0�^(�w0'��w��na��j"�Z����^��]4��.�{\	�.�S��P�X,�l �x��2ya�E%��*�%�enY�i�����p �x̥r2[<�3�,���V���+ɚ�|}a���p�g�T%�ɍ�/@�-�s&��u��9�]51y����.�ԅ�?)�S���0�`�V��%��������A��*������۵�V�����%KT���wh.^������_���X;`�oa}R.��م\��#k����v@<j]�+�,��l�hF�k˳b�q�����	Y���eVGK��dm���hkO;h�"WݪE6��52��Ƹ�/Y6Z��-�us�?�g�1e����*��O�H����jN�f�:�Xk&?/��Q(
�(��-���5�����sm]�}$�[ż�Ud]�F�i>A�]�g�K1�  ��f�0��߫N�N�{\���|�2th�{�
�%/X'):%Z �G����E�U��9.���\p��HO��p�� �ޅ$��6_�~�a�z�L�Rx
6���D���\�����s5Ɯw*����-�.�Gv��a[����n��2�b�/<&R {/�ĸ���Wh�e!���g	:��R�%s���ķ���Ķ6g`#�B��3�t��*���2�3ks!��d* ����-1��]�xd�sQ�|��[醱��(ƭ�Z`��&҆X�(D��>XR|���3ꇣD6�X�E�)݆��0�҃i)��b�V+H ����mሡh|���u��� B� ����;�73��,o�{�\B�}�J����v[�~��7�@�ڳ-��&(��az�[W	LRc�B�����T(��<cJ��O��rH&�$?����/������I�X�Pɾ�~`�Fn��0AKw?n[^T��� <S��r��/��ߞ`����ZO'�m]�1@|"���V������Lcqeߜ	�.U=����0�^���
hMqRbJ�&�ʧ�p<�9;����{`�ћԬRmA�hi�t�V"4Π`�~��M�S�R��ddڶ�o��rǓ�Κ�X�`����/"�$?�R�/�Nui����S�(�$�y�����֥��Db�>25�S�`��`��s��`���^�N�ٟ�Q���LK!;�|m`ƴ��"���0C�Z);��?��ԯ�u�p&�-=	����Z�`m��.��s�դ�t�oi/i"����1c�aӉU�T�jDEυ�DPF��0�
����)��P���.�$�]P� �e��Ј%��w��;��XSY:G��	f®8 �䊙�P+1e��۹-zd�Xv�yL:��h����%�iҚ2\<5SK�]��K�>�f���i8���^�T7~�<%��z�o���r���Ve�/l��*@b����+<�������1S�Qײ��v�s���