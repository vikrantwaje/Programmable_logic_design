��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z�����4��������8xT�(�h���/�<�F^[��V<v�Lz�=q{���ˁS�=Y��y�
��+J7�‿��(��ߑ��gƄ���'�j����/��b	 ���5��G��r>��T�CF����Yf42
!zEKǍ�>�e$n�i��F���C��T��:�/�ig�Aރ	V�j�e����@Ȋ&��<�RL.kD��JQY�q-9c��|�e5�P~+��q��ͬd�[��@�A{�����'���瘅t&�rX�����A���qr�7靽d�?�٪��|@-X�
�!Ȋ��88^��o)��n����gF��}���5��ӄ�Q~���afP��D��]�h~��؞K�Wm�O�gE��]
�(���L�����pi�d�b�;R3�! �yR]�H:r�T��Z�w��G
�-�c�r������h�����x�{�(�7Z���I�f<*Mל�~ȿ��B�z3��P��Gv����^n��x��D]LԱYi�Ž*BX�`m�gg�~Ê����4P�-��"cF\�$�i�Dؓ ���VK�Y,Q�R�WI��ڍ��!�ˑ�ܿ�lo ����O^�v�1�e���u�~>�5PgxF�.͆�G!�FL��UW�e�F-]J�.�ƌ�E�4������.�^������� ��;��֏ٌ�LsR� ����`�Q�#mb�]A���`�ED7��5�����H�6\I3Zp8&��2vKZ�/�N�|�,8�-�����B�����7r�,g<	$�t��o�k���֛CܢI���;_������~�7\��F�+v+H5ט�ԑ��*�����
~OP��;�VQ� f4�!�{�WB+�wtj��U��0㭉1�ͩ��5�}A�{��K�����ml\�bw)<E��3�0��ҪF��OJN����ߥ�������qD^��Yr-4���"p�/8�Vf7nL-��{�U��-@�Ӕ"��sh����ޭ�3�]yW�Z�쿺�ί�-n|�����T�Q�v�J����
�a�/`)�r��G�̲q�~��wi3뀖�:�G���t׍��814O�-��3g��X-U:��)�����V5 �>�H�Exy�M��T����aeJa�:94Į�"����b섔q�Szd�|�vQ���0W����L���D
g��3[������%����:��u�v]5� Z@����ƛm��?��s�R3�ǔ䙹��ű��ي���/CJ�K;���[�5�r+�/5L30�mP}ՙ�=�&�v��,��<��-Oq�l��(��|��!K{��ƱXIQ>v�+�B��Q^\�Q9��i�TSqփ�'���;�I��k��_1.������
��(ƽhʳz��QbZk�'�������=x�C������N"�CY�EരI��[�8��x摻~ѳ{��؊��"�t��4��|�z��>�x�� �a��>�9�)�#��j��T�f�fP�C^�[��6�T�xU%F�pH�?���W�TϘ��^4o�ב"�mx��|:��o�H%;ۢ��JU�t�L1��diTae�i�8��⛏���3�%��%]��2A����+vc@�0��Q�j��Aq B�{~����(+�
?^B�+�� �dJ�xq�z�F���[���^���Ü~��<=�r���0���u��ce���R<Fz!MQ�?����:�S.��*�j�i͒�pI,���ÖC����詮��nxT�zT���8��<���t7�d�c���@�:A/��zn����ı���F�6�z5����9�>�e[�IS�;OT"�d�(�C�Ӎ�X�&�f',	~��\	lo��7�S�Q�~�[_�?30i�ϙ6|I�o��P^�����ɼ�� ۣ�g�����؈�
�L�Yl: A+L����3z
��`�=���k�\��v��F��`�qlEO��o��n)g-3�w-e��l��jE����&��s�PE���D6ù�)��+hZ�1�� G��%5�FH�\%:H��}
z�+�>h{�(x�fc	S��/�Ꞧ(κ��R�i��f�}�^�u��;��LBO~���yYp� �"W�|)�!�����f��-�Z����?���8�H���+�L���B5=]˯�l�GK
(I��|'��.��	��^u-�o-��o2�zSo�r��:u� �k�`T�� �X��B��.��|#@�$�Hr��ǒ��ٍ��)�>��SU=F{����N������O��r�&�?(��h�����SJ#��CI����M�`�;?2*���a:��!4��I�e���6ޖ�S��0gX��Ŝs�x�Gǜ�ͩ�;D��Zq��=rc����PL���}����6��1���E�.g�_�(�u�Vk��%��4�n������$��t�
ԕ�I��� �H>�H��ŕމ"�l��S-�yƳ�I��~��&{�
�5���.7 ��VC�/�H�b#��ܧ�,Y)��T��F^�E�r��&��dn�S�p���*κ��d�%��!��
Q,����}uo�H!a�P�+U����P��\�����S���kG�S��<�e��/G�op�2c���'v)�=A'�d�*3�g{�3�	ʷ^N�s<��5r�c�$)8���g{��O.OK�l�Ą�׃����(��F��dx���>�}5߾$�F�zDE�=�)�ϵ��*;��*�+���Pp\4���B��s�~^�{�(���+�Z\�����E��������1��#�$Ԑ��bV�d�d��\8Gt%	�m���(�c'�\Ȑ$�CdN� 'CVy�1V��Z�������ݙ�VI�v���i�����o�ZLav�P���)`k��,��}���#W&���((��;����2Ul�ѡ�Ck.�h˚©���m�>��!�����W�T���\-�0?�h��b����A��I�i�qɒ5��*e�4������w�B0��Վ�bC�6Df�{�O�r�kW��-jT4���p�^ݲ>��%
A��X������j]y�G��兙#�#2%?���Mj�$S�r$�qig&���E��=�$)�)������~�F`=ϡKى�Z{�	�\K��xoa��.�&o	�3~��ʲ�#�,>���=]�뾡�Zmg-����X��z���}&^��,*'fLT�2;�<��qTf�Q��9C��b��GV�n�$0e<��]�X
�6��ˌ�Z�4����c����ob�~۳X���W�̢���a��������5�&�&6ŮyQ���PɈM>�1�q��)�pO��]�|u�^��>��[�Ԛ���T{D�T���W�t�VQ��M	M5�b�9Gl,!�&�9���yUr�����Rt��\m�9�[n ��y5�ۣ�{ߒs���zc�C�`9�\�*�SY4��T@���cf>A��<��fƽO��qV����p��fkUU{f����и��#����}]�^<Gdo݁�Edb��ŭ���q������(���y�l�`�h�I!��D
W}�I�鑀Ļ�4p�l�*Q���W\����Y
�iHg�����8�V�GXn+s�)c1S�����T?���,2��*X�׎�F1���=́;��� ��	�>�.��m��*y{]Vp��.Jg��f��e^@���4J808=C ���?,�v�U���̆&��%�9��G��`Nv�?�x���
���d�*q�}�w�I��H�RJ{�꧸ f�<�q�3���ō5=�M�Z�OW���H#��v�E^Wʵ&lQHsY��±�541��F䈷|t��0,Q��=���t��:˶3�V�%�(m�u:rqg�������C��G�>�ԕǃw��k�5?w��ʗF~�`3�c�G���(��4��r�R��KkB.'�5�B�P\��0��Vft4��ݵ��0=�!T�ٹ��C��q~�v~��\���V���F��+U�s���݈^6q	��=��&����-f�{}��f��?���<;5Fڢ�/;�3��?d!7�
��dJ���u�h�:rD,�a��7�O��j��.ۮG\:����xa8>����^�X8�c��@��$���gƿ���p�ܬ�K�M����lj�����ю6��fyl7 �v��-	0�ˡ4���?%�&骓�r�7_iB~N��4k������y��:9 �q�h<�/S��]��Z���/�LC��9>���5|�t�G#sjW,�E��!�6��?�A1�'2e���AN25�u|�1X1�2�!��)�`ț5�ć J�'�$�AUlBe,�UP�,F����HA���J��/�:u�E�\�:���U�aM}��Q�X:Яfi&J��Iq]ە�o?�c�YH�?rGE!X��̃�f:��r���ӪD��4J����bP��'��D%�p��,���,�*�\b_�g�P�x5�q�S�֌�A�t6��\��[�r�<%8��z���ώ�1��>:�4߫�1K^ܴJd�m.̬؞Y�R:��EP�i���\C*�݆��fmf�ۋ�[�������P:�D��܉��g�W��
(� �#k�j��o*qJ}m[4�,S�I��Vؑ��C����r�p��I(q��N�izc���s1�y���=).n��V�Z�?���r>���Ϟ����x��'�Y2�,����p��x o(��\��^`Y��SMeO4l@#+�o��7�3$f��Ì��4q�c��N���9S��l��M�R[rH��e8:�J�kh�]Y�����L�ѪpQ�g/��0���V8��'{���&� e��ݪ��r�2��*s�۹��$�	˲�|�M�|W�-�D�¹����� Q2PO��ἥ�]�JB��(�*�����n.HU*0N�&����m�_D�M��ݳnU��c�V������&L�����O���2�4���~�����eu���;$C|�T���H�ݦ(C�=���@Z^
	�c�
\S�x0�Lf�XԞ�f�~"�..ȫ%?��2Y����M��9�}�fXC���[V�hSG�X�[�r�V�"pH�U^5���Ŷ�����d�H�Z����bBp�I9*�J����'j�����?CQ�Y�:�bQ�w\wv�=`}x�0�g��suk<�d4�.	�Ol��v����;���n!�nͦN��&��)t���b���7�7��ڶ���&�d βU	���yU� YW ��������&Ҙ	T���H.Ȍ���(��z�c��x�H�4*N��5�;�5K��/m5�����b>QQ|q����:��L�t��Nj�68U��;�Z?lǴ}�p)!G��PV�!��
��FM��8�T�:��άՂ��I-��]BԊ��Nr@����v�DB�Ԍx�P��6`��꒯�ؐ��S��[�3�=J���r�8ӕ��%߷�w�go#��ko%�P�'�_<��U�yc>��:o�ٜ�Z���\_��?��R���1���� �X� ���6��X�YK����jW6�F��*�x4k�
���e���d؍�݋;�*����^M�C�b�+� ��0=H�<�\�o��R�+�T��Z�^���~�u�x��A�;8g���=�w�����@��HBz��`�B4�0,��n#{^_H5g��-u� ���?���9�-���2���/m�H
G��w������
&y����ȉןs���S���G4�#ua�u�X�����F<7��V(�̴�d4whu��?�� ۢ}��W��N,�_B��|&$�8��:�o�[��'�,�~��L?�0��4l�E3+��v�G!�O5`�?)ۯ@�?���}C�r������g�*���.8�>�����*&�T�:�C�߳�J��5w�}sB��~hYE~�t�]���`�o��錈)t�F57]0����ׁT5`ό�Y���e#���m�"��T�4Y�x�m��,}�$g���ʠ8��?�Ʒ����y���b���o�>�tk���pI�IpX�4�ӅX�*/[��Ss�Ba��4����l~�I��}63n���:ϣ�������!����6���D�e���%��^�E�^�ia�GA����+��ZTB�ݫ�ګ�g���-7��Ź����~��r�ui1��?Eo	��N�W1�-���%�w׶NΎOP��(O =EY���!���=��'�E�kV�D��<�|ͦ�
�P��4䙘��'<Hڼ����:��Go�2��P�%�o�8;K�|��b	fˇ(rtY]�K�1dXy�j��T�����?�U0.�X%�'h��T+D!{�&%A[,��8��.�4<����佘����Ǎ�zp�[c�fFB�x������K��&��u2q7#�4�vk���X�p�Y���^kM��W����c`�I����`�,h@�s)~��Ր���v��E%&ݽ��x4���U���i�Z��z��RsAv���d4-Y��yiA�Q�����%R!偒Q��6�Cz�$�	�8��Y�S���)
�Z�h�U\�&�����A��---���N�9T��-��M���C[�o�����΢5�ƈ�^1ԃ#�O"�~F���J7ݑ0p'	1�[f:�{��4Z���$C�(O�'@�a����C<_+-[��z�x�����Z���2��V�4
�L:o¨y�:��0~�c ��Pu�U_�e��_�3P���M[J%^]SJ'�WK5��ť[JnL�Y�ϧ(������V��u��k
X��7�wS�=�g�4���xq��e<yW
����@8u$�d
�y5��X�m/�݁������檨۾#����)�<�1
� Z�@S���l:�8=��N�H��&HF 7�p��O�%B�jIҾ�ʆ��Q��vXc�oVei��,�?F
Ĉ�6w��8�o�a�rñ�y�/�W�h$ S�MP�"3q��j���]5��u����1�xg��"]�>�B���Z�!)���������%���ѮԒ��=�or��@�)�r� &�ͮ��?������gR�G0���)᱊@����%;�e����y/�lNӮ]�����1���#�~!s�C>��i�'u0^�K�2� 38.�_'��=wo`/�ec��HiL���N�f>�Z�Z�\��6�0�"��9�ʒ�{�k9�6a��2
��h�y����*Ey�����c�O���`O��ۨ�S��U�
�%~Ől͟]�f2%O�o�.���|d��c����{/�mņ-�MXP�tU�FJߛ��=�-���9��N�\�p�vja��CG	�F��LujU��Ψ�9H�%T�!�	-��n-܁����w��� ��1w��rl����+1&m(��=�!O�ɣJA�M^�S�Ѧf���dG*)�	=m�5�B��b��#p
ኄN��s��]{ջ�B���� �FF�<�ϑ�՝�ц�x�ݹs�ڨ�k7j�*o�hY�J���ZdO��?N������1�W�#+7��*��L�x�����\]X���<��U�4���Ej��%��6tp�|޴������uo��W���JI��2b��~��l��$�<�j���Z~�)����5Q��:�q�:î��1���aS�v�H�X:
Ț�!מ]�$��"镽��Sal��kE���2���Q8X�Omi��1km�7�k����{c���Q�%O]�W�`/r�cb%"	ѕ>�|5�2��*�6/S�h)�hא�#�H�h&�7�a�j<��Z���ߍF^@.�ݞS�X���[�rH������VU@�;%h��N8(c^#��0��Kb<�ݰ�������{;R��7r����-]lF7�猏ЗM���M4^=��s,��B�����~��MY�Py��&to��a�NU]�y�f��%���yR��9[y�����s��Ѵ�����wHM�&���}d����J�ɴc��ZchB�o����֘��M���U�a'tɵ���ђ����'�MfFʜQ/�E�,� ?�!��X4���WY1���!A*Q������Ꮨ\|�"�2aS]ԝ�
����]��Rjc�4�%�Wv-�ƛ�����_Ue�uS��"�
Yނ���Ńr��h~z��hL˵�D�9J�FQ�w���g�����w��ҕ�R ���}��X�+b���ԩ��^M����H8ɜ1��6j{Ed��s���*c(�ѻ����O�Yޅ��N4����ʖ3V��Gw�#�M����,��+�=��+���ǳw΂����~���a�����g �� ��l�`�����FM�0��g&$�yo���J�����TC4���a��7��c�W�G�< жT��h�E�9�y�F�_�=��`�U�y�
��i��O��byy�Hf�-��7��:��(_,�E��5:w�Pc!�os��-�_n��q��e���i���aAקI���;,�/�4U&���4%��\�'{��Dd�����PPn$u�e���!6'J�*��)M7r/��� R��q����2��o^ᚔ��ҧ�
�2�L�#�hc����&3���I����Q��e����@�E�I��%�}�1��G:�#(�O�
b����oGM��2X�U�)NS���6K��U���ܭ)N�֖���$� ߞ�>�au�q�LS�aЩU�]��z��}Q�hrRe����[�B�cM�ؕ�L�lpg����A�*��\���~��ƕ8��bꣳ�WJ�;�j �$�|;��2�g����E�=��Q�@�pv<�����/=(���G��q�L�����У(�'�1A�4>kHg�ҵí2��>CV&���/Rlbk�2����X�������ο_;]������G(�5<�)l�F� ~��<[Zf��QZ��*WzF�����&2I�ǝd��5}u��a�R
׼�ĴS�,�����P��i�]@�f�}��'2��o'�6��k�ہdyM�m0rDz���Y�
����V���m>!赨�uj����R��."��l��%��E�3t܄�_�#�0�2�$;��zy�
�xC;�UB�������6�������j�%���4�2�t'�ʧ6~�g�\n`��/H�q�1�kj��z�r�#6H���|ҡ�8j�j�3�E��(n�$Mp/��D�NW��$�D�����W#n��=��\G�9~i,�a��]�)�/́:���H�J�����lt���{#Jo;�-��/2��q�G,)v�`0����g���u�K�rf^�ce-�tz��]�3�j-N�u�Sk�FA�M�����t��-앍z�� ������SU�����^5hOdsR��R���_L�Q��2m���Q����p�5�jdq�ň�z��w%q�~���mO��`cW#��P�m9��32��؋�|����>�ˆ�/-A+��?:<� q�a��� �|^ǋ�I�\ߔ;��ϗ�����pC2��$���cn��e���wW�8�)S1�����{�J�q�kQ�a��d����
��Z���c ���']SY�Pz��*w�N�C� `l4��>C>~O���% d"�w�K	��&�!I�>�ߥs/������Xp�\'���|�S����f+�#�G(#劑+��p�����i���v�̷�X���� ��R�&w�C�a����$b�;�V�2Tt�GJP3 6� ��?d|��"�K��ѓ�8��Է�J�����p������p���@`V�툏}3]�`�9��
��w��'�KQ��6	QBy~]��زq�B��O��l�9�^q��+	ī��_XFr��W�_�TQB�'�(��%B�TS`�kS��Y|�*���Q�z�'�-=Lb��8|�=�u^��=&��}x�h��fo�J�?�X9�O�nd��Mw��~�t���P�~돳��6�q��N�_�)��͓e��'����`��������ԡ���z�J�ug86Ba���ؑ-s��*�̌��G,+� DO���m�j�2�W�x0�%.�kd6A�C��u��*z�^0~����\���6"%�~�,ANx���'�ur��n�+�{(��"&�ȴ�������� �<��yy���ٜ9�q�n5����yZ��q#i�v.0pm���y5�'���)A�<i&���׸B����*�p����y��mt�^�����|�u9
����4�O�!�~~��!�dB|]�~��'���=BN���PV#ݎ�p�}���K ٭W+$!�d�e���K{bk<�;n�q�a&���?k@�
4�zZk�ۘ��<�|1&��y}J�aN/�jDr�W��ړ������ɧǔ:��e'[���ۇ��G�#�ɤ'�f.��T�KI>.O-{��+�M3v�SZ2sA9��������FV�ܮ��A-����m&��e�\�2kn5�ٰ�/?(?�]{�Yʦ�0��_��t`�bV��(1��Z�N� ;S�.������d�~�t����2�ϕ��N�l�kv����5�|�cB���ib���^R�F�ת��iZ7τ��V�I�I+(LD�A���Dj���f���!P�`~��@[�LU��'5�'��ɂcq5t�:
���YI1�yn�E�x�g�5��s��A���@D��V�$��K3cA7NF�1V�,r49�n;h�@!����=��������
K��oC�,
ֽ�xS��D(�pD$4HE�C~�;�ҕך��f��`��O�� |�(�TE��)rn_�d�W�7��;2Yu��G���e8:�]	�x=o�S�~$RȾxn�Y��؟�҅�g���t�0���%���|��c�i�c;ŋ��%�vH\��I��΄��`��&E���ec�+q8�'�6j���G߿��������F7�_���9��
�ͻ�L�kJsx�#i�,��6��#m�ʜj�����
a�U���ݪ�n6�3�v��w�����$�+�Э����Q�w2��<�*6˞k���� �s3��ɦzt�g$/g�{��ʏMFL~���V
�Fud\Թ�)7�X�C]��=�P��u�f�{��P���h0��\��US�Z%*c�K��,@�'�t~�������K��:���o����I�uE��9Hb���*I�>���Ύ�#s�eԅm�D@�������+��>��C���&&��STڕ���#�_��-!s��KR_Jf�VT_r�X��(�����9�.�p����`7�Ǆ��ʃv厀bVg���`��� �ը/�"�+q�߾n�2H����{-^����1���ǑﴦMVMʜ4��M�}�-�FծK��'&���!��ךR<E\��!~�8��b0�R���H������,iE��h:�j؟�ť���/_w��]�25/%��\�L=�85ْP�ժ�:q����Tkr�g�½�}�E+���J�թ
㸌봼ɢ��<�ࡀI®_�6���J�����5�O �����o�Љ��F��>Ryڧ�= m�f�D�$��������5�#��:|���,� ����2ɎjS �W� 7$n��EL��3��V�7bx:�U������~�J�jh��t����Hv��d�-����z����2XX��u��؇�8$W����Ae�n��¼`y��^I߹1� ���j�J�H�Qm�Ӕ����[��@��n��K \��������JP��lkA��АXևx�����~#K\�^_\�ɱ�J��h�m����q` �*���nd���~�	+P��t�W#�6)�
W"��&��ajA����>�+�Bf[8��Vxo�������%4�:49�ȗ�`�	bMӆ��j]���ݳ� �R����?� W�A7�3nS" L��%X�x�#9)�јz���M��̶\�_�zl����̊wu��X�/-�^��������f���_�v�(��(<���+��Q^yG2�����"�F`�=��~?+RN�1U��~��9�	.���k�̮������f?b�(��� ����L�����@�TlW�Z�6��{8�=r~o�BQ��&%�ؒj�~�: ����h�*�X���Sq���Q�Y|���L'�}خ6ns�G��uE��O����f5�,Ž��ѡ���*L�ǲ�߿���K����J��3k�}҅��V-ޗ�]/"[�h~�'��(RM큐�#��j�s��ׅND�o�c��L6���*Z9�3(
�;�����S~�n�"��Tvh.�
Ps_~"�	6pw��~Q*�P9M�ڬ�|���5N�X#��]��S_W�sg�W�T�}<�4K	��y��fI'�����/����(9f����_��i/�V�5#�*�,Ў��7��7��]3��goXG��ò�X4y�$N� �e�ܱ0������K���P��6��C�P�c�]�<N�e��s�AN�Y.Y]���84]c�ˌW�
�@�,�:��H��
L��1�9p��&*W�'�q<`x�{�H����El�o�J'��B�������u-�0�(��=����><V=��wԢk6E�z��և�<��Cj�~�����4΋$��'����	!���8˾j�Y�I��	���� �κ�K
)޶�o*U8����~����h��앶v_�(p�!����;�[6[Dj�)�����s�"�x;������Dw7�n��Ɲ���M{#�F����&N|Ra���G����U�zڂ;B���W��}�ӌv���O�`G{�>aH��hYT������'��N̆�!@&����/l�f�fKٮW���:��s:�R�ލ#k+�����o	ɒ��%���?~�������F����H|����y6{>Jo�*ͷ�޳�w��
��Z�\�wݒ�[r/{y_"ʦr6���	���G_�GB�(%WSC�;H�S\�	u�&qOk��)M����6B�z���`x��B)��l��*R��4�wN: �&{�p?'_���H-��N��Z���%����U�����qY�bF���;���O�T�d��JWF��NZ���N��"h���¢c���c��N��dJN�D�g��]����O�f�;��3 #�J7җX.�-W&�!�뤔T	���C�Jju@~�D�@��+��-���a�o�I#2W3����g3Xt���d&��Dm�zo�>GS��5
M�bU�e"+ԕY�T�G�l�;O2���/�$�ƨ" @xK�D�-(�L(L��oig��Ѷ�g�F�N�  �KI6�V��"����vd/����\��HA���-G��
܈�vrS� �Xh��޼�1�i���*�H�hշ��|��
�6�$f��@�6����J�oH�\:ED�m���OI���G	�� ��¿���\�M��ŞI�0$�T�+!)��ןjohp���|��e���qd>:��A⺾dp�e"��`N��o�FYm'�1�O�����k�-Dg�u��iF/�i�2�vzh�o�o��3k�ξ�nR������Pd�����T�1؆˾C6T1]����a���k�f����H^@k�A�#�$�<�x����S#{��7�:���=�y�i����U����Gz�6u�m4 �o#'�t�϶;Ѡ+c�F�_�=gH�9{U��A�d���kxkum�'���b�@��+1Ve���Wj#�4���x{��W[kЁ���?�:yt�pƮէ}�h��&OI�Z|m7�'�$#�:F-��E���_�`���*��=��_��[;���K���640h��WP�o�S�����Fm)�C����|�;ܛ �Da�}O��]i���Sf�8�r3�`p�ɝ�M.����A�m��`6��Z�G
�!���A�����{�".�6H��Y�@�#�1�h��7�"������Χ�LU�L���������
��� �V��G8���L�W'%<o�yip�`��L#h��V-dB���0����T ���pR�D�ᆤ]�5�L��q&oB��ɯ��p���!ik��F��b?��+j �L��;V�Q�2:}��2�GF�_�%ڬ
Z��+wz2�}��0��N�5ȱ !=닧w!u�9�W�_���(~-
N�C�ʦcj��(�M�\���?r:�0���8��*)ν^�*����ыm��^�ٶ|W�n�E���%7�'��g����ęI������b{��"L�p'Lޣ�����RL�ŕ���/x��o����3�0����"k�l��qAz��1x$_���s�z`��D����5}0��`h�"F_*J��/j����ڌ I��d�Ľng6���2uq��/����a*�%<8�>95���P��q�N�;�
\ˬ�ڥ�g�7ط>��0(;��v�����WX&����%����u��~�e���fb=��0!�leu��Ƹ�J���*\.Yfm����Y�P���/`Ͳ�;��WK�vD�!�Nh�NX�T� ��l|?(P�_5U�Jf�D:X}R���>o�����. �(��>��	�)�o�#x*���b*�K8(o��k��/�ĝ6�^y�J�-����e�PaQ�+�6�'�.����yM�f��=Rp9���.ó+�����C�ט��yM��)�䑼M>p�@@0|HK��
���S��G?omM�S��%^�\,8}#�EB�xp�'�M|��
�UR��'���`��u�@���ܺN�O2��1p� '�u���2��O�0}	���i�y�,iA1�կ�_3��Z��ؙ��wpa�&��Zm)��E�)�n�-;���_�*��&���	��?�ݙU��ϸ]�Β��� ������҄1!�I�W�?B5|q�9��%��C�Àq��?��lTTZ�v�j�xfW�T:H��-]c8��k���ZN�����ʪ�8|�u2��<��4:��6�+"剧W#�f"��3�$��8�������CcD��|y�9�a�դ�0���S�3�0�'����^�'�м%%��-IaD�f���Y���'���Nk(�[dT$�zʄ��@$�r8<����sy޴��#����vV�жcA�Y����$�����(v�r���p:� ��T��� �j]�$>�2�Q���e-�weY�3R�J�z��C8��rL�晕���˭����z@�����i-�|�������Ɂ�J'Vo'y��P��{���l�Q����*N��mI4H丸= �F7�KgjS��qL�{8��/��k�v�}kVȎ�`p4�WrX1E3V���Z�6�,�����&�K��Eg����κ�0�J�?ޱ�ٟy¼�Ꮫ?즙�l��w��ةe��sQ ��i���8[}���{Ϋra�j {���̝(�C���@6z!֊���Xg�}�0n0s�C3��D�4Hb5�Fd$D���{��R��p��XwM�B���>���O䴄����߷�Q~l�C2��3u0	�����v���}�|����%�w��@�}��Zu�g�I�v
5�u���V��\�$��o��3��eO[�L��G�a�v;&J�H������~@����oh�O�7-|�� WBw����^?���?�	}7`���cʨJ��mQ����6��f愸~c�bB���I۲n9? �&i��2�qSx�3:��K��X��pNcK,&��� f;���9a��b���"&��7�Rd�L��9��q���>Wk :=�%L��rl��B��IR�T�_��U��ݿ�'XZ&z���u�{�%�F�םF��惔{\�ܟ5T�KoNS��_�f閖5ǱA$啎ϰH���.��l� 6�V屏���n=<m~/RcE:�|<b��G�PJ|d>Ym��}(���'�9���
����K�@MT�"7�V�P�+/�Ol���>L"h5��^�t|ȶ|�ܕ�m�?��<+uY�Hj�P���;��I�pWLX���9���9�K���Hܪ����gǟ�Φ.S������(9
��U�y��Ɗ�{f����g�^�½�:C�2�z�� gT��:KL7 �;�#\���� V���f�o���_7$�x�,�s�<���
Os;6�˦./��(��rm4�g���מ��`��j�[�v���^��<��BL�`)�P�>Fp¾�p<��r���yd�<�w�Os�R��Z�*��.�6(�y�����6��_-�ߢ�*gګ�+p)�a����=���d R��R�i/AVl�ZF���t��{�uu:&#^�C _��5A',�w���������xy$�;5�N"�U
|a�^�̍>-k�$�pF�s �z�E�V %K�!=���;��ചЃ�����Q�z3CSS�W1_4�L�\⾷&�m<��C�����P�;��1����V�}J��>R�/����T�_#W?���6�j1`��Ds�:d(
%'l�#�0߆w��D^���?����S�M����#MP����>-�D��m�:Q=8 ?�J涒�B���ɐѡi���е���(O��'%�ѓ
��vQ��bPEӒ�u0�����g����(L*o׮�{,Tz��-�쨋��4q��%ގC���+MW;Hڻ��ĳ֠�|@{lFЂ:��"$������[w�;��G���c}ٱ�6�D��*V�)��,:U���=����]D�0�iZ���r�4X@�J�2c�7Nѭ\du�d1'N��z��<i�ũ\QX#��۔��T��a-���-��X��<�������f&�N�wT�IݍY�����+gׅ������㰫0��{^�~j�4�̋�t){2Y_a�l�޷�.cQ��%.Tw���H\(2�/(u�<
1R��;�H�B[��9��Ё�c�*f��C��ݏ+���i&�7B҇о�]�"~LyMb����od�
drč��;����/4&fH.���O�5v=�ꋓ����`���5h�!����>��H,��_ڏ;����_&=_����C�F�:��= Va������I�*�@��~�?�4+K)z:�O�$��l�]���,c����p��XG�f|�b� ���N��G��ɪ����ǳ	�2�Xp{ҹ$Ls#I|͆؞P˒�_�#�3�dK�Up����\"��=xv�]�Dd��M�� Ɂ�-�-���@����Y�{P�P���9�o�=�����G�,�I��el5���v݂ʬ�i�VV/SV:�������އ(s���\�W�؋&��I�
�	�,�
�k�66���V@��"�ޯ'��(����I�G{-�S`�JR�N����@w7�GtFxAB̫��YMVa�6"]b���?g'��hCE��r��3�B�����l���Л��*�۪=Vkp�ǋ`����L�Ģ��×cN�hޚ����Φӗ�86`4R�),N��q�K.ve`b\J��|)'��g`�O
�^eR��3�h�*�TL�o��|Y�q�y&ޑ��ŝ�+�����]N3eIRQ�3���>��<���F+�q�������>α�(Ӈ}@���w��n������齓�q��Y	 �i�	�?z��`0�F!\��?X���Kuu$�o,��� C�+=2��xN�z=׭�_���5JB#Z�6g�O�Zџ��,�/8�ewd���r��ϵ�Թ��Yx:B�߫���-� Sf),k��(V��A�뒵�9)�O��8�U���b����⃣I�vv竫��E&C:��Z�`��%!IvXsAw�phmy��DCk�T��Oi3������RP�G�PY���i�=^��G�e�7��C��D�,�6ܻ���Q����K�Ep��	*��n.ğ����D��U�:*�Kʆg�I�Fb�@Ҫ��5X|�h����k�q�k�4�{��p{�Pjú�_7����Ry2n
��󋿷�f��l�U�z�('�x�,p<�� �pޥG��7�t�X�2�lP������2ꣁ;�W��[���Fho��V "��cZ�:�|8��r��>����*����fU�k�2U�P�Ӯ1�JxRt�K,@�+3�!�zGw��V����K���<�'"��O�.�B�'���h�v�޷H�zJz������V�M��\�|��f�e/l�	�N���.����]���B��J(o�U�@��K�C��I���-EB�F�W�� ���D p��A�Ĳp�]ц��?�����Z��sV�W�lr�L�$��) |^:j+�0T��,����6��`>��]�oVp��;P���I�������Q�?���H~�nAE2o���l2�W����h�|sN������d7�޷�<
�`6K�shD[���\Nu�w�=<�,����S��&�s���N0�6����cŶ����y��|��/������AtX��>�A�r�"IX��Jy,�p[�&J#D�&�����n<e�����K`ό>u�㮰�=�O��4�o7��[ᑸ\��It�����aI�+����CK��ҡ&���56�ZjT�&�B�4Hq��4Jx��6e�z�����2=�N��V2�Z�P��!��R�c�?�a� 7 ����5��G�,�f)P�F�qd��C�p�1$���]�g�SEZ��*-=�sv��̈́��y�x���U�1=l��^�T�v�á�3�GvK6K��K��O')��u��}�3i�����V�ǁ�@Fx�+l��U��0����\����7J}J6�w`�⏖愞֏@�&����'4�;��Hb���XU\�"X���� �n�s5��� ��g�V����o�{p�^eS��$�͕�p`���Gy�yK�w��ve"�%C�� :���Yu���B!By���ހ�ek�;E�/��P������P
LYܻ��^�|�m��ҙ9+0�
@�����Ŗ���0d���-�Y���Wu�)���5���Ц�����C��Y�bཀྵ ʜ̤ ���N}�
�+��<9yU:�x;u��8�����m�ٮ���r�`�Z!��F����)��#��}���p�s�M莁`�6�� ����:
$�qE�'zy��^�&�det�Q���!?���<�m����I����#����Wr�Z�e�Ņ�u�����j	�h�LK�F�@ ����Jf�Bج^=�Bt���$Zf�[B����B�F6f����̽y��sY%�^�� ŭ����V�T_��v�x*�Ɍ����*����#cƢKP�U�
�gQ���j}6��}�vĝ���-!��x<�w��	�b��|�"���*�W�"�{�T=��D��(�~�m�N�>RD���Cw�3��a���5@�C�	�ۓI~��G�����O]X?�fxN�Y�s��Y��)�]7a�F%����I����b "a���3X }%l~�2�{R����&��f8m�P�8�Yw!`�rHEE��4kR��d���Fpv�x���� y��qx!�snA�_go3����n��[�.l�b�B� �XƧ*�^����~�I�]�U����u�X-�q]�̥v�T�j��2H̦���Y]��|��T���Y��M@��W�r�81?Ke���CP����y뉑?����k�yh���VJ�]�a�AИ�+��?T�$?�4����qK�R����`Ϊ���b�����gjO�u���"�h'�:��	"�>�~����"�����h	 T�qT�z�Z�C������<?����اd�q�o�0�!)~V�0����6F��Ε����P���wn��5���>�WJa�1�d7:8=��7�0��mF,��v���P�n�RźJ��ρ�#2��Jc������Z�KM8CR�5�Q��(jӮ�K���(<F_LJ�;�ws)q�c�(�>�YL��w'9�n�k�m�`{<a\y�/)
�K�J�9-x�TM�$ct���1I:yYɬm`$Ua\��KT0�[&h��B[�����9�؟���_�AO�̜�K�����}m�2����v��<��F��cن�n� ���f!�sT�R�x�_l/
%��׵,ui�6�į%���w�Ug�I����Y{;�����?�b<���rF�T��AL<$\U!TX8���8嬣	�/�ecW�Er����T��w-�R�DJ;���ۙ|���	�<����9KK��8�0I��z��7?P�S �N�V!P���Q|_��};/f�2�\��6���HKڋ�m�㩃��%�V
E�����ڲչ�y���K�-���+�S����}���x�b^|B�W29��I�|R���m��j�n;�ˆa�]Mj���u��z�ojf�.=Ƃ�U	T&�BN�ωZ���݉TyS^{dxΔ��s���hTL+�_��C��ʷ�����,��g���̩ r�i�(�n�,Q��MbZ@c4�Ws���&88�|�	�l�\��b����a�h�ܣ��H�Y�na���t���ձ:����壥�dơ����(2�`�� ��0�ڻ^��#���������	,�Hcw���ۃ�瞛z>�]E��m&v|�6���R�̋��>Fs	��":������!�B90rC�C!�"
]��?w�'���&�`FNϢ�ɡA��u���5m\m�D�EЯ�Fa�j,������V,�q#m��&>t��R �n�z�xs�cxTC�C*���_Ʌ��3}�lP(���S:R�'�`ǌ���P��5X���(Iե�: p��s0A�j�f�pP�3MX�-�q�M��AFb4�)��
Ȼ��֎Sf������!b�llŶc��W�jR>-}elD/�P!
BZ��*E(w(ѷ��f����2�W��r�qoT�"�!_���[\�9F�>2��}�~*��K��/����[���3���xA�f�b���ۊ�k�ۺo|��B��8�قĲ�Z��3Q����(S�r��3 ���e�c;��� wb�h�1ؾb�z�8��.&�/Ȍ��џ�w��L�{_f�3.OD��O{@q�ˤ���l�[@8 ,�ה�����#<��%���!�K���B��ʑ�����@�-���'`oal|.&�/��؟G��a�K�汘��S���!�M�a���G���p���3�iM
����>B�j&i�р�B�W8��_���JD��A�>7Y�\99K�7�F.[N [}T.$8���<���&u����y@�d^�F5�"�K��8� �2��y�s�ɷE�	�y�)N�yr�j����u �4)&;��+[�+L�e%�5�̍��4�k�}q�L2���U������Vp��3��^Ŋ��c�3�.t��TW�;Y3�)|����$V��N�y]]����9�4�fKf����t����wQ^H&-��3:�����k�p�Dt�Ji���cB��b��<��ƅs�o~�.��Z�r^���vY�+z@u�	]SDl�eI��a38ET(֝"2�0D��×al���ZD��Z��=P�����O����-wM]��	��~
n.|~Ao�n�<Y��D�A���%�AM9�V��N�a���O�E$Y���\� ęU*����!����D�Z�� |Ȗ�����r��z����g����q�0 ��fd�6Q���.�W $Vx(}`Z�o��tC-|�=t
��[5���ܐq7�/ �mM)
4z��@�{$���mS-f��>�v�@��"q���Q��}��=��i����
��驼����l�3�&[�LL���]"�+[����^�v��`����?/���$�bk��x8�O�aP�9F| y�gZ�B�q8��9����A��K�DOJ�P)drz���+ub���&�~s�_gy׀�w��+��D֛�aSZ��:�T�� [�ʂ�E�y�
��Bp/�|�]r�~�����2����9�� $��W*��>1qɋ{��o�R?��m��X�i';�B�ݬ��A|��b�,��gg�O]dR�OC�����2tҦn.�f\�t\O�5��us��%Y��Q�H�{1�Xm5J/fn;x��Z���j�w@�� ��^Ip{5ƀ%, �C���8��9�c4R�T��}l� P@p9O�JE��n���yJ�%�f�Տ���
��,\�}����2J�W��V+�9u����J�њ9.�h�	�1�E�����6��!Ȁ��t��V��X���R�=��Ʋ�Y#�p]qޝ�-�M1!h�Ϩ*��w�r�b�Xw˔��',B鬸N�R��2��H���J����aN��Y�ѡJ�n�̷���]���	��\��R�/�T�
�]�_
��(W4��e�d|���t�|����b���V�ɶ^�e��.U"��Vf缭��M�V$���W�[0��}���S�T�2eW���S�'`��m6���4`��R���F�S���P6��r������"��`\oMH8�A��q�`A
A�� C���uRO��vn"�Z�1�R�E�%�.��:o�O������5j�Т�A�W%`��-��#�˚���>}���o�F�l�PB���C&�l�H������B$2�rxA����[,��^�(U�e��T4���n��C��R�7:uδ@���:�N|��D`�u�ۖ`]�;��f�`���l�J�	R�d�ʩXP'�BH���Ʉ����޾��,�vļ���+�3��N�� �~X��M|Z�-����|�A��Z"tq�&�Бerqcɇ�"��*�H�t($Un)1�<yO�[¦�PYGU���7kM��q�� �sA�Od"F��N��E���;����%���$��&�=o.��L�'�<���&�����[2�8��N*Y1.�j"V��`��J�&p�E#����;���y���0�>�̥-�7PD9��l�;t@�����²M|:�C��F�rB"~K%�<�������8A�#Q[0&-]/
ry��'e^A<���B��,�L>6ce8j�.l`�y�ET�y��/��K�*��GU`�9n�Q�_��@W��w\�'�I�� &�Q����-*տ����J�rf�o��%��%��h�j��̞H	�I��0A���Dw��Db;M�ig�fӫ���4�;����^$��Z'�%�W\�:�3怍d��M�at���[���g���H��I%vgE��k��|T�h|�A��'��F(�a^�X�f�vZO-�� �j �賦���մ�C~����PI����H�88��YL�����5	�6uL�tmC�il�/B���|u.�{%1�(!����Fѓl��P"�=�����U��q*�l��j_+��s��+ܦ�����.CU�X2�V�>x�w���sEG�GMO���n�A�N��k�r�"< �l x��~뗞]i���3lc���������z��V���Y/@�NP���;꣖�� )�i�i=�go�!h�(O�x�O�|;����x��`��Ŋ ��H�����z�uY���������ֱ��%No�̜N-�Š�c-�u�5A�A��>����;���� +�dWA�P��2j9��rZ\]�������I|l���q{�U�_���g�-�s������v��3v\1r@�H!��{N3����DY�Y{	g	ιt��P\�	�Ca�\>
8���a2�9�1�'b�Du����~p��I6�ٞ���;��E?Gi�U���4:eim��)sí�n�~%�%��>pۉ��ϱ�`l��B��Dn��=���Z.&�C��y� �vt�xX�E�Ov��BJM�N3ͤ���n�*b:�bh��Ԯ\��!ƅ�{ְ��-Z���������>���2�}tF2!$�-���;aⓞ��y�Gݚ@��O�Tumq|�s�ֆ���突���͕#����Ȑ�r�DHZ�?�@$�)����zs�*�˄̮��3�;vu�+�3�l!�7��8�f2�	PҖF�L&��ő����������1V��i��C�G�)Nt�_�8X�ם��g�|�@����kIC�}��W���#~�U�:�9	[��-���� �{�`h����=s#,�9��;�?qW�N˄z�&����fR`vw�Z&��/'�LAQ�]����򿤠������Hh��$��β��J�CV\�i��]ìl^Ti���15U`E{�]�	d��O����Ew��W��?��z�����A��-x�Mp�?�$���)���!�E�^E���h�f�=��C�2�;.Ou_l�uo�68/4��ʾ԰_��C����+%'��'�ۓ|~���j�Q�0g�h�?F-+G)s�I��Ѐ�P�l���p}|�"���a�[V�ww%�C�G7	3��ĵ�nx��������"�Q��2��<&�`���	�ئE�~ݻ��եS�+�����V�\!v*���@��ɫ�}��I��ш����l]�9��QB�ބw��U�]�$��FD�]@��L ��ν����I��y<EZ�LLW�	�gR�R�Q�(�]2��+���3C��x�ի����JՄ�X����#=c"�S8^-C��I|uP�B��`7�6 �7�#92���~�4�O���Oc����(��s��Td8y%4C�r�p��������b?�F���y ~u��9-�Z*�#��S���F��,������q+H �?���a�0>�3�mh%���ur=�]n'N������ȴ�����\\@p&h	d&^�����6W��/xZJkBr���ѥ���wMo!9�F�<�C����[�6�ٍ�\�KH�Zdy9%BXp9c��@�r��?��{cɿ*w�{g��<=���~;7�ꈋ��_�|h^�ڃ�Hx*�h#&m��ڲ>���&���ˀ��ꘔ��~�\3w�򑾄�`�c��Y"M�$VT�б�� ��Ra���!�_ǿ
�f���eV.�rbG�j��m�P��ax̍���1�Ǖ��]���%�Qܱ��>?�)c��0~��G��!l��TH��0���ǋ1j��I���p:/#�dd��#x�Bn�L�,X�Ny6A�̆
�ڕIz������xϰ��!�ߕ����r!W}6}�N�}[���3@b�;�}E"�����R7$��]��N�Qy��2	f�Ľ�� �e�� �}�́}��(M7<��9u��X@J�H # 8'����q�R�0N{䄷�U��Xm�����������*�}�a��]�f2e���`Z*��)��� �����͞����3��39�4�i���1IsqG�h)h�R�>q��3��(��-Zڂe(��2lu]9":5�����r�z�X̲BYj
~�x��]��q<Ć���(�d��dt��ɒE��^�Y<�v'�WV_�F�HP�nr��~��1�&�݆4�p ����\D`�����H3�e,�X�lUcWyh�ѩ���s��2�u�Z�G��1F>�d��g]�����c��v���8f��i�h�-�V|;�v��R���͍Tn��ӧh���/]Y�� ��d���z)�[�IF��D�Or�oa�Cb-ݺ�������i~� �\~AΛ�ny/���Þ�|��6�e���Fŝ��룲���>��7~�V�v@�y�_L��u�'�ll��dҖ>�\��G9�ƊZ�^�3��AP��zç���i�O��ڢL9��P�ƙ1�{����X��w�T��Ik�%�I��ܛ���{	��*�&Q���|@V�D�s��r^/������@�)�{#cgFN=o�f���x^�f�!
�)}z^�	(e5�^��x�#�e8�dwR'2���I@��³��pxOQO�A
+�7�h��~��}YyX:9�/B.����d1[M����Q]���.?��Fބu԰\�7H=�=�WQ�:�qp<6�NAݡv�9�)�쒑���]b�+�G�)�eC��5?��6��^H�n��P�w�JD嘉Lx^�Lu��V8�a��u�-�ߖCZPm��ø�M���)wV}�{sf	MJnBu��t㖈��g���T��u��w�|$o:#��c��6����T/���J ��������6�Pf_�}}c�O����t��qV�=�0꣎�r�S���N�x�^���P��W㿥/��y��Z�bI9�Z���E9��H5�����-��X��	icvD�rO�|�����P��.�K�����J���������L�?7â�)�%!�?�֪�i=Nu�B��4�m�!��6R�%E-S`�a����V�����������&�����M�b�J=���|a./�ƘX�;m�����-�?���.A;�����`�R�����o/<L���WW����HE���Мo����ڟsVr��F>Dv��d�Ū� �f��T���,ݍ���NJA��,�������|)�7QU���]ԉ�>���u�G)��W�z=3;�G��$�F̟}��T;�V/�5���6���xOj���od	U�a�����kd߶�j�)��)1���D��ߨ�¦���,�'S��q�Qhԥyl�r�VE>�
���'$M#�-c(���Zb s�`y���' <����W�.�������Y�@Mn�(��K�I��-"\�r���Z�@;~�ȵ�QX�Z�8���(Bʐ�U����4��Sb������=X���9I�l��+�y�f����)䝯�e��N�fﬔ�XVԉ,_z~�l�K�p���뺙�U�?�h�э;\8$Pk?��������L��E����XNH�-�x �kA�!r��o�7� �#��$!��lun����j�$���]h �щ���G�x�}{��M�z'Fy��ۈNO�S"zKz,��`�����P�K�+`?ʟ讥Z�b@��_H�Lo0�P�%���@�P%<�N\�{~׈��.t{J�h]y�XwC�6��q�4q�Q%�����(S ���������#��&a�a��i�[�>w >C0�dy��@��g"z�6�:�c��`��p%b��L�?G/��Ub��؋���e��f��>��YbR~��c	�L�i��<KяrW5�mS�nv��gP��l~����q�I�g1�yH�{��h�0ރ;kB����F�bB˅�`f�Ni|����l^(0%H��C��T��<��/��z�8ǐ���r|�����w�w��<��/��x�r#g5p������b)G��x�A��?�{�y�:����LGw%MV�䚯w��H��Ta���1
��9�C�U��-��d��rw�N� �!\�ˮ_���ڝ��\�T�3�[�����=�GH�kXA؝֞�����yi��]��>}�f��W�'�"ݚ��K����%ȇN����K��Cl�,�e�f��� �/���Q��|�T�x��[Fzf؛3!ײL�(�Vk�wrUntN�ő�G�S �1�u��^��2�u��o��(i�� B�� �tIyٔo��3Z�m�Ѽ�����>TR>C:�x	c��;��݀����G��x�$��9�m����Y1���=~��d�J��9p��?�A�}F �Z�C������2�4�*d��<��b��F�a"�~v�9����BT�+Qל�x�tgLw'��=�F�u�{��y�+�h�җ��<B_1�:����FG�����&zJ����0%�C�v���ϐ�E�Ѫ�`f5�5 �AH�,�%��)�@���˶;�y����!%�M�[�1W��U�΅�����t	p���E0I`,�}��m��t[`]�l�+6�-	���h�����{�ϧ:�������`������#�%p�z	��<}�*@��Ȱ>Ue}��k[�I���5��9����ǽ�W��w��[eC��f�&����~�#��M}~L?�_�b�Jo��歜�Ь����İt����t�,R���*b*.G$֪I&��n�eO�S)�˴��$ ��ɎV���xmMM�o�����ExR� ��lw��T�ω�nj)d�A8������|a�T��ǫh.�����'E��PTc�{J+����*ZW�l��K���H��,�h�]+�Z���P�{�Qj5؂�B�!0���Գ�4Ci|���P����._��v�CǕ�c�JXx��k��aΚ�bCh%�ͣK��[����(7/ ��S�V�a@�A>I�ц�^��Q�6&-�����^����ᘣ�R��'����9�6����g�D�)�^�Y��s�u�'s�A�ݳ�ua)��7H~D5e$��ó���4&�HE̦I�]���ۻa��q��9/����>���(�O�Ňz����vPI���p"��c��a�v9�j�_�ﹾh�k���r6��������jָ=Y��C��� �x�9KNօ��<W�#�O<�^��o"'M��������w����B���'IrdR�ycCдJ��޺����E�}j@2l�#�S�s���ox�3n�d7M!0w�$jv� A�1����<d!���k �XN~�G���C���(I@�߲֝�;q�0)c�!�0a�%"2���2�%\fe[�|�E�����hh?
����` D%c�i4!�Ƚ�In�pN��LI�}�C3<�X�Bt۽Z]���c<{����������{8�4���kuϾ�nn�� w.cx���`�����`��JE����6�]�<&K�fl�����6���M�C�B��u�8�r�E)��4�0Ⱥ��W����D���9"W����;`z���8]�=U���Q�W}�Dk�~ɳ�_n�rp����ON�u��L�u�ף3�i���Ba��#�Ӂ<��a���Jr���4�dIJ"k��@��an��<.��u)��W���ES�0�s�z�rn��c���~"�d�t�X,uF?��Y������MCN,�`�u��]J�y.ސ� �Dc�v�T�v�J�pƟ"s��<9M�Nt��,v��;s��Cf��GQ��q�&dv<��p��n��Ó�z���^,�Z �U�v��1\nه @�ǛCޚ-�oꐇ�9������1B��{N��O$n��؅i-�����1T���<B�#�d6A�����*.�֯���7.RGl��q��e�Զ7+��|ڏ����̸�?ߤ��V_&���!�a�B���O$	 \F�`�F�'�B���C�޷a�Y`2C�Og2X�^��'.@O0.	��������_*9�n��a��à�k;�	OsI�v��ϥ��<o��`�zV�u�v��g]�bE�U��1�Mb(��>`Xjź��l�� �7�����겓�d����`77��s�>rboC�U�1����X{�1��o��9�vg��]K �1�s^<-�b�����~�l� /�?��Fw���`��H��>�0n��8�n��������������.K�귳���N���C��������Y�_���Š���!�o�i��~fo�@�8�뻇O����"4��׈�;Ջ/�m�Be7B����~^��B��S����v��ꎩϜ��j��p�)i�$��W"����*?�T"gp�`D��:F�զF��7�x@�3�B>Ga.� Ř�����f�L��$ ��[�>:rq���򝮇�Z�p,B�)p�#�=�!'!p��ԁ̙t|� ��h���D�S�������|��d��9Uf��C��r"�9-[�-�Qj��B�zJ���8���?A�)3��V��b"�0�{L)Pnl�ӊ��ɸ��C�S�޳L�s�ҭ��������U(���t�.z�ۼ��)�z�$ޣ*û�_Ėm�ӫ��ĺ���H�s7n7�D��z�qS^�L���&�k(?z�� )�%�'�}�����k_;��8�/鮾��F��O�����e���۞ϐ|�ZLI\R��In�J����U�	�]6��#}�7�j�^r�|�*v|7�{e�'vV�z5h>���^�}&L
��:�����R���>�z�@�^c0�J���r��;��?�JQ�Nl��T��Cf�T��n�~�/�}vYXʡV�&+�b)$^_��aX|��G"X��� ��t��"��>��=����tE���Xb���P�i�V���;�߶Sӆ���J�ڱ�a������e�����	�=�h>t�J�֙dA�l�fĻ�ɷG�N,��s4l�9��'A�Ǭ��PF,�����Ju~E/飡{eb�'	��,��y���ڐE^/���_����h9�_����w��*�&z1�A_ w{4V��l���=A
�X8Nv��A"ݔ!�vf��F��ޡiB��>9�����Y
��3�h����F���;�=���d�f�����ET���Lm
ú)��Lg>D�$�o2��Z��S�{q��5����	#]tS,B�����3	�UCL�.�������nf�"��n��ZLK"�
���S�H����I�Ή�6>G�w��{R
�Ϯ�j7kn��g�z�AI��7c��������,$��"��/Z)3�2|y�pv)6Kk@�����@�}sI'}�9�|�d�� �@�0�U4�1$Rs�r��/��nI9h�-�>��;��f�'0�ib����I�?eZ5K��UINS�G��l�M�B�ʸ*Lk��P�{�s�1߯��iq��qƼ�1��p�ŏm)��W �ѣ�dO�z*}�B6�gr����F� ��bH�|�`�^nv�Ѡ5}G�(mO��x�� e��:�8�H[ӝ��1C�#R��?.wU@_��6�0�i��O�#��I��֩�_�	���cgߚ�}B8f�J˙�ڟ���gi�t^�4I�-������v:�����If��u��5M8z�ղ�\�Y�������٤��F�M��U.�2��x��?�4�xw�Y��aP� �g�`Iȹ�q
�y0}�2P��P�X���|�r�z��������W�a�Ig�H��� t�Oʋ�0�[�l��^�9 ��9?n�����	�ϒ��DO��������́�Ĥ�P�{�x=5J�̔QC��sr&$V����D��a	Kz���V6H��e�T�6|#qGVU��e4i�"uH-� O-ڡ�+Z�(t�;^z�7�vܓ����l��!��֎��KF4;�3g�(y�[rn_)�4V��X0KE���� %2C/���	2(X��/���Ci:�8�O�so$��ړ��k5�b���7�����r⦟���ٖ�ƤD~R�Y-"fP��U�y':*�F-E^������aWo�
~���*zx퀶'�c����5e/$�<����h!6
Z��+Q�������I
f�I��&Ng��#[�;=o����I|�h��'�T�Ǜ��	V�'��٫�em
!P�rH`t PF������7Z���2@�g�EVQ����
�;4C��0Z��{�?�8.��Z�����Kp�7�Xf˘C��^� ʐ�o�&:VW�#��u�G��p�y� �԰�6b��*���w�J�[���po�/^V��]�W�xK�*u��y)�BCI��U���5�9�`���`B'��*�DU2u�خ�L��M��JJ#8L h,����0�搲4����?͈M �<Kq/76P�i��\�G��2�h�6n�@��-b�a6c�(���"'�������B��9mA�ah�fh�&/5��@����R�M�L��^��m��܁H�j5���d�$�A��<I�T��ш�T[pv[���_���U2���!J����yq�辕~�>��:�F� ��:�2�v�;5[Ĵ��N�����Y� ��S8>��~�d��D̂,/>�/+�}�Ul�� K!�$�) ����Z4�k��Aw/���$Iϻ�����o�j���J���Y�|���u���[��leq�(�3*�Ve�̿aVV�hZ���}�[5��\=)|4��e(mN%�џ����|�u��zެj	m3[QtE`W�[����V��c��A�փ-�Q��`Cn����J��.�[\YO�#��I�,6x0E�#��	:x�}��S�HH��g���U�����R�g�r˗ߋ���'�\�K�5س��w�Ɛ 7(>"��w� Rм�n�=��q
Yw]�e+4���q1;s�_p�,З\��eޢ��=;ō��$�FB���/�tET��p�W��'Z������f�\�h��v��W��8x��7��]2blE�苩C��C�C�#�b�J��� �~��s�a�'[?�7P�#�zT.��^���։�;��5�����
(����y`�����_�k�
R2���{��AМ#ǰ�Ԅض�!9b��qXˢb-�!᤽9QqRE3��pB]�Mr-��+#o��(�+r6��*��rěv��ốsn��@*�d�íD�r�^.��>�Z��k"��v���si?�Q�Y_{#=�QV�º��ٽ �T�y���d҆H�S��B�'�K�:yۢp�(�E+�D��)�����W[a�8��[����	�&���y�'��-��e�fsf\귣=������Q:{�3]�Ś�Z`�Y��z=1$Y��|K�fM�(
���-L<NwVa}�:Ӥu!�L:��Ey��3p%���t��̭��<�jh�%�Uč�������}�o4V����kj, �7��$s�pth��x`:%��`_"�<b�z}�u��/඼ }^������ɱW¦1���>7	#t�$�~��y�z����m	2<ۇ3_����ע��ԙ�]%�i�� �MNx�d8LZC2���f�ܳM��I`��f[ʿi�`$�Z�>�ʦ6���g�s�y�cb��:�R�2n2G �g�@X��`J�E�g��R�����L�V�9���X�#z�����3H��n��Jm�$~�i�6�{���B+$-:�N]+m�\퐿��s\�)ӹӇ���傥�A��!�zf� șx��.?�/��v��
�+Q�m����63cs/���������1qb{���m���'�r��}DD��N�r�Ǿ�s���qbcǾk��y�C����:(�?B|��t�,\7�+��Az��Neiq��։�:m��;z����%��WG�D��8`���͗ȃWӪ��|b��A�F�t$_�'b���q�1�|�����los.�QO���fM�R�/%�9�gU�.4�HKE+$�㟩�+�H7\w����H����9�w��l�Y�NϚ�U&q����V��!2���&�S�i+��(N#C�l��f�}(�4�sp�@�B0 �I����F�S�$�^�"�s��h�'m�L��~�{���}2�Ϸ�lµER��0�D�Gϸ�&���J+ϊ�?��H�vL�)Y�8�h�M�V<!Ae3۩NV���dxp��y
���~xڀWn�ͭ�G���ǯ�U�?���1��mMu`T��=Y�@��k�x�ytI�ؽl|	i��	��G3,���vS[�ڴ"Y�X�40r}�Z�p?�U�����N�]�J���������E������]5����; �
�}�>[$�٥8n��0�:��'���n��%�:Γ'
��ڝ.rx�_6GL����aV|#O�z���~Ms2��RR��K�r�|�Y�
�8�z��Q�.g�S��f����돷��( (%�Yˆ_�#[���֞��s������II7Jt�~nj�u�3!F�X�Ps�ێ��8��Xg/S���z����1Q3��cgޞR�{���lhx�c��I�q
�|���4�)�z�#;1҂g�(�L�Q�eB��Ы���v�=�;���[���X�A����u��W~��cgc���B�@ �Œ����ܢ�w���caz��ǂ>S�����Y�Қ�T����#D�#�� ��Xyz2�9��'9�O->��ߛf�<6�j�4�+-��A�kX�Ҁ���+�Zw3���i��*��Ф���K�]���o�)��aj>ZwԌP}��W"lJ�Az	����HEV5�SoO�,z���pa�w�V�Eb�^L㷓�2KACX=���R�</F�]�����A���H\j.�����_�a�-LE�O��g������||h5� �o�7��Z]���q��X��9���];[m+17�¹�#�#���aO�x�]��N.�h3!R�Ҩ4e3���	Ƀ$K�,[�a'��Pas�9uYt���̔'�є�I�2oM�:+�Mb��|gS�O�h�A��74���ݬEfiXfD?��Պ���5���jO��\,-�6|`8R&���9=󾞒��r�!������)�}Ua��0WZ�ׄ1A"=��:��YF�=*S�k���ln��G'���OJ�03��@D.,����9�
��}�����T���0&}�@ �w��7�D���ݖ�>���o�[�ގ�o&j������L?�:a�ce�HF���0~�A���'������n��6���c��M,�]��__`���^�4��O*?���K����hmة&� �������VP�m�����'-�5���e!l�]��۪ K.�塃�eq�s�Nv���;vYK��*ǈ��l�KX�7O��*��C��2�{����֟J� ����ۦ�R�C��V��J߉���zu�z�� ,�?���q��:v뺙'���
M/����^��?����-��Z��&�s�����������>���N��%I��݋Ȉ��Xn��۩9cd6�i)��s7A� ��8q��M��OD�Y�$�g��v��M o�5U�+�Vh��$�t[���;�JQ�>��L��l��rp�a����x����,��$Ԑ��!]��S5�aA螒ki�!��f�}~��M�}C�o�UM�H�<:[6��p��{3ٽŁ9b^21�殱ظ�O�%0T?�*��h(������,M5KϳC�=b'�61��sYK�L����f�1T$pP��%(<iwL7@�'w�Vp D�o$\��Ϲ�G�<�����_a�g�۴�h�._%��j�K�e`琺ʀ5_ďc���81]
���)V�'m�p��t�W��q�VD��E <fU�fj�t��*ʵ���V��k�]Ѣ>W���}i�
`��_Ds R�V����a��}o��	{ ���Ί^U�M���+��ރ�h�`ӓ5�؋iEY��b��ճ֒�߾�3��m�3�,yww����!�����5��މ���xm"�xj��5��W��-�UǦ�=��'�M���;�y~ݔ&�{wf����	>��E�����S��2�<FlL����+N�s�~Yi��vq��Gz�w!�i�$��W�fw�s��I�37p=�6���ѻ2���yk&�J�f[�>�e/fT���H��Ry��������X �kO������� �4���X�B����0�K�}ƽ[���<����a!.3��i�Lhj��K�SEd���h��Vʩ�n�Q�K�rQ0i��3_S����-|�	[9��8�.-��6��4���'5\���h]"��� 尤��x�4�o�,�%cy��ٓ����O�$v��a�x�)e�-؜1g�kD�I�f"o܅��o4��z<P\3�D���m:�/	�4F�]c�,	,�����ܼj���n�iz磅l��������H��TVr$��?�<8n![�زn��SZH�\���!��F���J� _x%ĕ�56��"��m2���f���ځ�mb"�{ۈwP�_�&���M:V�;�^vc��D���D�������u7�,6�'�^ռ�T���=�����������Ph��@��s�6��o���.-�X�k���	����J4}/��̯(��`&rڋF�z՘=]�"{=9��v�C0����C|���p��.l��?x�,�}U�q��;r�qڵD��BOh�ۗYV��!���N;Fϲ����E�k.�$�QVE�S$���<�X:�����&D7�8����0����l�gU��J�ֱav���cO^Sn�� F0���bĢ�ދ-T<���ݕ���YF�|�'A;L�^�~V$�)��.���p	�����l@��D�}�w���>D�����,e�|�W2�M�^�'2�G��R��2ߛ�}k���}���x{yd�M������<N�
���o�$FU��]����L�l�' D�+���)+���<��Yx��w�g���<x�f7��>�'�V ""a*U�{Y�V��s͕[)��r_�|��`�6 �M%��č#���h���f?����`�HD��0m���e�+�(��j��%��xK��d�'��ޛ0�tS��>��-9�4�|�����#����v�g�I�8��r1ڲ5��I3q��1J���i��z�C��,����F�r͉;x��fڈm�&Z'�5�6�m���c��~E5C(�|��F�������������a��\���}&��7����H��Jk<�*�H~
pZ�x����7#�fA�V� �>��`�R��H����/��'" �:�R.H#8(}� g����v&ԗt2�J�<�2-�r�~�
.�Źq��8a��Rb2g=ƞv�e�	ń�_�J9��}s@B,�(%}���Y
�~k�ӹ�����7,-�w��R>'�L)��}�a)�c�	`�8���L����ɰaR|蔴��v0E�Rs����L.Qc����&�R4?xz��}r�m;Jib��{+�����q�3��S(�����MJv��K�)+�2#�C.�����2�m��SL�歴n?�#�9y�9���g���vU�K#�;@D�< xR���H�t�ڋu������ѭ/@�ڕ�����h�?��,4GA�]-�+�zR�ٟ��w��oK�nW��n��]P�Q��������D��}g�ڗa���Vx�e��3D� �$C.�@I����/��x_��s��d��k>����ƻ�&Q�i�d��"�E����<�,��~(K�*6cQ�a���]=��I�Fd���ҭ��1�J���_j����-/P��f�^��s�L�ލE�/��I��{SL��U������Yb˒�~�uR��K&���ʁ�t�/C�Y�A�œ�����j��;�5�ӽ��k�f�j_���}�v'�P�*��ej�˺	�����졸è���<`��[���C�t�`��Fo��K1N.F�[��A;x��c&��
��e�����X3�N�s������E�p�j�}x��s�M�%.e�ͭ����OD���Ё�U�
#[$�w�:9�`��� �j;�����?�P<k)�T7c����{R��f��$ǧ�(fV#��k%�r��ס��Ӕ��(N�t�d0��}��H�҆?0\�"��t��z�KiD�ƃI0P����B�O�(�M��^
�B�O�~�ޖ��3P�����U���z0�T/,��*t��h��1�4��s���)���O��S�7:�L�E�E[�D��F���I��/�މD�x\	�]5v{Aƛ� ��c�CK�+��_�jS����A�~�\'4]�|��O��<�R<�H�}�S+]�{S6��x��5��/L͈��٫h�u�ꐵ�4)�h<�-�ot��m�b�5Ŋ��Arg��9�Z�΁I~A���2n͋���iG
�DK_��&�D��
��:]R�s����1�?�i�Rt[>��!�~�rс�����G�-�k)GvL�΂y�G.���x���e�T�����RF�$�7�������:#��Ȅ�I�L���[L�y�N [P3;Y�v坦��J�m <�L*��ˣ�[�uJ{�@�9�|Q�6�F�~ 0�X��X|�y�P�\���_j�AxlO�r\7�Z(�d�&�\�/��?�-����/����X�������Vj����	�bLZv�y�5|�C'W�;��uE*A�Eөw[�0B&�f��J�S�zsMO��'wM�#��� �JH�",�p*z���RGpK͡�X4�U�P�UQ�S�f�pB>U�������%�Ą�u�fS�"�&d�t��x������.!.3G�����9g�n'�b�U;G�q1���d�-S D꧛C�������dwQ�^u\n�re�"B�b<�
lUk
�! ��.�KVr����I/�~��4B��;Ѷ�Uiȱ�]��/������Cffd�g <��L�OҊaR��J�y���
�������u�EWO����b���ˤ��N^�?,#e��Se
pp
v�`�t�vo�cWċP�<Tek}@��~��� �T?���C�镠���d� 
o�4Wa+��iqB�"����eo	�/�sN-��G.��M�@dQp���,3����`��]�5r%�'�eh�$^ ���D)��o�d�s�L�@���6ﱂ4 �U>e�p��G���- �Κʘ)4��v ��_��������/Βr��#���)��lƑ�e���A��j��7�o�$l<+�p�����x��`t�ϥg'�ӿ���X�d�F��M1��y9�����x���x������a\ITif5y���ȻN����&T�4�l���U�.�
���`��0�Ĵ�?��?oq嗟��\d��o�[�Z��5tQ|a`t�U����w���8�&؜I�g�T� g �6�]WЃY8�vhK|���&o�F�	�������D�Dc�4��0�$l�r������]���������6K���ۄ��a��)���<5������yolk�q��m��I� D��w�3�u$F�d�q+���i�S�[�,���8����~r����/��	9�W�G�-0���餀��X�q��;[ Om�f�VI���저v��X>@�;��u��} <��{�	����']ԫ:���5����F�PdU����Pk��A@D��7̲�Ԧ��t���[2F�f3�OL��X����S	g�$�T��	$�
�lOS��*�x�/�^0�O��*��(}��JXU��丽28�	�����Jl?��Bb��D1�|<R��t`��P6�f�:���.�I�����"�ز�8BC�?��iG�z&��w����/�Ql���P����ũjo~/��B�-s��g�ju8μ1����>�(�{r��L���ݽ�9\��xi��R��e��9��,�F��=��O&kwU$�����	��5Nt���e���������������U�k�E��Rr��	�3��&��^)Z-C�a?$�3���T�geU�gǩL����\�3��Ծ7n$<an�m��!S�����Et�M1$��=�t�$��)N��o�4�D��(A����`3���s��&�fJhF��OI�B�&��8��k�Lb�]v�Mz�HJ��b��GK(����ݐ���H���w��󷸶ENq1�� ����Qu_�FJ��;6��w��o����M/`���݀DI��)�����1�1n��f�����>V�C�a��u�Jt��������w�e���m�`$&6�	���SP��F�`����W��t�Y��-�q=I^V[��������n�ڐJ=N�A���4	���8��
Yڳ�0��\\w�H��j7�)'B��˴f��r��/,�DXʴ�Q�ꎡ�l}J��#e�Z�f����]u� �=�o�������;�+g-����0j��c��B��t�r�o��3���#��1��!��+65�}�|��s�pQ��TQ[���3f�*6{���r;"�1�^�;�R\9'���:��i;R`�=\p|��H��a��^J[z1j)�t��&�� Yz�k<C�¡?		03~v
�izC���M��\�v�h��:�
ᗫ��� [���{Nn�KsqQ�-!a[��R�E�]��?��w�������orx�.̧c'����6�A��&S%Ki��_�3$���J��)H*�|�1B� ��>�n+ejPF��a"76����/��������#^:�[�{�
x�k�"tdϨZ��<`6V	�(���1w��w�zS��Q��8�^m���UA!�V���5Z㉭�ti����X���;�Z�(#4*���h[�z��/I�C��ED���*k҂�1t�{TX�R���j�2����=֎�c7��5&-H]�f
Q�e����$�B�����#�|^�p�4U5.��aOc�c��v	a�֧n�G���X�3��]ΐc�-�0{��{�����g�ӹ�%cRA}T$�DI
T��I���QJ��7�����E#@������T�n��D-Y��K�0_'�2¸��Q�+&%�q)�����⺌K.v�,�^�d#��?� ��T��݆�&S#Qv{�<�l��|jB����^��ԕs���M�Ou�p$�B3�=F�ۣ�$Q;�7����u���5��5W�3@�$&E����,lx�+�=�)5eI&�q��?�IE��� N���*���٭&����%g2�"��ܺ ��P>�gNp�5HƋ٘K;��������P;�+�C'���Ӝ"���y�F��	ڣ�����1���
���ӂ��T	����f����o�����O(���I��\����
6��l'��5���L�[�����lc�lW�,��Kąj�qIC��� R����	5$l>�|�8H���1r9��_��!.%�AOpusKֿ	�G	�d�A
��>�p��� L��lY��F�x�4d��-�!�c aC�}���o{.f]9[-k�J#䜺4��Df���x�A��q�i����	�ߚ|i�kfɹ0�BE�n/�ơvlz�%Q�W�LѪ��E5XTF�������n�R�\��c������\�s.�ReU���C>��w�W�!��O~	�Q1�`)���h0hJ��0��Sp`��ꋍ&���$s�n��g�<j��-�Nj��e❗8�����#	�?�M��7��eH��}|�cL�f�P����SC�U����$��Ѯ�2�5�M7�1�So�$�^q�:Ǭ?�~b��"nW�z�:�o@^�9�����0S*��Ҟ�8qy�D2s�y8-�����p��O�Þd����Y�ʨ��_�y�'�v��F��~��{ul��
U]��B�5����q�K2ؘ��E~�������,�%�k�ڜ�]���}uf݈��!������8x�H�R�-[������7ŕ��3I��*An����P$�q*��0H36�:����%�b��%<�?�G`�чY�m�5{_�JY��� ���Hu��x����!��\R��91v�R��')8#t1d-�$.̘Z��~�T=�k�s3�ep�iL����v�!l$�c�؝�a�MNS�/����^������6��tء$E/:#���j�ٚ����1�	�x<D�Dm�m˃pq1H<����x��n=�̍��0����dE�Y(�!���*<9(��S:��^�[�Ksu�2,�E��_KH���A��&�cX3�I�M5�=$Eb�<�����Q,�fwr�Q@W��n?
> 7v��N�W��=���ł�"�w�a�?}>�l�/Ks5B����<��ۢ �Į0\lv����#b�R�H�K&B_}$�	�����'e�㼆11gk�|�m�7s�x=+X�T#�e*����;���||�$���t,����l�X�_�N�~��x�&�Yb`4������5�'�_H��$v�|[rR�+�~�E	Aɲz���+�����w�Z��e��-�Qe�'��Te`Oe'�yu�����0�ɧH2ىf�d���1n�!9�,�i����h̍y:�tJ���EǇ��OΉ��#��2F��u҃�Ƌ�y3g ���<�t#��e���#B����Lį�����o:4(Jh- a��ʝJӀVR�zQ���%�>|zK��'�Q}���r�᭳�"�;�_��{�9���Tt�����+ ��<����1?"dR��dɁ�~(��ԯ��.�ڐ��@���`�>��F�o���j � W�]ė�2k���E��!��$��#xu�[�X�6M���X���<�9Ks��4�����7�l,��\O��Ǒ���7��0��(�Q.�
tAF��*�-�vU�Q��s빓�cE��k����K�,��GΕU�n�xnd�R��t-4�'1�4���Z���<&ރ�����;�S�8�Z:�(� ����~3e&��+�
� }�l�?b�\-?)
�#�ƨ-�0H"����S�*#��KN�+	�G��Y�XD6����n�o�'y��J^¶/8�i��x#�} ��Q��������?Jv4X}���M�U��&��u�3�̚� J�������q�e�,?�W������94!c� /[�_&�˟�.��ث��)�V����5�>c�� �?5���G3�?� %度��u���i��(���`~���}1-J�W��*���iK���'�� ��+���[mҫ�����ZÍ�q5o�`R�rtD�m�߰ug�GA�AyK��M���{��h�z:�VQ�I.�\{",ٿ(
}de�y6�SW����t����94L`֤�\�|�ݼ7���=Iw4>r9��_�s���ǎ^�/��f]dky��?>�?t0|B��w)������N~����,{�#۩�d�i�{�ݎ�_6z�r�lQԿ5�Fpp�P�����d�~��N�W��\`ג-%w/�s2|p��%*�v4��Aj����g�R�vb���«���I��(��ƭ���B�����JF���9����x�C�Y�>�Z��h�Z� �o�)�����Ż$�Ri��ʀ���m��m� z댗���lV�H���T��,[}��p7_�D�`��x3����CCx�ǘ�L^�~c����v.��nt.w��[�A�:��]~�&T:~����0�Ѡ�I�s�/l�@�mkp��n�~��L�9���e�>f�P+�ũ�MǸ�	_�Mu}�6�D V�Υ|�6o1�����G�G���P�V!�>o@$CG�|��h�p�H��S�\��RW��W9�t��"�U��wmsA2�;��ݘ/k��8����v��.#6t�| ��J̅����亀�����y�
@���v�&i��6S哢�)�O�{���=Z/D	���b)Qj�܆|����}��[�|��2�k%B}�]�#xbݼ_��O1��<^�k�����@���ܷ�pC�$W�L��'��m�P �,V��J��qB�4�m!��:,>0~\"􃟐���sjH���[�pno�A?dmn�ٴ����PէnM�vzdqc�i�$~p���Y�Y�G����� �:�[=��� |5�PVa$��fB���}ʻ�$:1SF%�l`֤lj���)�RSdH�C���/�ƞ�9F2�鉂
��&�X�h�7yQ!�}e_F�>��1%+F��z2�V���H��� ��4�;����㋘�ԸM�g�]ɺ��]��痓=��9��\?�.�@�Db��SP����44��� ���6Ͳ#�Ms�mVK�>�(�v}N���gC����\�-�l�뉙sZQPc��}E"��d���1��mn�  �Cg��K A�#M�H$��#(]m��p8����6�S��@eYZ�|i�2�O��R�xCd��6�@B{�������`J��,�8�K�u�T�
������3�X��;���0Q�8aQ���B4̢��?�FP�����'��ΔM��d~��a^R�3���s��G�T���m�r}��%��}2�P�פ�;�J�2-ٌ0-���#2�yl�(TN��J�v!�]$�yC�2�p/Z��>�����ڬ%�Z3�=��9۫�z'�g�_��!Q�x+�n�R�~C3ܗ�����%j���q�a��\ ��ё9��u̿�]bN���Q}@���jO��d�9/	��n	��ؿ������ı'�긏b�>�)W�3�X=h���)m��N�$��	�~㭖]�U�s Hn��Ey!l��{ն�Qo��)�����e����Z�ݝ��
�՟�C�+?���W����j:��T�?���Q��b�D���8��x���2�K�^��(]�ًq!�,`��l5'r}i����q쾕($�"�R�J�7��ŭT��Z��-\jKM�z��W�dk౏f���k��c�[��õO%���3�q��گ�a�]�x$��� �|�HukqY�����ɖ.E��tn8\��7�`��s��ۦ7Q�?��)�I����7yG��S���/?��m2�d����լS�2��B�W(��.���I!�#�ZaOL���%��ءd����rd�+K�Ѓ���{9�5b����i�V����P���Q�V<�)��U��=��W���E�=+2�� ê@�LG�����9u ��B�L��m�,��n��`ڸ^�kє���O	2G6����Dw3�@߆�S�C���٥ц ŉ\K95�H˭���.���HK��4}ـ���C��1s��G2b���Bӑ� �1�ۦpM��U�����'$� ���ry���y)Hӛ��ػ-n��Y�������� Z�GI�)��Z��t1n><w��;�^/`!��{�|TA>�xac�!,�j��'��\�L�*�a�F�N1�U�)����߬_^��ށ���9�:vg���0n_�Z��T�iNZ���m�: �HU��X�F�1�13�b�c�T��0��IiWng!H6a��F �q5'��\kz���;�Լ],(*%��<n�0���4]�2,nb�����5�Z��7@������(i`���,�]s� ����j�U��fD��0�wtx�꟝̷o�Y�	Q̇mzK��̀��z*g2c����}�S����#Պ	�ʺ�؈K������j�ֳ�]� U�1h��� h��BhT�o�࢘����)~�IE�Q�f���5k��0��0�0�^��\/��cBA5/.�*�n�W�L�eJ�D�h����u�}�z��f�׶�t�g(�ݭ���o�0-ˇ����HHv�{��4�B�[����-���~���CN��eѓ�h�4[�&rF��J��Y��C��մ�!����u���!��!��3��R^�H%lM�4���D����2`
W�NhP����iR◤��(B]���h�E�8�/^�!���}��/�V��:B*pb�*�1���Lo��8�]����ϨU��|~�T��.��RB�N��/wÝ�j��U����t�m��b�bn��E��d<����=7">��~dbri#���p���L�:���h�"?4��	}��Y_Wt}����(sxa]�.��ǹ�VF�^&]�NɊ�=�p�,p�΁;�y.�w�&m�T�&�qӮ��F��џ�K���.���{��7>`T�P�������x8��g�-W��(�KMu+#�t�Al#CO}�@�V���{�l㉋��FN7K�&�!Q��R�g?a����5��A��=�D)"�B�u_=�v��B�R.%Q��F�0���(����Aq]�R[��<?�#eAG�Y���EB�V�󲒤��O
�T����}B�¼RV��S��Xs�'���L׵U����t5�����R�j`���!�4`q3,
��ޱ��E�g�kU�umR����Z�'�S�(�5�k{�nݪ���kN��3�x^�����`m��I���#�K�h�9��є"FJ�������آ�h���T#>�nl�X{�0����i�#��}��d]��Y�o�<����A%$WF�߮�X������'���K<�x�HJ�l�6Q�M���X[s2x݁���/�܆�Y:�yn<=)�D�{^t>�)������$S����~�v:6�-A��Yܑ�h &�<u��mtD�7�U6��`�`����1��gv@ߢ��˩l��$��w+���R��|08���#ȱO��6�"CV��,j�J���Äӭ��˒���ƟAH'�����;��y;��vMJS���������[ ��w^L�䖛M�)7���r`x2״�y�7ɦP �ZGG^V��aJ�~/���]�]|��J�b���H�V�f��m�K_��������V�2i����&��H�>��7h�����.��0����i0|��&��IGh(��G燘������kfAT�E� ��t�_�NE�d.����f���~z���K8�|�9��S���,i��TPJ<w��l����MTǎ\�v���2۩7�9��ONDmD�v�6DV�D�a����p[�mJ��p�{]V��������9Vo����Q(߫�u��i\�XO�N�1���}?�@ߦ_;�6��C���,�c��z�-�Un����L��9��QQ�%�^��7<��	55��rOm�C��$���)���2�2%Q��=t0g%��k��� 2K-yQ�u�"ׁ��W=O���y��F[w3�zR(�D����G�q��j�#n��3���u��bZq��i�����"���ߴW��u})�ɞ�P�r��� ǢHE�	g�I�JEڌ��O����n�k1Y�8���;��S�X�:5� F�}yG��8l����u������x@���+I &�HCP �.p\6;v6���?�$~�*�L� �C�j�a��Ioמ��	�GU��F3pɪ[�e��~��Y��^���dH3��WD��M���eu�{��)*�"Iy�����׌7���F/Sv���ڕC�*�#�6�S��PGZ����%�>iQ*Rã	��1���}�;����Æt�Zo�1������Rc����['�]���C4/<�d���j����V�~�м���P��T��1G�J@&��b�V�f�S���X�\\�,3n˝��<J�����8Vo�L��`c�R��$�jGA �
u+^��s�ħ�1�<|H�o��|'�������l��<�S��`��BKft����C ��N�%�B��_1<�vbR��1����1���,�J>ЩNT����Z�N!������f���nV}oö}J��D#j-9�8&��w�2�h,��.Vx%	L���+;�!.IJ�*̠{r�g�e߅_P�@ڙ\p��� ��J2
X����w����o���R��M�m��a=��=D�Mp�c9c��s9�+�y�9����$�����`��	V�I�M��M�4�!�v����>��]T������o����ǟd��]+tW �D�^��m��I��4�p=k�6DU�-�!�Kh4�H�K�
ʰN_#��L��JrVE����ѷ�A�0��n(lh5�~ p�`U�z��΀�(��yD�c�	�Tp$��;�:��T-�b9NH�:"{h����V4��-���%�h�C2u�Z����l�-�D�]��b�84�;fIX�p�)
���c;�%��nm�������v$k
/�%����Y&�l��y6W�ջ�zUz�r���]���5q��'J`U��\�pH���1:�!�H��OnZ�2n�}L|$h�w��̙,hN�S%1<��ΰdWK�Z�u礢S���{�+M'h�h�7h��;���#i����h���F��B!���r]¥tޗ��\�Pq0����x�w��P(���b��7wu��
~����Ql�D���,N�H��-N�i�g�<������<�cOY���go�	[^q=>X�;i�v6�3,|Vxo}\Z������Q��Y�*�<�a���X���|������`jo�����3G*��F��_�[wF��D@t),ص�b�ߏ��4�b�'�������'M&Ƃ月 �@Ij�,T��i����cd%js^�"�<zMO>�5���;�Q�H�-�ȗ�LMnP7M�.F1tHpl�=���FpVn��
5whP3yF��#nD��mF%�G��W�n�=`xa�׸��)+-&�p�f��S�� �
\DD,wSw�?/ӫ�Lԛ�6��U5l��C��ż,f?'�`�pEC�-ic|�!�W��� �n{d�4��`����]���)ǎ�����[�̓?�w�@�Z���~�7����Ja�'������X����qߩ��"��ǘ&>��o.�s��ںΓ�~$k��b�c`�6i!1$��r<󛊸�1��o����N��"�X��F�lo����Q4 �@%_3��h4� ��5���ok���p�@_� ��h����0�"�FJ��6U��-?S����������BJ4��%�AeZ�Ev�J��2�+U�\��UWo�7��>�E�����g�e\}��@�7�S;XM\Y*"dL^fd��v��I,�V�� ���^��e_�I�j��
�����8�`��Yb���I�eor1?�&�}pX�sC���N�gJ"��S�#���JĚ8~��k,��~���X����i9Ez,��k�ށB&^��'���ڥƽ��0�SfY�0�PU>�9��|�0)��$���(��|��'5��]>�[@n4�0O��^����#w�w�WMcxt���a�	!�z�E�����F�Cg�FD3f�OeM�vXM1]�� $��a��2���˒�4w 0aY��a8�A�	X���y����ؓ1�I^�]��9����_��3&u�uq�5��P�
|���RY�9֋[��i�@��M�k�'�9�0"^r��h���#�)�o��`V3���	5�%^-�n�:>� �姣	�"J��&�!��W�/F������B�5CdexF��m\�qj�b�
�]�����:Fr$�ZU��(.	VlԡA[^�D
J�3C!�3�Ga:n
�m�@�E�?��T�2�$ �Q���jk�@�T�U��r����{�0���� &�����Y�Y�{�~(�b;�N@��)FM;�V��[vC�[#u��$��YݮP�j*񝴔0:��X�]��g��iT�4�a��ۅ������B��s"�:��,?<yl)�3�YN��aP����6PTa�iRI�_8P_��h����D�1~�ϔ���Y��'n�I?���7������Rg�8;X����7��#�b�`�[6*�0./���G=�[����}AF�0��XLy��������z���9s�bRHm���V���YRMz�Jg��g��ZC�*����ր�+L=`���f�/��������倲y+���u�H�{���pwzj��e'�ͯ�75�o+���,Γ򖵘�I�����7`�v"-B�Y;'@f1��[�<_\[�c��V�ˌ���PI��N��td�R�E����Γw��ϠiJ=�+�\R����~d_��Ϛ����1]�S����m��&�ԳSc;=C��=�D��+����^���]��R��Z[��J�u~���P�U)�,��I����A�Ns�K�����n��ױ���&�������T6��=�e�"o��rd�K��f]��q��w"=]* �qqYJ6����j�=A��J��a�D�J~��|Mc���S�����<v�/@y��%� �I�j>˵\}�d��ey�(��*T']19V;ڎE��vPH~+�\�y�8s<b���VmxEڗ2><Y�x01(��;J�#�%�&Ε�$�Z)s].����)/
��8������%\,�T%��z�� �˻� -W�	�}5��o��Ϡ��0K�'�2����țP����#�=��Sp��C��?�f�,�'��V���{��yo�-���L�k���v�����a{���֡�E�-O#�����HPEO+�{��	:ϢJ�z�n.�lr�Ȃ�B�M��ބ_�-���!�9;)N�Àl��̈�Dt����c�L�����'�s�e�l� �'��K�<O�z�s;%n�M��Lr�R֤�A��Ҽ�^���Ņ�ٲ�e��/�,m�@�����*P��
�t�� ��_��Ӿ��1x�$g�ܶ"\�3$()C-��ȅ �MO�������4�k�y����ZM(�#��/都��SsѾ��>!�A��ytK��נ��r�Qr�<,���1 ��w�5�
����T�b���!�Gi��^lj�h�y0�����m[*O�j���L�E�������l��S�u����Sf�W�f74�w�1Xl�ȝ/�E�y���Pe-�
;t�m�X7��O?��k]��֗�2��"P¾$��T�ZMԶ筆�
h ��G��A�����OGp����gn�V����������-���m�Q-XL���z�f�B��g�kG��W��5!u�0�n���jH�����S7&��
6�f>�(,��MF�s�j�!�� ߜ~\�iNDv���;pro?�
�6��R.Jv��l���d�Ν3�[�����&.LP�����Pf@]W�2.E�@]��-|t�+\���d)��6wD:��m��w�����7�*�HǓɀLNz��b�0��@y�ؾ���bն>�8�7��Fg��/�s6�z��E��Ra�"���}�w6.�n��@��ɧB���χx����$�\�!��o�E�
u�g;�m�>R#|�q������zvHر&�QŻ^�T����O7�,�$���A���!��Aƕ�������s�Dvϛ"g�e�=Q|���M�^�4φ[(�^�?�1�3�ւ��ݾ����H��ؔ��� �0��M��M4}r2㢳[�)2�ws���S��.��� ��u�O7LQ�l���j�������som�)c)���!�S��g���;Ks�m3'�S{%��\ ��z�D���篟C��H�l��4.n��i�R�&��l��T�?6�$����g*#H/	[�sa`��ŷ\�Ңƭ�92�z�C)D�I��r����֔���ET"��?�|e	FJ���Y�@��
_�.S;c��p��XCǹ�RRܽdIWL�YlO��Z�"�y�4+��]��R�,������5�4b��� ��cnB��1PW�ș)g_��$�<�Ӫ�M.,��-�²��&���ۃ���5I���/� �f��օ��N��7~�&E�{�pr��B_�r!�)�3����_�s����׍������(�_D��>o3R�w(���Ɂ!n���N�Ph�|�%��^!�p�����ar0�Rl�`L[s���6LM�K�\iR�N��.!�2m��[���3�v��Jc���j��W�>���S���g��Pn%\��g��&��f��-��������+!�����Ve%�q��}��^��O����!�@��ܵ.:�ɸ�S�hb7���OÍ�T8"3].��T�.I�`�#��jP
�)��ݡ�9� ��/{8�ԅH�Y��A�o�jz��Ӷ�.�L��'�� ����xH����y�x�����\K>�":�t5"���qS�-X��n˂kp�%尓�J	C'�����c�O=;(h�.1>WQ��{�1�p{��#�{f��D��A�w:���T<m�^��^������0���
ƳH�3�ޡ���+��9+ŁE1��}���2Сcc�*ϰ��!y,m��-��!q�;�hɛ�LG�a��`!�*���_���2ԏ�_A�q�%�%�i�8݉G�F���u�p���x�yz�1NYR�#���g��� Í�:�t|S���~<��G��(��cE�e����VM
M����)JC�c�6
�6ʙ4���64W�ȏ�DmNS��@���4�%G�*���k��*b�W`�f�����0n��ȴs�M\1Q	8����n}:t��J���"z������Sa��y���)�f'Ӌc��^��=�.����XM���;])����f7���CM���M�X,���Rތ�������^ͣ�� q��o�8ijG��-��]�����v�<`�l�#�/-���3c2cϟ{D��!�r �j���-�ʚ��o"�jq��>���������G��i��Z����
����@D�����Xy�F��.=�$�(u� �*'[�ݽK��͖��O_͘�_ߪG�Hy��@nL�sHB�@�
�=O�lu��:<	@�9���8eM,c��,{Ȧߨ&�l�yrr8A�(�VRz�re�.-�Z^��\�E�ֈ�:?~�S=az�7��������	k!�����zYt��
Bo�E����ar���Z���A
���V�`�;\�/�Ux��yQ� �d���kJ6�����-c�R����0̼ ��?�a�s�\]�l(���l|�v�*(Ɂr������_NH7��M����- ���'���46�c�3��<ιD�Ç
��������U��m��Y�TE(��._)����hD}czyP�������6�\W�9cz͉��p����Z������@��OC��;Қ��ֹ@m\�.�/@Sh	)�g(�~b��܆�;iA�!�j���q��7����,(қ�_oY�Ʃ%A*�ng�an�,P�1�<�H�RXVظ��pHm�J�<�I��fײ[8w?�=Z�Q�ް7��_ow���;��۴~�e��^3yk�C3
��#��^{�x[�R�`R����	���R��
9oj�yV�R��K�����:
��@�B��$�7#E���M��{�2g�피����v�"ej��R��(���W&n_��8j�O�r/��A�^"�m>�o�XM��1��~;,����"D��x�Æ���fAJ����CѮ$�d�eM>�|�Ё?�O1�qTT��d�x�?�� �ĸE�&�J�s>q(y�Y�(�Q�h���n���{G���Xf�n��'�:!�7�u4-� `ݞ��Y�u ����<�\���r��?�6�Sh�@�9���y#N���fN�V�R����堨0����ܯ@�����u�D�� �l����������֧�k�#�6�2��*O����c�=x�v	����O��z��G���LW��W��@\��kʄT
����WH)�鸄vǺ��š�������<&#�ml�y:�zۀ���D�Zm��^�&�N�8��X���T�K]�ή�{:��g�o�;�w@�e葻��?P݂S��7�Kv�v7��q<�Fw?I����Lp�m]��ģ[�X7�:nI/Ho^Ddwۜ�@����Z�ѳ��/e��R���j��<�����gQ*i��EL�.
3_3���ipb����N���ݛu���m���a�Ll�}Ax�V�~�l[�U9Wh��/��+�uՋ4���L=�xU��]��g�9�/@ѝ-��2�?�CL���Y�1�p�Y� n�W���)H��A�`L���D�d^�"Q/ǨQ���ےuO����)A��Q�Q��0T��䒝���2eh�1B���,���b�V�ki�s��h�Y8F���r]d��r�HC�^�����O~���@ڑ�YB��ZR�BiGt�b~$���(����:׊�Ʋ��J�ʽ��lO����?�ԋ���n��m�D�/�+
���\���S���_.V�h�jh7�(���K�W��w�
��̧b��܂7��3���*��:k
�u������Mڳ��-G�U�/�&$��VG�:�y�H���X&����r��%^t�2�l���
d��O㦅w8�A�G�:ߝ'�еC]{y_�p�OJ��~�9�o���f�x?zx���fF��m��և�>�ch�bg\�&���-0�'�ޅƚ`��y�*zوW�C�@�z�y�����;��?eb��`����Ӳ�C�n��b�jP��,��p1T�%w�&�W�z�X��ű��D.�!lfF�Y���C��L}��K�e)OI�
��Z؆���5	��6��]�ޣ]�)�l�g����̱C��	��*�s�6:�_��\��VfJ0�Ԩ�k��w���[�T�[�f���nо#竐���G�97�B���w�X{*^P��V��Nn�@?�C�/䒛(�Ճ������mװ��M�}�{�yt�Ϸ�`�-d��'6�Y�L䒭%��{2��,�%LN���t����E�+yA��&j'�x��	��Z^h��7�H�N��UXbj�>!þ��T��Q����K��*�1bg�i�Hfའ��*e��$
qN�݄���IT�R~J��Q�����8�a6_AK���A�s�qx���/���g����Л�6�d�?���&bG�%�:��k2rT̡M��o�%hYEw�6\���+��C%�ȍ�D�~B��f����a&�,5����]��x�k�6�D_�pA� �-����_�̹q�6�S���P,U�����Q�!BD���=��Pܠ���1v��9|^�Ո��%�8��T���nA:���_?��|Ӹ3vmL��x_<Z{6�kf�a��c95��rm�g=_��I�xҀ,�It�q�Õ�������}�N�u�?��ZE���=����~�6� L����(ӓ����:�Z�r4f�f�`�'�B�a�!�C�}���o&az�f]���4���	����`G�hՌ����S�~3����Rn�z9�]M�4q>��������ܰ��ޖ��M�ӀX�5��þ*�`�曈O�_��ۗ���.p�;s͖r
��_�M�|�{bϏQ{�4[�. :�x0.�E}L��m����5�V�xd�@s���te�wS�'x�	�i�i%G�����@%k��J��W�h�Ti�u���M&�o�mS����"���&��j�<�ߓ���W3��M�^�䫛^��<\�������xR+�Q�}]�����[�o�z�Bԗ�q�Q1�p��޹���_Yf���ۋԷu��	N#�Gܐ�w�^�~���F^����jT�u����Z["g�%��1t�D"�H���O���PW�r�Ww�0y�DW<�V�4Uط�ϝ?���.��f��Z�x`a����
p<5>��fS'K��ELt,��f{��k����4���!���%ڈ.I�6rԊ��p�ν$�]q~"�N�9:��8Q U�e?ӧ�9fJ�a��Q ��Lٕ��[y%y�������G���@�<��P���a�dm���`�C����W�>��V�93��0�r�w���$MC�h8�cr�R�m'{#��>�1R��q�[{Z�z�=L�k�߸5=E���6N����� \�T�%D;��
�iH+Ni���W����F��W.�I��V���?�}H*b,���w$��Ts��k��^b��g�YZʬ��r��9�iZ����Ł��	w�8��F��ً(�=a�{�UymB��x��Q��9��t<�����5�� ��z�IE@�A7�!ߔ�0��Xp�c,Z%Aٟ.9C�.1�I 7��x� ϊo��y�H��Ѷ0��}�̠�ʓh:d�#��7eaڠ߅��N�z���H��k�Q�oՏ�"��ej2R_6�P.½��G`w�SR�Q`8*Ǒ|W�o�V_��Q��$� �?5e�y�uCl9^H0#��� �e��U�S�ph��j��P���߳�I�YE��1�jqy�������̘y��{P7�#����[�z�
0%��������J�-��jX��<�$���S�r����wR]�Q���ߋN]��<%B���ߞ!r�/���RHM�(��X%�ޥ�T�qc΅�d�ݍ���z�7��xӹ��
���NP�e������wۏ��?�������p�JE�FS]eP�dX�#�F�=,��� �7M|P)o�ᐹGG>�)�>�[A:���~BtP{��׾�z��.���J���D�DN1�K��Ms��@�ݑ�JHk�)�Q�h/G�2��
˾y�{�s�C+�\w�SP#c4lz�tw�L�����$L��N�D�X����g1/�
8|�]�/�fJ���F�Z0��]e���4ƽ�L�#-��n�A��=���L�Q<��Z;X����S͏�T<w�������ƧA��ԥ�7�Z�y��u���YlX�9�x��A���"eN�:�6_D4p��/�} #�&8�0�[�fn����̡�-7�f8�aw���2i��l�R�1��2���L&6f�d���qK�VX t���{���¹���m��qF���������kW�U���U�:�m%��b�xH��aQ��|��4�&�[�S�<��0^��O��	�i��&˥z�;��8u�!��N���G	���и��b�B\��ۼ-˓j�#5��`����a�@ќn�fuG���:����N��'��0���A~&)�Ū_��Ni�`�����`_��T�V8#L�"b��fËL��ثЈf�nF�~Վ{c��Qa�6������8�:���c7�.h��M�cr���ď�s�V,����F�W�w΢��ϜM'\�ݟM�ڡ��(
�cX%�����A��'-֘�y0���Ϋ�o����X,���H��`��!N웶%�]d�]���d�8�9d�TZ�]'�\-��F�
G��p,g�y!�3Uc�E���_��b�|x����]�a 0=�X!	�����+-�sb�;��W|%%�VRh��i�E��S(�n��o޷���a�TU�ҊYn#6=���4I&�Q��QT+�g�t��H���[9�O�}�t�|�Q�\I��&��Yh�N�(�]E4\��0�֩I��)��Mk:��]x^����Lh�0���]��(��"!�'���� m͔��D�`e Ɠx߮��3d���K��Nܚ���:m
h�+��A{�=m�©�ƫ�%���XXjQk	�z.đWw�(�j|iQ�XJ���J�}�K��Kу1�Ws��G�W!�P�E��馛�L���am��ZIP��6�x+�Q���ZKp7x�r8	�KH��t����i�i�A��p��3.�d��0�!OG��,�a ���R�QVQ�a�F���E��Ax�(�@��!.r�|��ݙ�a?���W:��	��z=�]�,�\��O��*:���TVJ_�ilq�bud'�Y�ۤK.h���̥,��h�<��#�k(+ZeЊ���]z �|u.����i%yb�4vK�de�������C���������cM}����:^txrF��]<};Q�����X��K�>�̥�!�`ţ�U�p}u>����	��d> �n垅�&8�5��P��Dgp�q��RF��2���Uz��U��KBAQy�Ў!�zj��� /X��5��Y�N�!�YFX���q�,_�$R��rK3�fbD���w��Ք���|��>���1���s���i���	�y�����
��X�Ն�_���*sg�r i7C���=�������ζa te��r��o���^N��,A�O���v}��c�C���n˟��g*8�$�8�y���i�Rf?������(1F�q�([8�C���VY���y"�o0��u$��#<�Xy�Kx ݭD�s��U�߭�}�OkFj�	��K� ���W�R����~S�!�`�����Y�S�	=���hRW��o5E+�ҷ.#�xr�e�wĒXAԮb��E?��U;C��?佢�R�����i	=�i`�l��]�c�f4���m���*7���u!_h{��9�j� p�����A���P�s����]�NK�Q^#*����(�ا�\�;� ��"�@�����CaQ3�>�}���X�!0�L��
Ҍi�j;�*���vs+�'�ݩ-��ڹ��@;�@	dm1��J�S8���,pe%x.>��0[�g����UbK)M�1�۞��98}sӦ���S��%g>:�Q#v��t��lP�Ce�(:�L���9=�5ܙ�%�D|/CWMeXy��X�-M����,�����_�Y�W
� ���ev��7�I���H��<N����:�_v�*���L�8_��V��Pn]VeG���ؼ��ծ��[}�b�f���Y4�Unɔp����a�=��N8Ƈ�@ �<�&�CL(:��^��2�Ғ�Z,[�ȥ��b�K���_A�ݢcː&Y��s ���2�-w�=C�V��	�;�f���8�j&Q`߾p�ɪ@�$F�)g���	ESXG�^b��/3��ve����b�^0��}�Fl��=y�%��1���#�nA���87���U&�����>;��'~Vy�%_I �4�T����a��U��4�/u���}�.ӧ��E�N���*�b�f7cO|�Aֻ��B�
�J��H#( ��8�cֽ��&�������E����w�J�NԘ��=� OK�p�8�ˎu�&��vQ���Fn�>cR �ڑ��ֿC%��+
���>0�/j*��s�#��.������'<W�z�3�ж�ɤ)�0�*�����on9}�
;��r�W�� \�j��D*DXJU��b_��5^��F{�������� �+"��I�L��r{����VI�"#6���6��k4妒.�o9T���x����7��j�/חì���ұ!�6S}���#�jt/�NG %�����v��V�n�x���ܒ�V��X��>!��0���P:���x��P	HvؚH���i4�YՋ��Z��"�����S �ٌ����ݧGK����	��8�K#�o2_���������v^�M����O�K��"��Vh�y��ֳ��{jb������Xar��v�q��#�Z��f���2���n��"��Lg~�+�$8>kxsOZ#ǆ�Y+�	ǯ�K�
ݎX�Y�\��_6�!��=6��8Ke��<�����x=�Y�:QyX[v*��.�*��f���fz~`���l�jm�LA�]��f������������(���T���U���4U,����_{د�� 1V.��GJT1�%�\O���<�7��|��3�]�IKN��W'�8�����Y�/�%v��"HB��Cr�6$�!0�
Z��N
+����I��:����}a�:���4��Si.?�;*�GD��DN��� ޖ��D�V�%��{>)T�;�	XD���x�`�5$��U9g��h�.>v��o#a�t
'��0�Nω	ן�o��_K=^�_�Z�X00��,��`,���)����6�HqC��k #�@jm�8���T ��	͜(���b@l�@Au�^T��e1�5�1n��Z�ˁ�� ��Hp�ٚsCe� �����7�ev�%*��Bu�� 7���Ug.���w���?�=�swP�a�?�?��G/��I����K���_;H�{�m����l��E[��V�!tO���d��2�#��`O�
�i'���^v��8���b�A{�G]e���
�l]س�VtN����j�w 2�U��G��Cmw7��k�Z-w�sׄ\\�":���	�\7��'ԡ�.������F������rE+wE ���W^�i��1*fʝ��
�����S�Y��Ĉ�.��I�*94L]PZ��T�x��'-��CB p�,�fF�%pa���d�^n���	M=g6%3�%�CD�4�	<୰�&${��-�L8-�Tu�@�uy˾�e��s��~&�?�0 ���"�����N�����u��b�Z�#w}^��:�N��Kl�4���tt��F);�h�K�/ӻ�̥wzWv�$P|��q����Gzd�@.hs�9�'�i����������ځ+��D*�������N���8P�:���@x��H2�V����e7A��">@��>Z�b_���j�[�%�}rT�K�z�9���DMm��?Byi{G��[2�F��rt��ynD|_�>����'5,H�s� �y���D��D"��9��>��}s�oD���:�S&9y��O2����m��.�r `��u��4��	�w���o�PM��v��M��C�#��_^q�*�o����Fs����Q��8Pi�NCz��B:�a<m�$s���4~���M��G�gc�G���6�I�TZҬ����)�Di�ė���k��f�Ș)ϿI��]�כn�>��!VhM%�iZIuT��j@}ch�����Յ�Qpp�<��n5��'�z&�<G?se��RY�����F�A�1#��D3����ʝ;�E��A�r#|�������k׾�s�p"���s	���K�e{Wg�	.���������ܺ�C�	����"bk8��h�W\���l*h7���
x�����*A�a�R/Ǖr&b� ����j��|M�=�ʔe�̀J��uLH��&tF�`�	7\/��}Mռ�1�|��3D@�X�Ã���^�&��c�"�o�WQQu�x�;�{�����
��gKMb��7�\fh7V���h�6K�����;�"�`JWXڡ�Sp����o���7�#=�3��Y8T� ��8Tl�����:�)��YLsYQP__!6k�߈
�ە�M�o�H�ޜ��"bƜ�s6�zWH[�h�d�吸���y�M�.˯PH5?6X=#��^�UJ!2gTw@���n�W�5�?,m��f$k�nz�Md�0��;���ԩ�?�l E��Mo�H:�wS��A9 |���ixY;��C�8�լ@F�>�cY��J* �}�)'N)�:8F�&F;ͫ�B��::��h
n��w�A��K��ၖ�����^H�M�.1�R쐟��Xb�(<T���G�H$,9������3���)�Ib�'�Զ��	&�ɻx�f��x� �O���z<�i�RWb�5Tu���rd��"}N�Co���Q榴���"�ϫ{u�=>�3J�7�E*��ē5�����3O��.Q��@��w��6�%B����Q�����]8�o���.�4��2�ф��>KAm+��X�sr���4؎��voQ!d���>��I�?fM��mc�Ds�m�a-�Nͱ��D�\~I��3�Hh��\����?�!o����I	_yA��N��߉�HhC.-���@NfTH�y�<h�b.���!��M��`$��9��W.���k5vv�G��.mx��\tS\�*�3�r���cĝ��k��G�[�O�3��#�[R�s�g��������l�ғƴ�%S�h�I8O�A'�BPԖ��[�4�<������Wd���$�Edۖ�����x��8�1��@t��N��s�?M��PLH�9���[��q� 9[��t�慣�L�,����k�)�lob�@���P)�,�B���3��`/���F��j5T_�Ko�x�]�_l=����6���C�L�ݛ�AW�?t-2�SAP���t�=.� t&t�?�*L�C���z��?ސ��a��%A�"�댛�T6�^�vmG4���MA&L��5��0��_���$ t�Cަe~ިNa�+c�Ț5�l:�8�D��=�����/����J4l^��)Q1�2�=Z�{��>%�pt����4�� ''p�ߋd!�XY�� 54_�7��{����<�������_lR����)�5d1n��
fm��v�fo�A�?�5�X��գ!�� mѪ"��5�)�m~G�� (��B�hJLW�k�vW�\���?n���<����r���UKۿ :[�SQ���庪/�+Fc���,�
��#�:k�*���yu����O�d��n�#$�c?�	
_Zش;i@8	b���"��{��L�o~��ъ�n�z�"�?�����HRǔ1�izV�4<%���oM�XԾ-�~��Xg�׍����t�;y���Y�kR��}PC���bڄ)�32��j��g	w�?Ū�r4���:P3u��sJ�X������
��VTz��~����z����3
����w�&�ct�]K�6��s�az� a�oO�
�z\M�tv��t@��q�2��w�?����-�,�Uru+����5`���%�3�-,v���W�+"-������R�E�^�}$����+�k��2Uv0r�;.�m���l��n�(#��4l7>!�;&�G4���"*/]�ʻ�U� �Q��0
H���{1hZ��TL�'W7H?�ٞی��X�3�G;]�&�8dS������٘�#�j���t��Y1���tb{�����D�#a.��(3<����"���\܅�[4�L��|Ֆ���A�4w�p�G4oDXI��dA��
I�^�BKa	���Ih��ʩd���8s���Coޓ�q6c�����Yɘ�ǟ�D���������݌ٲ�w��?���H��WG�E�c�lo���wH>G�hge�8�P�2�#��5d�τ�$��j��%�+=�@A�FC%)$A�(F_�-t˺6g�[�un*��7Qk��E�O\~����h�1ϴ���R��P%Fi?hݣ���:⹥��O%{����hUk��ͥ;;�=����ݫ���PP$�nx}�fR��v���0�h��� �>�^�jM�`�����d��e'O+�-a#a���p!�H*#�5�V�6�~'�s�J�����<����4m�Q��.�a���^xrZ��R��E�	���O�jj9�o�������Qy�p�3��r9���-t�kc
���$ZP���]�S�:���U���_p�Y_1�[��A�Kz�a4� �lszG=zSI���y�����C˓�<k4����6����#���q�1����Ҭlc3�o[�,|�kQߙ�~u:
��w����[��F���Gd^�����Bb��/�F�h�h��#�����)?����y���ĭ$�_�'D�T2h��@S#lK����F�DL��e�(���  lK���/{�2܏�-T�ٺ>�|;�e���DNy�}�T�C��Rh���Iv�l�(�_�����A='lbu�8C�y9ʒ-�F��7��mHxD��w� �0�{��/ژ�
��v�*!;6:�6�t	a�C�5JK���)�	��I�/�=eؿ}��!�Q8ܭ
����s;�§�}yS���2j�O��
���z���)��'kG�
w��`�T;��q��b�21qy-;ڧ��������ͼ2���{��[��s��F�(�K_�ey�>-��[�>y]E�ոF5�B�>�E#�(h��������9�0@%,	aŗ�E�aYL�*�LCg7W��x����@uL��Y��GG��6~�a���^�*ߎXA�u)�6ο����Y�/�B�3r���/c��=���L� {]�����n����
�"4��n���3��|�}d�(�֒]!wh�J�`���M�L`�nd7�o�!����F�^H�?N������9Ր��c���,�i8��`�'����y'�12�ȀV��< �Hi�8�cI����Yڝr�'!��94UO-�I(��Ԛ���9�MEl��.M�>��~6�ۡ[�aI���ЭݡY�BE�3��S,���&v�&lv6����i_L�}/�)5���D���^���H�1Uh��S�vZ���ѺimJ_�N�?6� lX�\Mm��F�0�y~�4$�ra�B9k_�O��7,�y��N:�4��/]�	y�t��*p��x���F��U���rl�*���IJ�S�?d����.D�j%7 ��� k�isxZX+�H�#���F�U^2�,�������� PU!8��m�oc���^#�,���4����n>w���O�z��={�� !�^I��I�o��cz5�/���vF�b�'�u@�2�v��65��J�[>��� ��4�Uy4+�..���"��.F�u^6F{�)�V�	����|\^��h��Q��D:�˧�Ț�B�:d[�īV~8�9Ab����r���޽��_ƐCu+�W����cR��3��j�-2oM��˾ 7c���$�-k�bអN]�K؏G�N�3�Ĭ"��`�)�'Jχ��2�k]:s����Y9�Ѐ�#�����fE���[�0������7�5��s����f���\�y��e������?��J�m��15���Я����@����R�q��'�a�HQN�d�vC�c	����v;N��* ��v\���M�%� pj�PR݌���tϒ�ʴͯ.l�_~n��Z���@ի��B����fa���z��8�	��[�c�Ԧ�y4���F��GaZK�Jg��G\���E~{�MB�﴾��]�ľ3�ޗ�QO��6�8.�Z����̏}�3yX�)�]�����6�����J(᭑��39p���-5Gg sˁZ7���	�z^Cj�,h_N�j�7}Sr���햘��h���j�vH}j�O�PR�@����c�8��P�>x�'Õ6�\m�����:˝<�C�=�d��2r*���s�,�c���ѫ4�����q��W�7�`1e��m����R&�g�Z��/	�p���E J/J�e_��8��aM��?��cc�ܥ�X�=����#�G���lz7�o$��A�jP�&�#������<}̋ީ����AYE��HM%Rb�?�L@�a=\T�4��/(���|B���t�ێr����OV��!��Z�3:0j@��ʺ������m��-�W�T���mN�(�>��E�1��4[!�>+�}�@�����P�%4�/t՛X~kw�W��I9?��������E����m�$���y��t�g��G?�M����0B��4E�{BK �=.EwLSKc4��$��@W8�Rf9#�`cE��@%�jX��L�^yl'��{ܬ�~r*��K���il��$���|Λ�654�:o� ]?kc�n��fth,4rG�K^*���x_O���7{5��O|yp:0�'��@ �!9���Ej�/Zͬt˺4ޖ��B^��=��I����0�E}b<S�N�``�����ˑɻ�߸�{ք8'���R���O1uP`F2&����������)O�\Sʠ�hq�ꐉ�hF� ����4a��A�ݘ�"��֫ZicIq&�.����?/���(h��� �x���"��}fHt�h�%�Y#��,�C�(	�~2>�Øz�^~h=i��ͱ�wi��:K�GK��@E�t���AF�N~C?���[���rU�0NY�0��7������(%i�T#,��𱩤39�]"3���_3�#sޭ��C�2o�
(�q<��G���s���.�y�P0=%��$W�	��e�t����	���0q
�b�9���� dc�c��x�&,{��Y�,@�6H��d&T��]�rS�u�f�����[|��7�kmt�>籍X��0�����Ʃ�כkچ��}���`~�}y�A�����=�ݮ��0m��<O<F q�	��{�f"Ñ`�0��z;�3����\��^��p�����VwB��$�<��4,8*���ߙ��nk�x�«)�����*�-[�溱��X��y�2P��9������I�/�O���λ�oH`3���W ��t�lq����爫�)��U���!jX�pڑ_�C��6?Iߗv�����|g�3����'�I1�A�L�[�Yk�������hc��W�Zd�r�!�"�㟍�@}A�~�2��ah������Hlvi2�!;�"���?b[�n���1���X#���@��
i1�=��,�KyU�[r$�������3g�����<-ZJ0KG�Ϻ�T�U>H5ODYBh���0+W���e�_�$#Eo��~��?�5�f��k��<W�S'	��U�|�}�u�`
~>k-1��a&X� �3��CD����M���y-�
>>u�\�1K�o�_,�KN���z���O˙>�W���{��F� 8����������+����oQ�-���ED�:ž���Rɥ9����p���B�"T��o%���x ��TW����+d���
�d�Y�z||�����pH�f���eg��\��d�,L&�5ŝ��Bxt��j��q�e�;[*z�N[����j�"�����"�v��V7�:���օ,F*��?�n�c�x�g�����T������6�y���-(�
�cC�u'��=fM��"��"��Ѣ ~��_G-��YY����r#�V�B���L��y���o#پ\[�n�D�&.��lY��|,~0a������j\iDc_OL�*�'�ƴ����\]�0^#�\.�a֜��{������l![j�S<�,�/t�.��S���n�������UHns�%�����r,t�C�B�
���P��t��Q�C��o���)o8�W�H�Ɇ-�6YH2P
�RG�o0E�M�\��R 3�o���D�8+fa�a4�ʓYG�h$����wB��b����mH!�2\�e�"��0��*-#K�X�pŽ�K�/t%��/`�𔗎M�g>�=�L`����}�|�G�ʌ��*�!�#]��/�g��ފ���"���@��/
rXS�#��
�~���N g׻.�H�� ��I{y���r�S��?�z3UUƒO�O��޴eAl���$8iؖ�iA9VсAe �o���F�4��� ����G��Ss[xs�8��y���3c��d}���C4k�ϡ�&��<����!_0֕�f_�ږv��xM��-v��c�Q6\�_μ�NIl��/�+e�K~�x��z�r$��!�b��Җ'	à�:��n�g�i>|D��>=�Hh5�6�κWa��:�E��Wp��4��Е��e�C��0?��q�6�)�)��  ��e��y��L9���5���4L��x�)��p��3a�l�f��w�O���]j�w�Oъ�2NКB����GW9����Ma��4��X��|U�HV�� ��/t�K�S��������n@Z|��Zf\���J�S;]^�f���:.��������֓OA��`ͱ�r�hY_X�tH���w ���L-Le,�k�'�Q�����1�5]�|�����go�W�g�Rs��������/��W'�ß��+ôt����GL�t��D8C*��l�L��%[A8�����╀{�h�`&`x���*�&*�w����T!I�E�O�y���Dc���E��&>*�b�F���1��Z��<�g��(���|�>j����)]�B6;(gj�ԎH;�*7b,�t1�!!��^@�,����y��#؞m ��6�x�C��8Y��l8O8�."�G��DTQ�\��N{Ĕ�q��(�gH�f�;�0�K���'��":L��X:�9�#��<�&�;�<��ebm�����0a��j�4,�)4b�W[��\�w�iPy�3}
�h�/]�Ep��O�?�����Y�M�B������[��\���|6+��2R���=�������CNɂsZ���Xo3������@'H�5�ݓ,�W���ʥ�*� )��W�Y�b#�����B�=����
 
�8�L�p�V���I\Q8�3�h`��HJF���EF��K�7�-`4T�N�X�G�$�Sa��(�*���2���� ��2���˪]�$4��Ӳ�E�lt���D�1�g�n���qY���{���C^`�i9ӇL�F+���		I�].��n��wQ��"��w1��ϻw0�*.,w�-@�mlGi����S�.���?R�G sǮD����K�p�_����}h��iD~�x?z��F�ul3-����{�v�q��$�LO���&}�"�����T�� $��ųY����H�� �2�
o�t@�\��J�FDo�����>�v�d�Q#^�g�J���<Y&w���$��ee���VM��ɒ�C����2���d�r���D���{U�G���ʒ����\�ao���K�=P����W���<�YT��ɭ�T������BxԮ[h�3�+O�g�c�#A��`c-� �iIo�Q>1�4��H�y�&S�'ީ��������i�Y����[:���e<���w����}x[U.�P[�Y{sI���3�񸹊�f_߾8��l����!�v��껗4�r��D�ް��9^<4�9�1�N�"����&3�^\h�����k�����>;X"9T��UYG�v���K3��/������P���o�ʴ�6��)E����h��+fd�l�8��9��\r����\������w���6�5�ҎD�,n3�Q?��H�jR�=]���<���z��R��tqnq霩2��U� v���(.��I�W��͚�8�R�Pf���m의��h&�S��i�}��R��S��QZ�ZGpm�$�'�o��JM/���K�="E@5�b�y51�ו=Y��w�]ԑ�E��q����󰀞VV������wND{��+��ቭ�"rF��q�Vb.�߈�nf��i��W�Qz[��?���5�ŀ����`�%Y������k�U�����%�>��9�Lf���Μ�4_oP��H�fA��H|��U��D'��J�LYφ���f�d�A�v6aS&�-&�N@-�Ηy��t�ݦ0+��#eMHi_/,�C&u*6��h����z�5;U��D�ĩ6}q�/U�Q>�E��<^]ӗ�ceN`7ID�vCUU�d�p�N�w�<?��O�Gg���a�"� �2�WNt��5K��$�b_��`Nx�Хz��۴6WL�u�P�6u�g� �I�.�w�����ǐ�N���l��6*ɏW�����ѭR�`�� +U3�i�d:�颦�&��&�<1�ʗҿM�(HH}��/�м-L8� ��Z�IY���ߪ���хS|������N;ɸ6$t�>A�I�B��<�!Ⱥ\m�#fr02N�\���du/��Pl0,�(�p���r���������-�D��ǲqK@V
Tc4`^/캮�ƽ=I�ǆ%��b�-T�F�Ռ� .��B��TNVP�[`Gh�M�Љ�6nkA��e��r'�l������/��2S�1 &�YzÕ׺� �Da?u���[�,��l"K_���/�X�')�,��}�c��Ze6����H���qZ΃��O���8@RE���P{O�Y"�N�3OߙX�W�;��>�|�jh�0����ٮ���,��Zϊ'û�Qy�M����ߖg< �A��Y:l
o�b�.��EC�Bc��׏b�Q�A�-SI���4&0��?91¥����M8z'����ek[ý�%<��B6���������-��oP��aA:i�1��/�T~�z>E�#�,��zFg���͡΃Q�f�(�,�j�re��M�����B�Yi�������oޫ�o��8�����#�9X���V��n�d㕼�=�+��d�S1��@����,��Y��n�=����2�*�V��C�
r!j�˼�;NBq�g�PɡgGL�g8� �1=��tg͡��C޹��V�Z�u�뿡�H��&׷��Bȩ�[q?S����V�&V�|�8��0G��ə�E8��_�^���϶��F7,O��+��{�{����m,۵��܃T<��[��l{c�8�x�k����;5R������Ω6�
�����E��2X��	��-��l�5�86'�����%f#�\�_��y�R
�� �bM��X삺Lϔ�@��7X(Q=�s���|<A����ʹZ�7֩w��#T9�L!.D b��*���O�	��mN���HdYx<�%���� �`��\�,-F%���#����̿V�hP�6ߒ�V�@wLg⹗�,�����1�J�2f!JS{q��XD���K�7��;J����.��'Nas��W�Jfnu��wfG��qK��}-Y�h�s�=�=�������G�>;y2G�p��
��8��߄��X���~_�������Px��{��iR}��
�8���]�s���S��bsb�e�D���T2�%�5tL��U`n��qW����� �痮KX��h�&(�絖���Ծ��I�0HK��g]a��L�l���&&��e�4D����v�D���l�YI"`�F�"�4b��-����%��z�)����3_h��<�.���V@>1�C<(?gd������3"���rD/�lU�e10I-��e�9`�s���f�[���6-q�$3�s���9ٛ��z����f��d��Z��E2P� ����+�-i�����^�G����$�Ya����i<�W��![�k��������z�i�'rĳ�oA�;f]{��;:@�x�U��ڬ���Wqem�G���X����S�6�5��d�>-4T��҃�C^�nk�v���`���H�nD7?%� n�]W�N�?�l|Xx���<��y��hJ����U�YS�� ������?��a�S�m�B��L��W
�B+����������K�q�]�>���y�-�N�_o�'�>�Cu�0�R��]u����D/.4FZ��'l�v7�q>2�ʞ��ߥZ���3�R�S@����QT�|�)�P\Xu�X}�~��gN�l����ӝ�d�k�pD�%L}��~
f�IN7&7�`8�A7�Dx��f�]� w��T<m<����|�\p�����8 Ӆ���y|�	����	�1����$����vP'���*�殝̨��h��I�}>��]H�l��"~,6�/wtK��?���������'Q��H#[iҔ���w��#;��� ��Y���+ڳ-�fYۍ5����� [�q���m=^ǭq��l �Q�1�����X;p�F�J�:)����茤�*q���[_��#������n�J����V��3�Vo�cu�y�$G�t�RJO����P��]���X^D�~��k�&J��|U��m>��\APa*4� AG:+��p�Z�.+��Kz�"�啐ڢA��{�*��N��f�ߚ�����:�-mZ��_�7��u�1�F!��H�b�C��u��]����;�d��m7�I��T�����'�͈����Dh3���-8a��M��0������9�L)��Z��/�}d,ڇuƊO��#'aD�^�~��T��8am^�Y�B��V�D�^�@�1Er(BG��U��l��87��¢FL{R��W"�0����l�b�e�`��	t$����8�O+�yu+��Ed�yOY�Q�J~�"����G�)2�<���zϫ~f�s���>(`�g<�"׉|�q2�^x}�D!Q�p�N��X2Agm�I����s�4�B{����!A�A�6����ɤ.\�����#�x��+�B���Q��^����f�#e��3�W܆�_~�"���{���š?R>���&�핊d�)���ȫe�g�O��9���tv�/�W*�w%k�5�G.��y��{�M���w�U�XMc�U#s�?%�
�ꊶ˲PX���J-MpFW���>s��Sf5�9�� ����:�ax���������18r2R��O�*���a�@[�A��M�yp���`���AWP��k?�sq�:4�y�N��)��䛔"@�XJéXɼ�Y �j��MU>�+��F6�n�S�O���%ذ��zڕ!.�H�_�Q�ÚϞYM���R��髦eʖ�s)F9'a��'s��z�`�?[�)����eD�Nv�G=3Qfr���[�?7r-M�Iv�@��5 �}V�k�S~� �G��vmӖQ�4Vܹ��W�ǣ�~q�-0���~���D��',7�����Ox�5������N3������l<I��"�z���ݔU}����9n)MJ!��:���s��F��F�xοX#\8<w��m�w�?�gb��6�[��<����g}D.� ��yH4�9f�=3n8<O�Q��@ߝ�w����|�bISS�v�w���.�OE�,��K�8�h�C�MgUb<��rQns�/NGv+b���j�B��ր��ۣ
.��Mf7:����I��C���=Y��������Eyܶ��Bh6p��{x�v�H�T��#m�5�!<��DX���1�)�m�=�80;I�A=О���D�]��Y���D��r����1�;��̥��f��*˚=¤�4¼�A�N�2'�4��+�3;>�-0P��C��;Ax�Q����H��k�qPK���%�v-���?	
�La���W�fνl  fȉ�F�06?�O�@�?5SA	�o���7N�g��f�tz�뀁:a����6�=z�	ҝ�ԎJ!O �2��	M��ie���{�߀lr��u�Fid�_3��x�����R�vm��S�k�ε���K�f>'��W�Y���+�l���xg6P�q:��rM�A�z���7j���c�皨3�`��M:F���c�}>{.H$!,���<�6�Pj�@Q�,s����tp����Ӡ��P>$ڋ��  ���l^�H���-�L�Aވ���*���\��Y#� ����iM�h�%�,��YZ���yYO8ܸ8���$c����rb`�{@��Fj���؟�.�)�*�hNT3D��N�y@q@qҤO�G�i���X+OYn�*S��Z,����=�d��'6����@����B��g�*�u�s��_�-��ق1�dʸD��^q�SUTBXGh�:�A0h�H	��R�45]:?
��c�\�ؘ*9cY|�H\���8�z���I���W���45+-��ˌ^�D�]�R��{z��-�
VK���IG���>�ci�wN7�U��s5a��� (�;�U�3���jR�8� xu�<݈����I���:R�����8��XH*Qp&�҆X�����cQ�#�摛I<7Q,��C�An�m�kY	��54���9��[��p\|C�·ԉ�XL(.�ІUD�?��0��|���Z˰��&�8��E�Q�mgϜh��U��|��J��B���y)��x\)���R��5��L�g٪�@�%QI���!�1�i����z���+�o�<M�U�]��)f���x�Dik$d,�B�d〝H�8\PŞ���Me��^�b��+ ��2��P�.���F��O��-Ix��j1K�B<�gE�K-b�~e��N��?!t�G�Y�V7�)�cXH�N�Mhi����(�=�6�Ȭ*=��cC/�>�[����c�a�c"����W�+�xs{�=h��5F��>
�����ڷ7���HZ�Oo��d��5x�����)��[;"U�S�Ό>�r���a� W�����,�L<�0���'f��C����94�4�mݘH��Z1����	�H��m=kt|�)/���K�CI�[�^��O�(V8�H����9��3q0�"��Bc-*��Y6�s��r���b���^[9�����X�h����6*ȏ��>ՠw�Ӡ�Ώ0���I��To�l<D�DP@
#������,|̞[�!�R�$� :�_9i}����lح�h�oˮ�o?�I_S���z%�wP�*͆�&ܝ�P|��>�T��Ɉ���$��!�PD&�oTˈ{rz�h�~�`{[��]f&�~��4�����ksկ-qdyoq_*�)�']PN�a̴Y� L�RB%���:4��Q~���#26\�URd���������[�I-S,���fC���;3�Bq�����P�n�R����3�唤k s����+q\�o,�[7�eQ~՜/��|lR�0�){�}=���}��k�DaX��7���"�u���Z��M9�+]�n�ܤU�M�(�Q�F]YA���v�Q��1ηi92�B?.W0��ng,�����vc*S�<6�Z���a�3�Y��1s��zJ��\���H"�>��q)Ϣ�nS0��6��OE�G̎�\��b���껎�rC(��}.��0!zU�-[vi#���<K��Y�ӡ�L�jF�&��i�	b�\�V�vj��Tbx&p-S9�3��<���xπ�d���RG�D}UI��@��f���s���~fp�@���:��aI�u��͈N�G�&��y��O��2b3�R�(��8�%	@w&������!H�'ϸX6�ٌjW=��7g�x�`g�Z��P�w��;#+7��8Ƭ�=�p$x>/�?dP�B���6��6����//�+
7r��,%O����߬��q���蓘U'��L��)M�Ӈu6��ߚ�dT�ʄ�Vm�UV�C���C K��N��)��,\�N���X�l�6�7��GC��F����Y^n�\&A+r)���etuٛ��È���2��69Չ���j!�vW�'���ݧ�z�5K�nI�V�B!�OB�k�۴��;d���=�O:))�9��}���'A�`��M�&��m/�	$_iu����h�#}��Ȇ�����ѧ#&_�T@��i�I�ۡ/����D�%�Dw��>�gج��p���k��n�����@%&
s�T��cO{�f�Po��J;N�>����R�8�����]�N:_���C$�; Բ'�YS�!�^oTs>@-�c����!!Ioae�`�Ѕ�/-M!�:��'�r��;�lR�76$��{/-~De�պ��'*�Bǅ�r������w^�F7�Xd���wO��;u_��K8�l���Wf�+ѹ^h��pQ>�m�Ϧ�H�Έ�K�5����2����AW��	7��3_Z�s���k��ݛS/cx^�ޒ�Ok�Ir"���Z���8=��ي����&z����_?��t���~c>nR�l~G��Z���ќ�S�M%��8O�O����oXɈ�{9�XI���U�;��dݵ�L������&Ԫ�5�:�o�,v�u3����@�L�5�_�&�}�Z�	��Iל��{=sq�9���!��(5h_��5���@���0%�%x=���&�w�[����M�c�';�+�yj<E�[ی��UC������&�_�}˓i!w��4G8�"�<���J�ʮ�!�H�ꩇɰM�ԖF������q�fe�t�[6�fW�݊P-
�9�R���!���9b0�U��%Ч�u��Fr<�ꮾog�SA�%��g�����}ox]6�-S�1��̍Y�$$o!��3Q��&{w�ԃY���$?Y�!��� ����>ު�G�����U(�{���Ɂ�S�4��� ��,S|�9���'_��
�������kVϾV"F�L��,��H/��8��j�/>
��ah B�R�$��3���0ž��P��wŊd�3���-:��k�#�kE�#4I)�< �'0IHL��pGm?�GĘ5����j� G#�W��m��|���t����xN���C�o���
�'Y�0������>*y�f�T)��������hW9��o*�b/�D�8pS��n\~�ׂ�

rtҶN�,iR�� �<ʭ!�j'U��¶�Ш���DFÛ(���p���熲��k�̣�/:�m��7W�̩d��]F%����=��/��.WS0d��uĹe��/1[	��pR��2��������b�VV�ac?��>�ƴb�(�)��b��;���R�c�A8��+"3�*�)�x3��CD	c��w�̋�746�f�΅����ý�+�I�m�r\X�ߙC����eK�]3Z���t���6����Ў�/4g�^��r�!>�2��Ŏ���7�w��w�b= ���JHcH[$s���w�^��M`̢�Za�ȕ��a���;�sʜ�iS�6����1���u��3ADb ����J�v�y�A�W���5�LQٮ���-J�`�_�F3AoÈ��s!�����ybn�m�3�m��&�H��6զ*� .8>S{�~C�0���Q2�A=Q���_�ё��g�Q��A �/GJ�.z�EN�h�2!�Ϭ�!.FGp�x�@�n�Zjx�d��&��xߴ
!0��@��5���o�fŬ������F��0L�>����-�Y��,���J��O%C]*��^�lw|����,v5�`d�(k:J���q���