library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY LAB1PART4 is
PORT(
C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
HEX0: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
);
END ENTITY LAB1PART4;

ARCHITECTURE BEHAVIOURAL OF LAB1PART4 IS

BEGIN
PROCESS(C)
BEGIN
CASE C IS
WHEN "00"=>HEX0<="0100001";
WHEN "01"=>HEX0<="0000110";
WHEN "10"=>HEX0<="1111001";
WHEN "11"=>HEX0<="1111111";
WHEN OTHERS=>HEX0<=(OTHERS=>'1');
END CASE;
END PROCESS;
END BEHAVIOURAL;


