��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2��@l$�~�@C�.��Ep�\6�Ҡ�}�y&����9e�vK��3%D�a|8��ՊH��JA��_"5>�M7�[6j*�O���������;i�w�*7�@��]ᮢ�mHxn?��Z9)�`��h�4�
gƭzűW9���\�Ѕ�J�9ר�����k���8�{U*�it|?�:Ք��E�]i���A.j�?�&婏����H���:�C6	�Ow��<�BvE��*E`^~]m��x��
&�o\��������0����~
��4ځ�%�؂\f��/}���z���4$:v��F���J;Y0D^Z�\�b����r"���X��*m<l�Vje�-ԝ���X����j��w��cA�g*/���Vq���7��
,V���=�G�7�Ja��su>�u	�'�z]��,���"����C,A�&���n"��6�B��Ʀ��;�^�����Ioĥļ����M��+��'3��8ã}D��W�1/!�a�>M�m�)�����_���E�ND朢��)f6 �����0�����Jtf AV����:g�~N�k��R��H�b�:伣mί\����FJ��L�+�WN��飘㪓4��S��1��jQ y���f�����ҨJ�����$�p���Y����6#�Ր��ݦF�O�z���/�ݿ̘��윶�N%�+���7	���s�vV�,P����/FIL��{���F�������O��ءU^����U�\dٝS�m��	t�@䝳��ۛ�9�2�x��������c�p!�Y�r�Z~�˚����_��]�[�3F���n��D ����gk��D�7�T�U�a�v5\��	�n����`�H'�I�w�ꊎ%�Bϣ4n�븹nl�x�9i����d��k���r�蚂�IG��Kt�X^�
��[��	���9k����9�TQ��j���(�(d�d2B����E;���7E����2r�uM4�Ä��CH{Z�������*oK��t2~+?��S��2b�����������|���@�3���.�'�Uv��ْ�Q5�:����jD�5���e1���+&���䦰�\���8����;���7�]�ŧ!��[�Gv�&�v��j��\�2VA"I���X�g�4r����};y�aR=��l���ܮ����A��t ^ ��	; /V�@��{gX�P��*��}푅
��3����ǋ}����s��,V�z���=���Lˁ�wb5NՎ�W���ӌ�R�ߞ;wֹ�T${�k�os�U�:��[i���採������0����B����}�	��I�*SK�� ;+W�p�L��ىK�s/���n��X��3���
&.{�Qz�o����YD��\�#���Pp��R{e{t�m1�V�������Lȟx!e��^��8�u��ȇO����I�B��j=xq�Wȣ>�>����S��ܝ)�k@ a����E�糎��:�ȭ�v���Iq;y����+��ӽe��0o�9��aG���.]�9�2Yώ�m���	8����ax�$��y	����=�y��oH��f�6�P+����;�o���<����W��D[���Q��j�ؖ�g
2�m^D|K��m北��+��:}��E��N��������D%�b$F8�I)�8* �Ha��ߩ�s��h����{l��z)z#Ow11�ø6����n��'�fPTg�;��`���W�-����7����%�t�rܦ\7b�m��&�����t����C.����2���� ���������M�Y��&Z��8�B5�r��J��R9�԰�Բ�=pD��Dw֋�]=��IW�_���핓���1`�Bd���}��=����G��i��DǗ��ݝ��pm��'	�Q�0�c���}Ch��J'|�a����� ��|<x[�<���Y�b!*�#�B���|����l�,~��������:�o����-1��N	�F��[v���+�B�`ǚ-��H���{�Bͪ�A�� �x5��~�Hy=u��ӣ���fI��{e{�J1�E�P�h��u%�6I�vF������$l�HfY4yK���ubL~�P	�X#$�c���Q�~;Nz�ܨ'���?�$Ͻ%{�1�W�o�+5~�����4�ÝV�;c1A�>�����j�����#�n�C:��wl������L�E���f��:4s�xɉSrl/s0d(*����Z�ޑR0I򆂖AE�4k1,�IC̸��(kz�$d(Im)U�`MB�s=�A��"���t�&����(С�����!��2��5�W k!�ՙ�5�0>%V��3�p�h�m�����~�2C;u�K�ҭ{�7��chޑ�N�:Et���1i��[��N��-rnp�n����}HY�L�r�8��Q��hZ[�%�n��d��Re�6�
�{�ܙQ��,a��J���_7��$\���>��w����.8Bq����S-��xP	ä��]�8��Hw?\�֠^ÿ&��H;���m��j>�2b^ϛL�b*����Jln�c>a~�d7�&��!"��1���8�qr.܋������F�>�x����V�ދEŧ.8L�׽��q��"�Y��(�I8��>XMXF����ǋ����a7���;�>�>+�{EEk��5M1J�����Ҕ`�<�t��Q��F)�Iđ�<��3#F?>���1��C��/z6cB��;C�`��v���lEՔL|!�S�K)��"L�s�>G�e�KI�D=M��i����S��l粤����t��N/�t�<�;�G`滈`�����H��J��C�?jd3V��^&�t���8LӺ���6m�ck�Dq)�$?�����u���ܪ^g��_�T�^�[9c4�"�����BY��#����;�0��`���˳������a�����R�������qHgǩ����;�N��
&����NL��X�)�/'��t\)�M��.J���
;yZ����X�zs��%��=p��޽cKD��C4�B��-�S��i����4d�z��`��m�r���-� <C�y���um�Ǯ����H�p�1_6����N�,{��%C�w���ǂ�Op����_y-�����CЄI��h����C��DDjf��THj��1Tl>ʭ[��p�����	}� RKXB���pB�����ѹJ��9<y8������8MU��C5�\��Z�:�0F��#l��x�Wd���r��Z&��;�n� 
_�a���ءY�:���S"J�D������X������d�l�{ۅ�W�a��;�dg�iH˪�jI�2j��'ؗAv�n�<��8�i��������� ��i��,�c6.&���2Y��o���"!��`�?*x�7B!��=�'���=ծ��@Z��b��񳚍�备hbA42���y�d�}��U�Dv�t=��D�	���Ifw����#�ߙ}�\|U��%�����F8�d��n+X�_[��fp�Q��a���GRh���r�₌	����]��"fSf����s<�!{N\���H���@ћ%�\��<�8�/���)��C4%ߖҭ���8�.�S��>��V0F;.�Ev�B�w6�#�s7����;� �a�/S�UlR�Ѳ��lF�M�
�"��;�$�m~=�C�K��֖"v��rn�#i��.v/Tj���|Vy�o��n�Ԭ>ԏG/#��'T���|>
y�����E�v�@�#t�|��tT�/��*�V�(JYɴ�@��"�z��S�����o����c]��5�8 )�dg�G����jP��ѽ�#g�Y �� �%
�\0vx���09<Lܠ`N�p����p����������v�99Yzl� �/{y�~O5�0���vc)|30ZA~�T����:mk���|u��Z�>#U��e4�F��ۖ�zMrx�c�U��ixԍ%�kb%3อv ��w0�6��E��ܶ�\ ,���8.{1"""r1��bf4������3��-V,�L��X��Csi��}���}X��hf�|��gB�5�'����ca�,�Q/DQM'�k�j�i��.���S�RNĵו=>�N1��t���uo��P�ƣv���C�j��"��	$�!�6�F���ם{��/�BI��o_�����.��F&V���,2��[��<|�V���F����e_/ns�+�r���R����"\o�c{�\�b������#XX�O���k�A�G�����G*G��W�،?οX���31M.@;�γ�/ŷ-L��NW�����tů-�!�r%ZGR����q��%�j��B3���*Jڂ٫�����Q �+�j�K�ؽwY������h��Wj�'d&tק`1nĊnǺq$c[�$�_#��$~7j1>Țyj�{`�Qv4[���d�o��tmw(��,o�9}"B�^l�e<@+���"��ǰ��EE��iQ<"UE�zBe0n���Y'%�Y:�w���.e���"����5� ��R�����J�Qb����y�6sVJV���T�h����� �ՠ͍��t�(�;���ߩHeϰ;s��@�F|� ��0���^��`�ȮX�a���������yڍ�TlL�BO�?�(E���w
r�'q���5���D�
�@�-:�V$�H]s��O��j�q�ⶤ*j؊�[��ܘW���.4b�b���/��-���7C:\�u�9�{��$�u�BQv>����T� ���vb6 �ϒ/�x}v�C�;N�L/ju�\��Y=f`=F��2�`|a����f�J7�a:��+m��]X�k DF̉?�i:0)����г�8|K3�Y��S���!��N��W�i�C`�/[Bn��\���1�-��y1'3�P���q#�7Hq�Ģ���;��=��k�����5� ��%ް���)F#%Ą�D-q�SVP
��V�r�@�Q�!�n��Y 1"�aB�u�}���g��A�V�8���G����݋�&�lat���XV�Ƨ�v�8�:D�<�"{�3<�[TF�Q���傼�7�s�rY<A1���Yj�V�����p����S�_ũ�ߡ*�:�R��;�Ʌ�D$����D�f��a�<�1ˤ�b��M��H�%��|(����rՐE���u'/ �6a�p�fƜ�G��L�a��6Z;J.��A3rO{�٧�n��{��(+NA�s]#RH��RwD+�02:r�E��uW�\8֪�<?!��=�0U���}��-��k��c�t����X��_�xd��-�ԅ$�]��E������
�N���!o��zg�h����K3Ϥ�B������sm⚡�q �;ރ�T«LhRzD�TiHUﻋ�W�歽�2����!!�K{K)P��܅��VgT��m������+.���c��vf��B+��Rґ~��]y�,�r����VE��(�6Q�5�o6I\'����I|i�tglJ�k�4�����U���V�<
:����(���E$��� �{���r���GF�x���nI��l� �N8�}���w��:Zh��zC��%�^}�`ai��e���$�$��ꀳ
���0��:��V���wN���є�=��l�썐�L����C ��)���3�H��ݼ�4���\鮘8ޣ�:��J�C���
��٬���c]#��}[_@�>� +��Iu�x_%�ϬR�l�u:�F;�Z����AF0�Rf�>X�♕Bo��%������WV�����$�7V��&�b<D�ߋH�B�~�)��X�/�R��Q~��ۅ"Oh�~7:� !��I0[��@�,H�j�={^�&4 �՗	'�_چ"�y�ئ���h{�7ߡq�}�˗8�_dl��j��A���9/�&��sb�7��r��mJ#���0_ԅH�����{gdi�}��0�� X�����0�/z��%�C��@��$a��)B�����J'�5y���XF',F^@���<��-}W���sx�ό��#�o��N'~,���L��`�p�e����hC��h�������eg��B[�2j�SC��$��6d(��i-X��0�u��K�$���Ի'u����G��A򾟈G�h�&`X̸0�n���n
��)��&?�T'��qI�ؓ+��,��4T��N(�k{��g���6�S���	���p��RK����^J�K���wU6�-#�V�"��|�"�|}��Q�X�4���o$i���i��ݻ�g�{����օn�,��Sv����Eie}O���%��E�(�q�2#CS��{��_�#ȋ��.�f���� ż�(�����B�[��RI���ABU5������zb���u����l��I�0P=*_�<�Q�<W�e�:��;�+��]V����;F#�T}5�3�@��f��=Q�^|�kP��=E�0��IF���B�IYAT�D=0��V�
���æ`���,č��K�3w.��3ыZ|���A�w�(�M�?���1�.�}�F6�be7����
V� [u5OAB����8��?�\�{E}y]?���@�H0L�E��CK	������6F��"�=����ᧉ��S̟g������\���`�,.7S����1"5A��3!�UFƑc�-Fk<��A�cfKhT z��L��9��Fy�[P�ˮ@�eI(�t��A���{�a�j��9Ű�K�ߏ�o���S̿�3ز�ރ]x3�^삼��/8&=2��H`-
��S��|6��~��4{�Տ��.��O�P�H��)��T��򜷌1{�>]G�/7r��؆e�G�j,*���Ե�������=g��Y����B�����������	���`w�,h���jgv-���l��~�b7�}�T��b(�cZT�	~�K�����)���J�Ը���/�8��:�p�R�~�~�+j[���4�2�l�J�Rzu}M�/<����u��*,4�}h���;]*D���{[�Xʼ�&��^M�U��'ԟ��3�Đl� �W �{��<�2�ە�@���e�����PR�~�����X�J.X;�p�EL�C\Z�]~X��;`�D:6������.ƔRD*\9�t��t7�Fs?��4��7��J��b�h&.!z��8C�E�r/��ͬôP�FZ`���%��:�/5���0��z����4,zL�w�e���2�f���aIK���\ܗ$�XnjDd��o���8b���[����Y"'׻oY~�C�
+��s�~\�2-�0�����8��RW����`��/{ f��)N���V�O����l|+�`UM��Z�/��֖��P@�[��J2}�NC����"��މ���rkv��XE�V�w�П��6�B�A}�� �`��ur�PP;<휫ݣ�s�E��� � u�ku�vL;V�e�]���[�����R�g�� �sɔ�E����Οm7_�è�  �r�iJ��<"��H=�^�Œp9?�Ԗ���/[��v(w�6�0����
����U�GA�G㕤\��Eʥ�y\���L�o�O4'�UK!����O)��%�Z;k+�������T�����.�B�����c���M�l(q��y�rl��������#s�#ddDB��]�9rϣ�#8H�,a3�y�z�]�Z��-�%*�/�`><��)�m�N���l���	�Ή����b ��� yK�09s��䬦u7�W���<n����շ{+ݕ_:B���~{� ��$������/ml�41P�U���|��� 2v�Y�N�a�:v"v@�ݸ?T"-���^�X
_��
Շaǌ��%PzU�cq���@�i{ѧ�YM��0t�,����iۂŠ����LRچ�3��Y�#O��gq^����_5�9S5��8��z�N��O��A&�D�;1b��u�c�+0��� 1���_���c�P�A���+�ygJ���y͌���7	�!hM�ݹ�;	�ׅ���n�y��M��5�JzK��JF�@�t�������VΡ��C��Ý�SM�SXV9�������a�i�`�����F��[s����ը:�Gi��~;�}�ҿ�7��|�_�*��Ń9����^��D���Yl��(�l���%Ы)aHZR�Y	��M�dNɌ���o�͎ӳ��ķ�Uoio���>�x�V���\5C��I��.ZN��+�����qPMG��86*��@���E3��,�!<�zb5Ni��O񸹰��.ʠ�	��T��	��3%n��C\uO�I��Žۣ��~zomy:҃��UI	��g�,����%��g;띈��ĳ����gj-��X�X�g}'���S9�	���w5K�EͿ�'��э��Sb�-��]�@{������$:�B��ɚV�/0��N*�[]�E�G��|���-@��)��C(Hng�yeLA�
Ｉ��ܚ�l�'��l�����K�5�m�xbm��jKif���@�oﻨ_�ۣ! �v�}|J��0=e��$Xͯ����@S!.����_Ze���ѝ7qǘ'���0�oL�қ��l�,a��� +���0T�j�M��.��{;S&����f"���?fKB�-��2��8܂J2�@��Y0b���
�$��$�ZY`m���Bf|�W�t����蝄�j"s��U��� ���g~�b�C�٢F�'�gV������)rA��^3��v$0u��hM�f��FwC@�
�i5�JY]�S!���[��qcX;�%c���*�ش�O>��:�UuɼR����s�!���!L�+���իm��|1�G6r�J�����'h�!f���I��FM�S���0۩Dj0E�5F.�g��y)�eM�if�ݖ��~��5���j'RB����*�ో�?23�*�� ��H���K�zD%�ϼT#s2:L��f�s��@���pl���\X���?.ט'��i,'�F�ߕZ���.�Iw|d߄��cW��pa�7S�Y�)�
2xC��Y2'�x�r����6,{*եl��6�	e����Q���fTGs�TH&u��?�V�f�@���G��=���V�;@>�sz�)l�2�f��M�zy��2��.�C�;�q5kJ|���(E�ÿ+Ʃ2O{Ű�����u�Z{|��LE]�V�a�rBQ3��|�!��d��ҶM�$�T몞7�6�jreN�^�+��9T��-��gV2\��-�Y�;ہ琉3ʍ�/ �ڌ���4��^�QX�t/2��L��1����鬞D���l�F�)��1�>���,q��*�O���%4Y�!�Yf��0qh>v�Y��|w+�ęߜ���Nlw.'!<����p
lp�u v���Rl�����YvY*�����r^ c]o���������t�KZ�͡�'f���y�>ux�95(h���A�8�y�=Yŭ�R���$�8� #�k�v�v��[}��u���ُ�r]�^����m���5�OXpk̽���BoP��*Î�բe�p�����	�2C4���B��\h!ȍ%_�$�ݡ���Q��Li��r�����7j$�y��N�b��[f�;u�����g��y�-90%�!�qc�R��BX0Ҝ }a>�#�	c��b��z9s���}���6þ�'m���WԈֻ|�2^�pG�
��.���*Q����Ø�hJu��_V#RO/��%�+�ޙ烕sQ����1r���/4i{�6�j��.y`LrWX�?��P3F�H~�i9S�Zo-D�* H��n��ˉ�������<5ޘ�W���8f�ǎˤ���UȥZ��)��wdv����e�'n���4��8k�������YT�0M E�E/�q�š���b1�|r=z�E�^ ���Z����Zf�%�ȑH]P/�fM��{���.^�F�c��J�Q���s$�RR������/�}� ?�T�Ŝ22�Ɉ.8���=^s�I@���e�enp|ߴ|x�h0����?�+�&���XÕ��=�1�S���f��7%E������
��菏 �Ï)����m��G�J��!��;$$Qg%Ɯ`s!��l/����"��R�����2
d���~B*_�%��.�{����}���j�wh�>T�-�d� ��^hu�$�I��w��Y������X$��A�s^���U�[>Q����_8K�f�{{|�;a|vc\�����Z$�g��[��oB>�*/W[O�q��9�JU�?���yiAS�k�L�ѿܛ�1�wT4�G]��y��"X�{�r�g*$N���:�!3�&=ىVmܟj%�*��(��N��M��;a�Xq맽�[c��@��K6㧏�a��~���o�j�/*�� ��.$����+����$���^W���^��&8��:�7�0��o��\~��͗��|vR��;��D���˺�'�ə%}vg�av�>[�"����^t���?r���řu���8z��P������Oͥ����Q*�z�h4Y�M�j�����!P��� E|}:��M3�B���̗'?�L��'Ǿ,Ǒ ����޳6�A��G�čnG��1�Ĥ� d��j��)��u9Y�l�J���-���f��k֍�;��o�!kaP�O�$W_@T�����k�_��`�[����|�ĭ6��6�K1���'����v���V��P��En������Ga��>�`�U-���em�T�/W�b�����\k�',��܄L��M^�,�l-]��໘� ��H4xv����E���Grc+����=��U�3V����:/Pee�Q�7E!ޙy��P^J��v}�7�|�ӛ��h��j��s�S��ǱK!��\R���M��[�s�I���P��#��G��|$�'?9��M���t�Al�}?=R��'�Vm7vE ϳu�����S��9��OY��������E�Ï��o�U��M�<*Q����B?�95-?r�Ġ�n�6�ɋ������SX��gZ�W)��� =&]:��xY��h:;�pRX���s��̂qD3x�x߷�����B�kl�d����Ա�.��Q��m��M'�.�	�*�/�L�:X�Y�/�EZ��#m�N�k��sO�T�{|��e}-4L#����,;`�ݿ���$���L��Uĕ���Tg_���_��h:�P�=�f.Q�#���s�D��x������}��̀�o�G�!᭠�nd�D �h]��|�}�`�+�����n}b}!��Y�z�֯�
8�Ծ+��Б��S��E,k�Z�Ǳ=��+zh����}?KՕ6p����ۢ��~��Id�sp(_��[�efhx��Yߝ������O\$����������A���.Qx������<8�h`̒բ��9�����&���ꮹ���ByJ%����a�w}/�H
��߶�x �Ib�.I����C+s��� �S<��G�\�dX�^J]�<��W�nb����'7{��LR�:!V��i�x�y���ߑuF�U��֝�*�õ=,��J�M��4b�xD/�\p��^n*! �ۖ4��e*��V�t��@t�#���9�f�YK �����ݝ�9�2��^�B���3+�ŕ�rݶUԉGbBj��l���.��n��e�G�c
.�6z�ǇY�����9t��5�@MS�G'W��smK�5�]R��6z�FV�8�'e6j���JRK��E6�В
-� ���f�Ӽ:J���}Q$a�9��~FN{Ӱ���J:�P�(M���&�^2QA��z��UƼ暙J��w;�&Ȝ^r�Pw���*����cr�XsDT`��b��f,-z���F��e��WT�=���M7h�ڰA]O]��B�+X��뿿pI"m�Mm���s��+�x�®�3-q7˕�C1l�p:X�@j��{o���F��S��t<6�������0?d�Y=�S��"c���C(�WT�«��s���F�|��r̘\B�#��1_�c�a"я.T���0�l��iRY�.���Y
 p��+f���p zuWa����01o/�(�f�������L%��|!����=������DQ��j4ר�P �VCGw0��s�3�]���`���`�ٙ^J�WUFO��h��.���,�6���5�'�|�MZ���(�|�������`�X�G;�>�ڑ&k$�J��A`��9;�+��[����t<�q=�M�{:��g�g��t@�5²�F�!����4�$��A��(�h�0����7]Ҵ�y{z��`2|�+ͪ�S)s�K�/���$(`rߍ�u	������b�8����zߊGDZ���B.$�P�%����� >�Ț�'�H�*�/��ɟ��j���|-�	�[#8s��Խ�iJ�0�d��Yl#]�o�mb���K+s�
���:,8�_�_JueFU�n��ݘ=eE�[�T8r6�9�����A������?�0�Eh���B�R�28�uw<V��D:�C�;� P�!ӎ �o��m��;�����MF���HG��-�����K���!�^u6�p��#W6l,w;MO�SHnL7Um����|�At۷�'����y-�v�"�:�w��$�Z^���C@�ݼ��2!ϱ��<�{K^�o����6�wo���*&��MPoj�lF=)��L%Q�p1����W��}hM�a��{�4��ID�����FA��NM���R�\�_1g_{wI�
��e
i`�"�;��!�Ff�qHmȝw�d,�`x�y���q>�rFc��F?����A��ŀ�bjܔ��0���=_*N�����H<��ںl�s����&qI�w�V�@�[�o�̈�d�C���F/��.%17Q�z���!��}Y�Q���*≨]s���Үy��5&��s5Q�5�j���J"~DI֭�7SnI�C�c"�Χx%�L�9�^e�#eZ�)o�Igp�(�֨�X�#�)=s-�^Y;����/�՘U����l�e#:T�����u��:F�����z��5G�����B�rF�V��,����.�f����� #b`�����)�Q���҄:�U�� �G�g��x )��<w#��X�N�������D77����P�bL`^Ng�%a~6�����g��qL�#����
��Pz���y�e��g��4�ISj��B
���A>��ɿD�� P�P��v�(O(�|XHw�O)�^Pè�i���ëȇ~N�PVƓb|j��@��ɢ�����������L1�P���9��e��Pr�j����w?�K_�`��3�g:��zzו�RW��u�J8۝��\�>l�S׻�/$���D�ZgoI�g�o�&t β�	���"���u�6��3\G�Ő!�8�$�x/�דjMt�{vb?���!+�8��"V �� c�������M3�yj��Q�IFLt2��������4Q�v��QD��O��p����3���6	���fXk0i �B��tuNn��N�&����I��&@�蚆�G��nM�u� �I�u��U�FjL;�yK��4.q��-H�F���2|ܩ?�ip���ƠHjRH�>���n����w�Ԍ�,o��KaՐ���7	���ﾶ�o4U�W�e3|�<��������4��Y�y�����'��4�����T8�M�S�R���|WwX0��7�������%t�&u�|4�^Z1����D�M�5�l=�'A�aq�8[X>�l������ҸذF4P�!W%��C@�7k�����D�f^nDhȢ��%EMȬ���񥶡̼_�?QϠs�W}S��\@�R�~�ģ6��*�&��L�u������w<tA�ґ�� ܧ�+��+�6��Ή?��VO��!J
{i�D���+���Z�с�x�������A�u�}���,����;V	_���[$�����E��Wϱ�}�,�Mj}��Lj��0���<��M�O�4���K,��$���鷔#dF��S��>'9�d�"��~<eSG������N����lا���I�n��4��O>�`��i�����z\>l��!�c�-t=�FS �Ò_�Q��TNIj�Y�ô/�,�>�5���f(��(�+�1�G�����*g=z�Ԉ�UA���j�7w�F&GL^U������,b����/��x�Z���#;��ެ���d�����8[�r��A�pb�ƍ�?��SF9�	U:�3����j)[x��ۀ�PR�|��v��	��e��=�&u˦���Rט�et����
f����`]��*\�S�i
WN+�i>zz u4��Q��:.� M��`��ͤ�n^���iP�?8X8��Gˏ-jwm̂N�_�@[���Y����f��ʺ�Cg^��2`m��5���ϐό�3�^&��=(����6^��Z�J{�I���~����;4�0w#��9��H�����E9�< �<�Ȼ�*�@:����c<��&�A����^��6%�x��c���+�dぐ�͞(�1s�_UQ������'qVBm���sOl�(p ^@6t��g#�D@��&7�j�s�	E(ш:�t9X5�M@x�ў�*G�����ڔ���]8� �GKY_}!G��5�Ǒ��?2#o�ˎ�	U'gL7gQ���ؗt�/��[*g�ڹ��r]H�n���t@;-��(��2�u[L�����ۤ� �A�x�w�,��ե�js��g�!����b���u$\���*R�
@��Dt�9M"��^��Tɗ����(͌H��x��zm#	���o ZB��p��ҍ�n��,�'�6���P��IuH2��	���Wdߒ}&9�.N��c9�ZuH����U������8y,�R��F��^xA�IN�m�-	`F��	�n�.(��o���m�C�+ye���M�H�vöқ�@p1�G��>�����
�*=_ٯt���4zh:	�r�|��8|����2�:�!Ңk�U��o������m=��R�g�׮��c�*ގ[���,�y�6}���	���Cx5t�\&$-��t@` 0�����Y�okX�É�c< �)���������0�AR���z��u�P���Ĳ���;ǘ��5U��b�K����`U�#T�ZGv��o�e����g�
�[J�,�.��G5�zX]щ�DX�o����*$��<0�+ܩ��[�KM�	9�$�.��ŧ9L9���T�!����8_�30��n��\<V���t�&��8�m��`��Z�����lcr/( �c�:�B�j|(���?�
�	2 �Ӥ`�m�.��W���&��O���i�ܻU&QP���jh(��O�( �=�E ��:�P�լ��1�S�ʻձ��7��x���;��R�~!|���R9ܼ�Z2���Wd�l�����Uz�a��\o+��)�c^'|�1���Ÿv��0������NiY�*XpO0��Z�#.����~v��`Q3�m�жS��$�	�-k������ �cBc�ϏI��zT@�B�8�����}����q@��Ls�)J���]�U� ���=�[��Yo�gj�q��j�����or����>J7RY���7P䶴�fwA��[��ץy�N�v}��le#N��;�v���`��b3ۊ�}*���i�`�'�!L�@N�!r��K���OU�p�x?��t�r��a����$ �)Uթh �C\�B��k�F?�m�>>\{����a������
�gЛ&8��3�e�~YD4�1g9�c�yP��`q92���E�碒3	T��2\��m]���<l�RW~�e��a�F"^S1� �+K;��lP^�=��Z �ۭ$�W&�:e�-�/���\���OH_����r��2��S���+�2�`Ц�zY��$` 9�[�%�eeA��Zr9q_�m!e�m�g�d��6��(D�\�Yn�����`��qu�Dn֢�!gP�w�=CLj-�!��C��w�68}ؒ1o�؛����$�_6P	���j-R<�ɯ���<Wگ���8�H�e��VZYc�x���n���m|{/�]s|�oH�\?��r�s*wX}hS�Յ�Q�&E��C6�א�᩺�xg3���h�Z"Na�:@�s�`t;���6���1~m�g�?�wa�p��!��#DA��r��c�,�*bG�v�@W#�0�6��<5��/x�����`��j'��3;xi!����"K���|������a�zA���i8^�i�Ç{��:��Z�����ҳ���R�pY��ʤ���l��]x:f���D�g9������w�m۠����_��s��l�t&��L,ǆ��1㤔��!�����2Ri�*�@��V��XX^v�u�E��������уM$p�|vk4���@�4����H���*�B�VŅxcրl0"�^�E�X�FBoUB8  2\�Nȹ�u�1U"a͗$!���\�\�����W�n��4	��A\��i��
�#p-�V��o�/Vo�Of`���G6�L��5�bMEF��%���-�T�" 0�\��%�5�
��������Ճ$Y�Au�&#�B�z%CD�:ىh+H��[�88�#���#0��- �/3��E��tG��������Z���⛙�������ޙk
Ҽ�>��A>x%�-\_�����n՛��:4Y줋��N��8��E���t=ˠ"�9q%��|��6���-J�B��<HG��1-���pWU"��}��(7���
smg������Z�<>��k+���w�EHc�f����	�k�Ɓ\}�2p��M�r������[E��~��{�u�̾?g��7��G��ո]�f�����eK�\���5�#�+��:�q�WÝ�dQC@��@\{�'��Wp���;-#\����1
8;۠n��3����
��,ŃN��;:�CA���P��u�O�b����b�h�C�f풵���F�څ�F}zhZ�e�/����oM
e��P��� �L��Nt-�	���_!��D�\bg�r7^���"p!�S�&H�k��-�b��)� by�x=�u ���j��V�[z��?���=��B?z{�M���,�>9�E�.X�z�~g���QV��>{F����ңcU�C�_���W��A�R�h>��X��S���T&�h(H/˼�T�����e�a������]���2^���^�Sp�w���`��1	��[S�8z��n���A!�h�A���P >�oF}:,� 1~-��,H�����T�5�_K���|�c+�����zq�-��n���
ִf����»E8��T�-=�Ir��L9���a����T�af_�Й$�w᜵���]�.A_�D�[�vrM�=S�)����^���!\Fy�;Bv�<�����7�qGߨ�"�Or��T�.�slx�u�O��EjY[L�=��zl�1��7V>�g����D4�Nt�"�i��X��:�����9����<�I��c�<0S���Xgp`����!'rI���i+��ȏ��f�nq�|ջ⠁�I�χm�c�V#FW�.��=��{�J���U���:gCȖA��o���n�\�)�h3��i}u���#%�[�k�]M�Izy�B�^4�h�9�t�+`EZk�ѽ�@�%mj����|91��6�N5�'ѴC��RPA�T�����4ר_�,����U0[�@;��|�'Sٚ���#�֢j�	Y�˜[|��Z��M����n+�Q�t��t���6�F�R���h)��̩��:���g��3xM�6��WK}�p�7�>3ق�@�x��K���d.��(w�I�f  ����t�8�i�=7n��Vl75�2�\U����̈�h�E�(1/鳵&�(>�Q�ۤ�k��KZW��9rWZ@�ΨVu$��j6D�]0���h��h��hـ����D��iBA�;?�u�<�)�0�[�0��UVLz8ݐ,�ѕ�8��Y�ʢ�@�+��kB�x�!R�$��w}���mMU��2�Ӯ����C`�E�xQ���ۚ���W�cY�d}T�Zc=�U.���]	;v�"za{v��:��~(|L�C_��X��(Go��"J����I�z[D���y���=M�GQ�����7Q�WB)%J�;����܄D� 	LX�͏�l�>�_��q�t; �F<�X��o���3t�E:��oW�sť���(y�؇���ESp���{����C+rS{k��3�-�K`Ԅ�A���j��	��>�k�l=T��:���N��a��K��Z�i�����M+�����m���KL����YR����׺d�M��RJs(C��}���tP[y��4mh1Y�L�����]�ϖؓ�E��>~�ͽV�f�M�#�ޖJ߇[��w�փm�E2��m��"���u��n+���ꆢ$�`?ʯ|m�t5����כQ��Ƶ��J%�@�w�;��Qㇷ��/h"�������*��#�&�+l8;q�X*A0h�ΩV NȆ��9�_g����<|$64h~R����l�S��S��OӁ�t/�΃�iy��*T3�r�Z�j[��g�N��lX%iH�o�ї;N���X�����kv�&��Ո��m�w��kX�����s�1��{"�bd����q�k�ge�U�]|�a=��f1{�48���t�e)��9=����[$1�0�~XFc���H}����"���Wb��5���<�/�[ޅ�o=�"D�ʵ���pj������7U��nr*��*h���MqS?v�O �y���@�Y�}{�qS���(��$�a�����Gw1����T)` o�g;6�F���72`�"��� ���r��C{��᠁��8\Jm��}���&?0��\ �u�����|8���Ai�V�y�X�$�R 8�_cg�Y�x�ːEy�dc�#u���kq<��K5J,��t��\����^�Α�:�rA�䃵dPzzO�H:}�`[zә��pYO�n��	E~+�6p���w�
q�1�Qs�&t@�0�;D�	�6�1;���u�<�i�p��@x>'�O��S
p����
s�R�١�Ek4���~6�:E��jsC^��ߐ0�'�Ƙ�/�a�HE��Xlۀ<J��0d��� ����ѐ����ݢ���f5.���E]���X��J��*<.��S�u�A|&��;��:�(�$�4,�K���F��.n��;Ɩ>�s���5�p#�V��m��3h��۝⁸G�1*����6Y�(C 5�샱�ug�_�%j�	CH؀~�Z竳\��x��3�j���О�8���������H�Ɇ��M.U㳕��[*"��zd`��8�97r~�#{=��)��#Pq�D�nŴ�~<d.��}�*�N)���oy�G�&lIVs�B�$=����n,
�5N�9eČ՝OC�@Ը��>z��^��ܛpȯq8���',�~B@!�=�L�oMWin-Q�qOAǈM�jH�@��2gұ�����Tن���2����D����%��J��Ge�W�mŸ����|7�`�h��$�Eg�ȥ5�{�#�Y׉��Z�1��n6����,�}�1]ju,�F~�<-9>���X���A�^�JV�8��yPf����8I�̻�Pg�C1�Pa��6�󏳠k�^/O낝ٻI��(��1V��~%���SK�P��˾��Q#�oڂrh��Br��Ӽ��� W�����s��)k����@�o�G�8�^�>�9)��W�$��&�}<��G邳B4*^���1Ѣi��!ԭ��լ�������k]f#�"W�Vh |�Hp����$���9{7�C,v�EO��G�KuL>)�xBq��q:�rb�����F����ݳ�:� w#@'��o�Λ�.�Y9#��m,l(���s��J���Xz��#�Cn��Gy���e�I1⇑��K�/����4vw�f�T2˿1Y�τ�䁸bh���4;��*��%�`�%���
�r����ZКgy��}���e���g���z���Չ�6C$��䎊)�a��|�J�у�o	��a�w &�0\��?oeN0�)��VH���pP���&;����ˊ�N.D��@7�9�<1%V��q^D׀��~I3�a��=�B����3 ��"{g��|�7[����#��5�,���"΀r�{g�H������.�5^�xRtQo!��H�� ���xôH�ȷj�8mze��X�}��2I~[G�@����?g��Z��$.W�	�BS	���Wݿ'�v��ιʒ152���/"�,�M.�c#��G~�z�"�z�FH:L3Hw�TA�0;,��j����U	����w+�#��#������)���'I,Tc^�}LR�Z�$��kO�%�`�/a�
r�7�,3Y�����UG�P�h�{�iS���&��aQ�P��\^�������,�C������;jBH��_\u�^������N�m��嬨��l's��
f揇����G�j@�*��oN�m��_j]�P�쇅Z+C]'N��nlZ-"�N��c������zQ�(	�V�S7�'�aCY��N�ڱ
��dֱ��'\п�\���r͉��=�Y�/�"u�<��5�� ��봭�B���	ҩG��ܮ��~�?��!�KT�c�A#nT,�W���慼::��G��QM�">s�������
�py����Q�Z�3I�b؊ThcTF][R���7E����c��n�[�Y�@�����Wr�8E��������&u�z��j�d�8N���#&�9�m#�+c�Ե���h;�:�b�o6���ɽ�Z$���}��
X˄���QF�,��`C�Y��G�o��iV���i���p>Og[���^����d���)/��(3nr�J�)��I�J�F2�E��t��a��8=w����.�':�J�L���K1����Q;��3/_�(^t��<tZ�uwg|�DAڲ��{͡�D����jǦ�Y��7_Y8�Ky���!���Qh[}L�
"�b��e!�y $����F�Bc5:��wN
�c���D@5�J*��{�hZ�����(9�r�zm5ӂ֌wp��Ik����^��x�歭��
���ɸ���*׍���QlD03�}���߾e+��
�ڣ��-fP0���c K^`���L6ǡ���h����S�[�'nG��斜��N�e^��'��ɞD/舮H��V]�y���j�WJ�����H_׍I�cr��I� ��, �+��IO��t��k^.F�nҬ�8��FD�x����ު�8o X������IW�������=�,)�4�B�K�����Z��JG"��M�.b*�;�Č>�e13Y(.�����V~��j�c|X�D�8L���M�4|�|A������7��9^yȮ�e�_d���A�� ۋ��3���ꐓGl�����.����+��6��If�� ��`�y �؈�k�EL�,��Β=5��'Vnsq8�f��~���y���[�L�Y]h*��W,�%�:����8��Դ&��N6�\��P\�	���{s�C�]�!�Iq�B�3��XU�w?p5>*�m�*�`� ���*Sy9=����V�Kxr����F
H��$P3X#T 9�S��!�
ݘA��J�C���FW�Z��gϊI��b6(@o�f�!pU�	l*ݬ��0ǅW���J/)ו�����B¦� o?�bذ�ͣ���*F����7�o���39�4��F����~��s������ j�qdK�8ψd��(.�g�Ĵ8���� ����	�l�b�aeцD�.�K֡����;���&%���Y���n,.�@�Oϝ��((7���<���КE4��M���ƴ����ig*%4ӧ+�J�)�/�-��E;��0����/MǙ��O��`�msB��r��Uk��ju\�G�mY�����q��UQ��@��!�4�/BѪ�����r�?,aojx��z&a��g�!�#��t����уI�Y��M=��c��;���H���x�#hFZ�t[NG�4���F:�RR[��r0�a𵦖�5{��Bj��m�R�k�Jd�TNva��By _���-��Y��&�E�{�l_���\x*�X�HͮR+��M�����?�8(M~.ȇ��a���A�s�|Qu�%�q�kEm��3��~O�1Q�&NK�^m��XC���_�'I )
�K�]��Dm�Y�]�:1W�d%D�_��=�繛(�y�hm�~���Rg�������[�r�,���Kd�� �J���~p�S�D� �������a�����7����:�-KKt��B���N�5�S��Ԕ��0)��S(�DB�}�]�o>�'�!4Lo��Jch,9�ؤ�Z��z�t޷�=asMN���Ƈ���r��Aor��^@pV��g�
�Af�Q[߹n����/B���b��I�uR� �������?�R7΄#��b&m�(�F��E��!+�}�*���{J��\�`N��}�'(��5;��)���o̅Q���������5�:F�V�(�-?��pSK	����=�N����·Y�2�[������l�������T�d��p�J&ey����ꥱ`�
E׹����wX�lR��`�jdc��Lw<	���/����8�T�?���#�<l���b��p5�������Iw*ʇ��d�s�K#��Rs�k	�fM|G0�Ú��G�AxE%>Δa)@ � �m+�L;�U�b�O�-�����EYXk��*RNp�u�oy��t6��p��q�Y.U�s\(3�eu��r�h���� J��P3O@xm��쥔[�2�����@�̛`Ӈ~R�J[Jsn�A�Ш.���.��������/E*c���}��ۣ��a�;x���θ�_�?��a���܈����<�TW7�W���M�����'�݌�a"9ϗ�����@��"�Ǖf�����X˂�	��.���zoA���/�0T�S(_:5�k���Q���X�=H��aI���O���*'qA�����-�*�(�6ה7��@'�)I7�e���t�q���[)�7F���|�mk
!�ڷ�ˎ��O��Q�	j\�<8S�� �lܗ6F-|�U!n0'���釈	)Vݫ�T����Y�Vh�l��x�9M,7��)���^%H4�w�U����_�DT��v�������>`�Z���AIAhx{6�ʙ`��45n��Q��t�[�#2~���ߑU�ژ� V�zI��l����7T�k��0�ک��y�E��1ХXyJ\��H���xOtu���P�")���G))s�Ag��BMՊ��pl-�O��ɑ�L�E�:��3'��%o8u#l8C���Y*�:B�ۢ:Y�|ŋ���f�
�F8,�O\$�I���F=5�����J�7�#H��=A�G�Dg�\8�odb1I���v�G/ZS.o���t��瓉�+��n~d���!��.�#7J_�QoS#G�5۷�O'�7̶L0<!������&�W?����'��32?��q��	�3Ƌ̘��.6KS��=����6��h�z�g.#S�f��
�TD���4�@��{ ��f�M'�x��:���ϸ��R��ģ�J�)�d�[�aٹa�;��[3�+ĵ��hR���Q6����e���1hs�^_���C?����'�,6>D/ۑ��<T���\b�
N0ؖA���H��^/p,!R�/�y'g3Rz���i�Q���
�v�qr��_�\�s-��_��S��Ш-"%�CZ�UioU�U���tT���C��"��a)�h�^��!�\�G��^bx55)iфk/��JL~���X\�pS4��"1�P)ƸR4���@�F8/�^_�N|@�2�U�Z�HO<{ʫ����E�����6̦֗o �n��J�*��'Yn�q�~1t����[�d�-7D�U�#���rzh-��L�<�<�e��3�����8�_�y4��:�K��}�I�d��c�%���"����ś3�O�+�7c(.�w�����4\-���c��ޅ~[��d���b�����D�'&�*\�v1h�t{���Q��B��:F�Ώ��z|���0�K&D�ʠ�:���e��朡 �����hnkr[m{�{�z�zV�^�Chj�cm+�������ii�َ����{��Ϙ�g��W�:���H�����w/Gj�@���&j�I�g*@UX��������D��c��Z���Đ)ʕ��ib���<*(-�~|{��G���{%��y�ۗ�"�F��H�k���.�|-��C�1 �;u��/� La��+ ԗ�=���4�u��J�vZD�դu12/M}J&����]�
W���ekVcיl6O���^zF�*��2U_8r�d&��O�C���,Uj��@���fp�b(!�T���K+�v�͋�\K8��b��C���R��TT�+c81�EeE֘ l(њ7�������FS�����T��Ni�h�}N�	���.�i�ַ�W�!jX�@����6d��5�JXU�>p�r,�/	�G#}i��%'_|в9X�='�x�2���"�y2���T�d(~��?�MLq��ip)��#:̡Ej�9���|sB��D�A��γ`X�q	'�l���I�7`�})�>�b�t�|�qڸ��#�Ϯ�s�1��aƻ^��7"�$lW�ˡ<��7H����#� ��w�9��|�?�^s����D���?a=)�$}17�Z����o�-'��רL.G��2�ј�0���;F3y�MQ#~Yɯx櫜gmC��_6�c�g��Mrŷ�j �sVV������f8b�b�
�-�I@f#�;�o�Z��I�᎜r�vI�a}�©(�|��r�� ���h�Z��?MV�H�o4�wɍ�u�TQ_���
�2�5=���O��x]OqzV�l���V���(�`�d��*[�7e@>��&Am�������s�G�h8��/���V��.O�8�������:Y��,BI2K�%e���_�����W�c�����hdw�6�Rw��I�Dl�vΫ,���� C��������灋jt<�|*
��S���Ҥq�e*�+IA�&�HR��	w_pρ���(KgGN��,�V�s:���9�p+i#�gO�����	��9N���SbkC�`�[��Z��e�I�a��w���K�7�vN���"m�����	?J������p��x\�$�2�-8	:��*:D�cF2
�"�]evugdGF�YbN���]v��HI�A̲x����f���+�7��@$⡆٭�|�\�;��T�؄��ʚ�E��iee"|,�Qk���T�E��Y1����˴&�9����ꮸ`�2�M�o`G��ZU�
��I ����]��r�)�<�rj�/xȨX��dp�=5��w�<�	�;Խ��].�r]}h�(���N8L���F%q��2���g��9�%��<hPK�j��,C�j��K	�� ��m��:�֒�>g��!M����dm�ʼ���vT��$VZ�.�j���2w�;M ���H�V1�p�A{K���`���
|$��� �����d��<���u�5���E$�S�Z��ضm��D0]��?]�]oUh!ZۑӹC P�H/����I�6�g��K��鰖�3��ޒ��"�g��6i�i�Q�4MRC*�-��rBΞ�H�A�J��S>z� ���Lʠ����|=l�q}�.�'1�C�ɦ�t8i�&Cɵ��E;y@�����{at5����C�r3�n!7��nQ����ˬ6�֛;�y�m�Pn�X��B:�ޥ�<"9VV�I��S;d�GXzo�����BW��<��d�m~�9V���Bvo��ϖ(+l�@O9T��*g�i.>c[=�b�2N�5�S��3��ل��G�dX�á����_�/�k�^n� ���n���Q=L���Ƹˑ��r�<�������b���*���9�l]�
�Uj�XQ���s�jxQ�ކ����[6���-��� �߻ ���OC�lV+��ɷk�lE�~ˎ/k	����UIPR02q����
�k��ph� «�BS_u�^gh��Ę�4W��3^�p��/�K
�lk�<�CVc�}��Xx��۫1uA�"��7����׌s7����la������)S�oШ�bwvo�3�T�Lj��Y���Iu��9����1��J�p�0Y���0�?H����O�<7e��%M��=�x���`Ӈ���q�Z�P�!A-1�����u*ӊ�c����[��>/Q,h((�a�k\ngu��!_�<��j"���:��.���OVg��P�Fa=cu$�R�j�ܼ� ��L����0��@߹�hx�e'=�	�,F��J�TsVv��h.��E�1���lU�؉nE�>���gf����Ͱ���9�^����K"�H�uU�����@X�n� �\����/l�8SB�`2!�MF����^%�����cq'M<"�-M9P� Դ�rR�S'9B�觞q?mq����q��̣W��D���gck����i&D\���O���W�4�k��H��jO�/P9�C\?HO�b^����k&'�ì+ϧ�̮i����'`�#7wX�����"�Tv�Q�Udu��g$�+�i�BA�7�,Ȑ�r�;���r)�Z�U��JOl�qFu$��n�1{8-�E�e������Mp�6h��T�{�gv��'\�]kI}�:�r;����C���M��N�R�i>)�
����Y�n��g�=�u��F������xW=G)����!�m;yY���D�G
2L�9���S��\)B�{��Q ��ޒտ�}��89[�x�n�M<pگ��;b�L�������\����ȇW:�h��wPY��\v\!�zR�+j*l��c�(��5�qF�;<�3e@w�g}r�a�?��p<�p2��@wF�u��\��azh'��K��X f�K9��^��V-��1���S��e���?���(��#D��u��`r�qS$&���)��УT��f����WN��U��^�
@�+��r�����|e6^�<MV4t�6z�c���ә�lJ1���WB5N@�� �V�z�3����������QNˇ�{��4f��λ�?�t�!���^Nú�*0�~�^Z�1R[*;c5���*�u:'� Ɲ��8��.�}F��yY�U(�������%E��&�<�=�~�Gn���- +23�?�R��
>���Q����(ݓ9*i�4P)b��מ����<S��	�l'4rOqg�]X��^�b/Qg�|[��-ݵ֨��H�W���-D)���}�$�����mbi���&?>U�Ki0�D�q�ׯ{���s�J�ē����3������,���X��� ��k�ml :�>@��s�L�)��0H���",!�`�;���4�8Ê�?G8���Z����s�G�M��Բ�pFw��ڲy����-L�a���]JR�[гc_v��7(����R�׆,���9[r��vƉ���Y�T
GߗH�(��q&R �:��{}���zfb��A!���C�L6Q�#ey�zPn+��=y�.�f��b�AE�2A�mZ8\��i�j= d��'��ä��ji���LK� �w����a�N�~���� �~�nZ��µUu�l�Ɲ}q��Q�F)� ��u?�j�/��O�:�4ވr�z�dyi@K�0���W҂Q��3\��m2�jg��xU�zi����h�]�LW
O�&RH!.�U`��Q4�ȷ����l��].��?]��up�i-�U6=����6��$V�w6!��r#M@C��b�d��V�����T	���eN�i3׈*;�d��w�﫝x<��d���t�Lu�ƹ����d�A�4-H��83�iS����j��?}] G��9x�1y���Q��a^F �ȨM�a/Z�Z�ݥ4~,�P�;�T���p����	�Icg:���+[��~a��t�"�T�f;�ga�z�냄j ����'�Q@n{�7��=8F��|����A_!G'}�R RE%�Ɯ�M"�ٹ��h�a=���C]h�t�"8H�ΑA�&�mj%�}�k�L�ݭMq�~�keA��ǃy��!8Y�&8�
����]ZY�.kd��Z8��F�?T[�-�7�V%���Y���P��hTX`0O:N[�'�L�:��"aKl$vi��'��,b;�IH���ѳx���Y����8}�S��b��	g��܅P/�����7Zp�>���+�7&��T������;�H
+fo�܎%��p�Ec��X��C�6�1����#@�ǭ��[nW��w{n��	�m�*��&GY����[%Bo�.O�>��1�N>��G��9����v�"�LAR���a�q8�0b�TI�5ԷMT��]Sl|�Zޤ��|��\�gf�v�&ӟ��t;ߓ.p)�]�>�&�=�,�
����]���p�����뛃�Y*�6�)����)�7�����Z3��k����%��N�Pb�xn�Vc%�'cq�v�"�~<�$>�ϭ�MR2�"(i'u)j��Y��'QR}��y�*����&J���q,Vۋ|��˵�p����>T��52�z]�!7�(^#)�Uj��j�p�T!c<��d��>*A�%7+�@j��'��[�7��:�~4Sp��oO�E�j�&�c�D� O(G%�$�vc^��K7л'ͯ2ƈ֫'����՗���ْq����Y�u�ي�Ի�k�a��9ϵ.Ƌ:���Ⲑ���G�:��	�ӎQ>0�p\l����͎�2���rjBvD�̌e��L2�.y��3Q%Q~r�2.s,���CN�����f��E8�{� ��:o�6�ǡP��3�bR��y��Rz�(}A����aN���唩��0���K���[~+?��$ K�cL��vH�q�o�pf'u�{�{7�	?IBE���
��wQ����.�#1��Q���y�La��xF<0:�}����0�b��Z|���Z�v����U��N�4B��Xu&` $1��;�mֶ�J����ƛ��V�n����9U�	�j7k��X��vÎ���7]�������#�xW��qF������7=)]�ҚP��%��|pکIg����z:�0��G��4:�2@o�π��i`�|���̠�l��EC�r���.�ME��}�i\�O�:Y�������s���P�[�:	 �_��.Hz�Q�@O�;��x��PˈR)���k���<�r����s����
K��D� ��	)ndQ�E�Y�̞�s.V얦|�E��8��֛�Ԏ�<-���v*tCE�㾒n{����QY���9"r���k�S����k~���1w��$-9�)��d�`�^qҡ-��3�m�s���9��eP�� ����wț��y~��A���O�	� ����mƸ݁�o|�O��FΪ�<9��*��%���ۊ$��$�j�@w'A��f.9H�,�y/GS�3�6��=v8��ހ���Ŝ�N��$�Lu�=��,p���b��(~�:��4�E�`e�B5*lx�6����ޡ41�jF쥴�xh��y��N=�� ����:|Q�JNK�4�(�b}4��;6�rB
����P9�:j[�<n��c�7��7#~9k��x/��Ez����8�u7���b#�g�P��2�28�Ղ:�qQ����U^H��Zs�4�k��E�l��">�W��
&�D�t �{rWrC�o&z<�gE* �a���WF�2E��1�6��j/`� <��ɽ`���)�߉[��n��?fcԂ��}��z��a��](��� ̂��ɺ��3<dH�� �ðS4���}�"z��7����$[i���3DY��uL>�	�����w��,O�U%�D z�h�f���<e'9�����1���Ȏ>�/��� F��Cˉi�ˁ�F7����T޴ҹ_���W�9�����&���Cp&`��}y�P��Z�(~���CYg�˄���|�Lͦ�(Sa�i�x1:��eu尅�)��F�Pñ`��
K�rU\�YB[N/ �C�%Ѷ�E]�c�J��O��ɱ�4�6���1�z��hnM4ތS\҇	��ü�!d�uov��8��9�L�?8d)8m� ��� �����ꑈ�
E"�{�g�7�q&7�aQ~��ȧ��z�h�ªd��禑6��FfW�<�pR��,��mP@���*�r\�%	��T��tj}zi�R	�� (��ڏ�i�K��`ލk�h0�?���*�N��枃&o򻖁�z�<3qҪ�����m}�������3K���09Ћg�w�teL'��"F�@���]��F	��ky�JB=�`�!^rB�j�(F�gk��ƌqR�%,���S��#��H$*��~}n�Q�;b�V|�K�s��_�)`�u��#�0"#��ۈ#��X�r��s��/�����:�'���D�ަc<��؋��o�C�q�x+����g��%l���
[�:]�8O�
�ROAT�.�<*U@Pi�ZI[��r�2 ��Q1�j7���F&��S�8),8� ��GLL<��,.��̆�:&��T�2(Qŝ'GK)����X ٣��K�pQr?t!m�*#�1�-����%��;��^��ƞ�x89,0�v�4J��W�+'ʧ����,*�Q�&�S=`���b��F��� Gr1x�c	&!��� ����Ӛ@�A���:�M��bK�-�b�e�6���W��|�O%��{�q�����ʠ��zY�`� ���dU�F�z�ŋV�0ǡS�ָ���|���c�s�|�=��:2/������bbt�m���3��
�[K�*9�BS���@��G�±��i�R`�I�-C�>�U��R����]Jö����Azf i�0@KE��[��A[���ը~�����r�n@��S�5�"״!��k ^���=J�Z��<�=ggPJ��dl�5{p(�q�Z�5��_d��!��fC��W׽]�U��>@��'GR�w�&�V/Y��U�N$�C��c�#t�}»l@x�-��6���e��H]/$aF�O�`��lv�=�HV+ʲ�xk�N�@���:qk��*u"����Ƿ�:.m�T

0���B�8���vj,�v`[��'���H냸��~���[NE�R�`PS�>p͆']���<���Z@�����^şC}�C�����%��ϙ1����df8�sIG��½�����Һ���;��ګ�����ϔ��b��Ei��Ώu�K�)�\�>W���N��B��0"��Ư���>�l^gT\z���9��Xw�*��>$0 ���q܂�8�o����J�Յ��bD��YK`V�u���k�V9GJ��6�Mn�4C8��0t�������]D���Խd5���<[�����9�j����L��k���i9&�H@��O�<�M�q_zm�tR��u0��3�kB����lE�49-g�x��{�k�7Y�+�!�q��y6d����,߿g��#tp偒rs�S�Ӭ�j�n���E���
-۳`�'�|`}9I�FP���d�L6�̾2p�J�$���y��$6��W��rV!nSwzY����A�7��Ԇ|[��QH�?�M<�J�xފ��i͔ta�.!\���@S~�e �	��Um�m��q��B���I��)V=.Kg��X>_��s�h�/,�.�bC)z�
=۵[��,PP��:�A��N��X��8�ZfI��It�7ы���ǾT��B53�%�ʨ� ����Pjy�㢩��v�D�*�դ�4�{���ht�.y�_$�����4�
��3��#�Y�����Q9=�S)�MpZGQ^Wl�h$
b.��
�3�]�{�v��w{ZWWT�i����_kؤ�6؈1��Bp�2gT���7e�a"[if��LGQ9Q�:�O��䇚�܃f�<�jEYa}JD�d&�9���Y����3́�����m�tr#��-�
!��0h�6��"��q����l�Z���ڹ8���HS�" BI�G�WY���K��C��,ªVa���Q��e��_\�n�-4��RY�n�z�"͠b�H�M��)�:�S���	ׁ��A�^v��H-$\!}���ih�������-�͇2��k�5ĳ��Z�+e�9�(rA�
;��_El$-y��s%�#J�ۿ��F�dg2DO��0���/sE:ϗQ6a��*�kh�6����D�C٣�}�Zv "g[��?���>�D _ۺL��5e8ݞS�B��#�B��F���N�uJ�-/�* ~D��Z>u�g�e �ۻӑ)9�`'�����3�)�P6���i4h�@sܚ��h�V�@Hye"pE�h9<��SK$P�*6�會6ãbQ/}3�QD��9[��2٠�d�b���e!u�����O���$x�#�z��X��&��A5|�;�qV�� mx� ��c;VT��a�j�㮝�J�P흚�U���;vc7�Q��1�<�T�ذ�x��WyQ��?�29I�� �aw��R��V^�ێ�?}X�Ο�Р@�:U�j�{�զ1�&��!��3�m^��:l�����D�k��V�d��z��k�roED�H'�����9��W,�X?�R!n����0�oC:Dٌ���ݢ�ܢ�Uˇ�oY��d�]v0����1Q�A4�h!Bc z("aD��m�St.Z��Zd)/ED0��F���~A�eʀB�Eʇ��* �ܕ��h�p��U��x�۵��LA i�
D`�����$L �'��Y��N���2�x��8k��!���/ 3��V���ǀ T�m2�;p��Z�O�~'k�6Lh�'f���1�ı8�'l�6�P��S���A��RɌ���(�Uu{��'߶T�{ �#�6� ��# ��x�̿,��3_�6%�Zj��%�.��M��`!#��о��E�h�J	�����]�Xp-nA��fPԓ��/@��k}0�؊��������9V"~��)���b�^<BD�����Pǎ%�Zn1�a� =�Osar��so�yC#Ҽ)��\�������iʥ��l�e�Í��Dޱ����+�Ժ��e^���pQ�n4��O�
>�bѼ��	.?��pQ�;s;������i5s����H+�#�5|���j�-��+�`��w]�p/�� .s�=G}ɭ��mH�#4�w�!�����ƴ<o�*���}l1�AR��e�����%bEqF�`J
�����,"7UE�yw[�/Am��	��9���_
��n�d'?���J�>��E��5�|����(8[#���"U�u���!�i4�Җ3U��Z$&�.��3��U+��5�)��r��p�#)9�5���0��e�M�ARo���GXẃptYCigM����m8�) \`7�4�^C��_�R��a��r�3�X&� �H��m9���<n��)䟶64�ڱ�8,� lLms3i;�� ����QՋ���v����Z!���ht7�T������#EvL�ܬ*����}�)!���4<S%�� *�v.����"�-��a���M�Di(��LF�URh��r��Y�j��H� 5o��b���|��֞�t^ؤ�碕�yU~��egQ���_r�ڜl�|p�O�{0u`��B@�M��^�bS�6�	��3����@D�p�";��=���8x&��� ��;���~��g� z��؛���A�H��Y�+��|ž����.P�0� �踡�,L�c�9��ejN?�JD����^�,3!��%�ܨ7�*vT�W}LI��~pg�w��րt wԠ��֦ԁ��D<��$N�<��|��ض��JDJM�+��n>�~
��%1N�K=�����_и�U�KP��E7og���|D���u@��c�b\�$Ix��y����� ]�*���/����c��<$U�<T�e���q�����5H�R�@�!�����v��pH��o"��/���