��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?F���P�T폖�f�[
�F�/f:�\�C4��r��7h�S����B��y��R[R"ox�o��	���3�3��
|��`�gWU�d�_�гU�,�����D��(ۅ�gd&w�,��~�W~ߟ��oQ�?�&X?��]\�G�����j��-�m��R2���}��������Z��E���u��7+��W!����
��!�59��Li�' �Ù7і�w���P�DL�^t�;�A�d�FU��lN�K���gY����%X�e]8�����4z����� �6���m�z#Hx-���b_�5xMô�b?ώD�#�Jc�l��ȕ$(��
4�]���^���K�+�#��n�W���d���F;�!i.�W|@I<,0 ��L��9dҫ):���eFi�
#UmyFh/8Z����89<m��nZ��*U+*�<�G�kwN!�+0�����8L
�����Q�]d�0E+�55�GUgby>��K���u�Uk~�����bSV8	h��r�.r2������	�J�~�M��U)��́䵨��1y�XW8�;,f��%|Q�Y���F��c.�46t�<��'yn��sn(�z��X�ccʐ���bb�(v��*fr����B�wV,E��
�bR�HO�R�vd�?�h{�ڎ�xm`g�Ǎ���4Ц��?ӢqX�EB3gI:(>�4^�3���8�ccac�������Ma6����٣�Ye�WJiN�s����)�Yg�ב����s.ӊy�eȸ�wS	̽ԁ:Oz��9��f��i�q�����
�P2;�U�z�϶[2X�I*u�n�������%q7�^�:��������i�Cre�Y�&��n�W^�ܶ3'b1����h���'k�l��;���]���=p��;xZY+薠!�s�˸}28:�1�x+�5wRnlip��wY�S���ѡ/����4s��$�`|�-.������g��3���>�GF��� ��@�X�N�gP`:�G1��.�{}��(?rZ��u�/.d�"=�{���Q���}�
���*Г��0����?фa���ܰﳪ��oۊ5&s�Z[k��l�W��C�����-��|���	�V	�t�t��pa�$���Tg}-P���ֵ��?6}�gu�3&�u�< |�-�B;����[O�n��p4\�$��*m����W��5Cq�����i��'�S���(a����O�|}t�t\Ž��{�`�Vf��D����#�+$�����5�����AA��J��K�7�:�(�����>�Ds�Aɸ�\�!糨��vXw���b�AP{����W�����N	٫H�ݗG��MP+�����s�p6�v�9�p���E���f{�H&RƳk�$�2�t�L5�E?)�|l����Die|E1���B6F����B;��ɵ�'��z3��m���3�$t�J��s���>�e����G@/g^%�Q�#֚��f���`�r�"5��feb��:�������ܭ7��pL�Z�1�^�g�Vc����plΓ�uQg@o�2D��IW^
�ćJ��9�
�T;�Ӥ�P�g�1v
�#���K��j�"��C�`�	d�E9�2�;��gX�~��{�K��:D�s��b�GiĀsu��T���O횦���"�}f`VѪR��,���D�N�B��f��%h�J��͍IkK*�	&�W��*� RSI/F�9�A�ڢ��
k��#W��G"�0`��_�7��D����;�O-a稬��/CVB��'�J��V��u{ o ����g��uiV'���i5t������f6��A:Z�b��Z�3o�B!��wB�3�����	h��n�+�,g����J2�Ln��D��:��s�`�|�4�4Q��䶤�$�M�~#T��m�#���!��'��($�<!s@g����J��0X��J�!Dn���i�M��.��u�v��j C�D�"K<�u�4�/�(و/O���:�,����Y}��W���$N�a�qqu�h�nV����65�8��ا[���"�����v�53����JTT�DZYU@I�t������?���!�_żwe���V$,�@�/��Rk0��[�a[�(/�M�WO�	�_���ք��g~=E���Eۄ�e&�=��|�Ӫ'n��+��vC�w7L�����7%��=��Kq�YW`[z�<�ShF���M�g��ՑRPY���2r�|���Cy���P�sjp�6TւK�Vײ=BN�Y���<�#��,�l��	����?O����f���O-�>�#��ue���,2���&�}���,m�bH���c����`-��[�_�S7	�c�����h�j�G�?d؝VR�0j�O�'���Y��1���33
��+t�@��C5;#��ڒ�Q9x��'v�w��F��6��]"�d�G�?�	�U M&\�*�Z��4�4r9���g������j�PB��nt���|~ֶ7@7{�@��(EazJ}�t�}�a�@D_�����پp�lY�+�$m݊�ٽ�g����9q?(�i�Բu�kJ�^s0��d���*]��Ff���X�>��	3a�Zc�A��	a��F�����}=� i6�} B&��A���*�a��E�-���£P�ԁ.���@>GVw_⠭�6F˰��9��o�9]�+K\n�jM��LS@��u9���Cj>���&j���4=�[��.�������q\��Jv��؞����������S	���2c��HG�y�/��ie�$�>��։y�zJ���gv�W��շ�p���/͟��Mj�W?�B�D�(��V�@�V���g�R�ˊ������ܫi�6\-:t�{<N�Z,�;����s�s�[���2����9g�>&�y�G�+��^�@�K�Kr`4���c����������7����=e ���$ҝ�I����tu+�];�ܜ���SH��h�N��7��R�-:H_{Չ<�_� �|g;I���ڎX�9%n�Bi�s�G�5/]�[�X;k�̯b!2�����>�m�m酽^�kqu��ڔf	(�� �dO��ً��/1(w��'#<`ټ-�>Ӗ�|0$>◂��:h��ԭ�g} MW����J@����x�{�dd��
�{�1N^H�Qi�P\R�.�I�~�{��j��Ww�X�jR�4c׍f�te]}������L?\����<�;�O`Y+�%E 2��T�),gx$!�M�	g�r�[�!�����V����[�W;�i�s�ba�������K�q�mA���]�M�n�rX��;���h ��rk�q[�Q��8�g�,��
���l-���p%�:v`�n��b���I���B�E\DA������f9� �F:  ��a�~4EE��ѓ�4�������O]0Ⱦ�])��O*���A̻���-C�L��u���.�a��(��^ �	*�'�������SG8���S4^���n����ؿ��*�hi4�J�?u�v`��+�q�	��&�NZ��e	x/#y8�$a��4/�Ԃfm��ȰۼHr�9����^}�:yKx��Y�	�:��0���� ���r���
���+��U)��h�gq�Cs�d����Ĥ��?��S���Eߨ�l�-\�V�?5�:��K�<+0kCa�Έ�{Fa���vP#���RO=��Z3
�րM��b'�FS��=�C]������p�+�(֏k6R��,ͶU��j���Պ4���Q�{����P���I���Ș�T�]}�%\y}:�7���hVw�z��tb�%��qXq���5�EE��Y�!���-J|�V���C�����ߛj��?�.Rz]q�%��E忊�գ�v�P_�2���	��T�Y�.���x<_I_�]�	9'Du˟�+k��#'Z`�ԏNb9��!|�>.F��L��{�(ˌ��4t���D	e"kN������sT�b��weY@B�,W�tt#��a.䙊i�0��Y�������yWh~��{9�7��˩�	��JUw��������K���ɹ}>(r�s���[X���i����eM�n��� ��L�Fc�IN����.h+��l�1�F�:��)�-��j6�^bo�"8����X$�8���0� �� 6�WB��.0���.�'�H�k(�e �7HYc﷣J�_�{]�����ըT��q�o�yn\��e�c)����z��Y�lN��%_Κ#��9'�K��h,�"]��춿� t%M+�%^�!*��1��,�3h�nd��^&�
�� 8k�yY��.��=*%{�v�!�t�P:�Uj�����:����P�f����Rb�UI��e�O GwY"�D���1	�"�]0jդ�"Jl,WY;�C��f����h .ȻDK��KS�簇`��
�#����W[U�k!�k×/6za���r����ӵK�T}!��W���ߙ5���I���Z*�������T�ݿP�'nP�aS2H��c�9�R0�R��NL7�e�.��^������4�Y�X��iu��fy[� ��/��W��Y!Z07��j�N/����I4=ҭ��nf3�~��A�䭪�Q�:���������>%�������b�0�'{ �<K��^���ld�lEVu=�!8ao���GM,�Km&��.���7�1Rv���@��+ϲm�<T617�r)�6��/wd���Z=��@�����}��f�.3��Ύ�-�|�)�l�ÌЁ���b�<����'&)cC)����*{/[�'Ԧ/3_^�s��!f���4��F�{��8�z�!Wv��.����:	���1�s����lK��cT׾#OC(i�S�T�S�aw:HW��X����؈�j���[p^&���B��o�X�|����S[d���)��"�q~���ӠF̀�|����e��C\A�h[wdH�7�ǁ�R���9������F`l���\�$D��~�vWk5e��.�\4�!*C���I��t �_7^7m�
�H.h�,�_P_��/�]���,�}�w�k����|5@ll��w�(�&Dk���Ǳ���.�"下ᅺ�l=�{(�DK�X=�Ώ�p'.Z���# �$Q݂��14�b^����B�{ХӧJ��H'�57B���B;�$k�Z��Ø��3�쀠Q{�� ��0�nv�ɸz����w�:z�H�$��}E�.EI�����x�8w�pw͛�r��Bn�ˤ��&��l���}A�Z)j��؟2�mڡ������&J�mO��)����R���.>*	Ɣ��c�M�9{��(g�-�}�p*���q����x��I��X�b��K}��E33Z�1'�����$��5�^ @�6>M�a��,�ħ>��� ����|����ik�Z����D�|v!(�ś�`���<kel%Z��To@h�t�w����Pm�Q�3xA���������G�)KЖ���_�y�+�H���Vp\�	�SB^6��3Q���}���&�:��Ǩ�3L��������>sJh�T����GM��@�K�4]w>ؖ���SF�U���U�����qPp
C��}��(�T�l�WV_g�[�s٠�7}��3L����"/�hp�ܴ�R�ޟ�w�M��ܮ˅{B5<8ԡ7�j����⼄��po��������ch�	� ��g��Y���B��xj�}�R����d�OƩ���,'D���/��Z'�Yd�3�٘8Τ�J"d����X��1��s�G&�(���ʷ��D��T���}�>����&C&�_�5C�^�QM��)"F	��B<+��|l缇��;�E�W%S��� N��X�
�\�W�W�VI�+���u�Td)�?	[�&E�,�!oM�.�MƳ���H¡�\�#C"]�K�A@cj��rʻY�b�v��CF���װ�l�6�y��Q�C��%e����P�EXp4&��v���`��-�`�����r_w��6ï画˴'�Z�ۏ��֪-O�㾄]�n��\�ň|'�l�Y-��H�|����0�&���ƴ.Ʀd������@L�,WBT,���u�?s�WL����PY&B?����1�λd ���la���_�sp�-��/p��Ɛ7���F~y�Y��j���jo�v�d,P�x���5�Ɏ�f1ٍ"��B�������S��H��Vk���m��K�@O�g$"t�R�9W���K�N�d�q��*	"��)�ÁG�H�&*���Kv*^���[�DJd�r�*Q�:�j*5-��6D�p)�Y*R\V��.$q���
b�VFƂ����_�ɠ��p6;�x�4Y�-���Z�z7��6�i�(
�kJ&~�.أŚ�B
OR?2���g�7A���{���o\x _͢U'anK��!-Vӕc���OD07a�����%�Z93�w��fq#q ܎7��7Q�����3���B"�?�@�5k���v����e���9�Ƴ��1y���m?^bi��U]W�_SѼfg+oĨ���P�B�%��I�N��%
�1�w�ϋ��؁��JD��}1~ʇI�g�\<�1TJxl��ݜ߳��X/�e�������*7s�nb�1q�!���/����2q� �۴P�y�&wP��չ�-�L��D:U�]zN&c�
�dܲf?��`T��H���D�TK�J�NV�o�N9ܪw��z��4_����?hj�'�&jp��NMF�ƣ^��	�\	YQs���^aJW-��g Ckkv�9�"��40�En�$-���?;w�����������F=�Uq�+T��*�b�ά�J,ي	��ᖔ�6�8��5&Mq�"lLiCI��GF��A}%$��z
��qɔ�	�y%藎U}��8d�*��M�D�Y�J�󙦇�k���ê	uή��T�W��R� ˴ W0�g ����+KS8����ϑD��;�㚥�3zw|yH�<n�i��sz�� ��N�M!~�����M�$���į�%�dӛI��������uO{��S�H��R���Ԃ�8�b�i�'��/�OP#��?�3]��v���񩽅��{@����݊�Btj)���5 �j����I��>�:��i�v��wE/�Vw��Z��y�k����va8�4�3&S��K|�ќ�Υ��Ҋ�w!�� ː�iB���~a��L�>N��(�N (�{QS97)����%yß�ÊٴP�A����Q�t�p�r���Z�K��!�|׏����|%]�=nj5��-��" oຌT�FƉֵ����	������RV��[C���>�T,�H�Տo`��Bs=Lj�a��X ���(���(��!H�i[�H[�c:߆;&1����VN
72�Vm t�WJ�{զh[�)Q�/+��I��ﷆ���xr�o������d�P�,k��u��^'��H�&K��_C�s �[�{`W+��U��?b6G4v��i� �x@�z�|�,[���f(�����V�gs\�PZ0�̉"�oH�Y�@�%q �2��b%�(�_�7������i�(Z�k\�zpL�m^.<B���YGқ�\Vr[�u��|,q�l��gЕ��|�{�B��Jz�;p,�Xp/#[}��
���S���5��b:n�]�ެ�e�.�H�����+ډ�\"c��
��b����4�Ў�H���9: ��:�k��e���8�Y;4��������G�b�f�b��f�1�����.�Ft�U�!쟅�4!�4�0��tI�g���ºڻF�.I�*�H����=�눟���%��J�q6�;5Y��֜JQ�Kf��\0��pؙl�;�����(���N�����mw�P�V�B���ʜ�{�@<�O�_�(�;�Es���|?���H��x܉s1�ޝ�����ĩԉ��9ˉ
��O������|H��ZF�XX4m�@<�S<�}�ka���m4�Sp軺���x�Q���@�&�2bGA�����k�\7����H�KB3�~�>w5����Ex�Ñݨ=#��X���'|-./q��puf���o6[Wz�vASsF3Ԇ[���0�n�Э%�#/ \6�P9	r���G� CxНux���ެ����/�JJ)ĵڻ����� F�{+�B�vv؁6*5����Jb@��x��C|��;�����B<�d�[�?�����i��L�v��'�,��^hF��8ٱ"��1��r�:�<�-��HEg�V�l\J��� ��Νܖ�Ӗ�<h[#�e���qM�r�
�AD���I��%�R���^��H:߭�����<4*Tt~��"�uՅ�*��Gg�a�-�H�E�^��k6�歬%�&�F+��`��TI��0܍Xj��(����Q̖G�w��>���I�M�uYh��B�*8t��U:FT*d�]�s1�H`�jE���4�����l�u�4g���1�oe0ՁL���W���oe�D� W��`�G��i1 �pRo����ܹc��L�͖~o� ~?�z��'�e�=�\�S*�ߋD���z��16Zp�'��k��!�8uBi N��cff�^\���&_O�e�c��I7��0�|/�c+��X��؟ږ�=�b#�"���4O�S���%�?�NK�.��~�QX��|��6��o\NyF�~>F��;(D5Z�J*ϻCte����L .Vj�����g^�"�,竈�U���"��J�~�	����IK��ңbY�bO~�34���Z�F�"���o��m����"3���v��Pg3���^,��}�Xڂ����i���+5Qi�؉r�خ�-�9�e�Di~��²�ـ��ŗD���+o�;��J�6�x&�,�A.x���euh��R%a
ۛ#�,y wA���C�jx?k��#�1":�D.߷D��3���=F���+f��@�'*zv_�DH (aМύ��	�;LHNb�	�����t�!�rCIn['�Y��ef RW̴}{+�AQ�u�)w�J��?3��`gQU��g%f-cލ��v�+X4���l��b5ň)]�FM]�y��G�#q��AF5�J÷��3~8;T����?�G�3���'�"T�v:@�d�2��y�����߸�T{������-���G
S��v� ��&	�8�p���	5A܀}��6�#y����7p��C���C3+V���|i��N�V�Rl���}n�(A��!����*�sȓ .Q$�&�ru{K�.|����c��{J�[d8&P��muɯ3�w���3�m��*��\��5��&�r�A'#z˽+���`%�x��q־�k�1\Nj�k}뜻��e�0�G�:�"��w���g.6��̑Xm���F��EU�+�'�|~���x���鯿��7\.�2����Hx�U�q�u=LT�e�\�tb�摁t�w���IM�5#���rNw]��K����Ţ�)3�)Ra��&�4���o[�p��>� �P�9��{*M~�XE*n2u�.['T�`��H&���3�J�>�e��E��{�:`���t�ݔҡ7+���ܗBZ��/p�O���H�\]��Z��@�8l93�5sJeup�2������9Y���E��(<�s��M舯<xF�N�x��'iH�>�dJ�|�}p"��q�@ߔ7��S�����'ƣ���1�¶֕z�"�qO�
��ReHV���o	�s#S�0V���+B4n��0��5w�]V���TZ�w]��#F��(�#�h]bQ�SS���<��-s��ኙ��`м��0�	���`S��I�H�a�,c���P���bHч�	��g$�� wd��;II7�7�NE�m/�%���o��߯+M-#x���t�~[��S�-�j��}t��a
,�(�!�3����i�
d�t��T{�~zJ@.p����u�*BOǖ����C�^�C�Y���y陮T�����CI����>Nh�����������M���i+46�(���
���G�M_g �%��M
�b����Κ���9+&ݱ~QJJ�c�,���S-����^l�Jel�}��jP���w&�W��:	�_�½�[��lK'�n�T�i<�#!���MV�"�31{�~
g=sSL�����)qڌ��(��vz����.H�V�n{/yei��>sQ:�?h�-��*|{4��!R���w�3��N�⎂?��#���^�:�����^��*MUg�9�CY�(�
��3�(��0��8�b܀�!j�-�Q"J��%Z�D�V_qn�J�����R՛�K����;(!W3Y͗w6�_�&�hn9:�X~\�\hld���ߕ���yl�
��擺2˚�q�n��h�)�Ģ*��KV@H��$�F��&*��;����)Oǁ����j����S_�PM�5����V�wg/��9��vs�|
�N鐤�y���X�G�+O����WY���|��D�ڶs�U�5P��25w�s)"ҁ���ǲ����Hw@�65M��?�g�w/� �_�Ć���v�|��tI!H�	�y�u���q �vpqT��Q��|������E%@FY�5F?�6������Bn�3�A�԰ex s�C�i���$��aO�`&|;��K�8*�l��o�F���|X�)���M{ 
��*=����q����9n}U�?���@��ș��<���p��E�F��(�)�.��o�V�R�[DIZ�F�=�J�R(�p�� w����3h\��:�����L�;�L�^O���A�K���b.Ĳp:�Kc.��_���fp�D}�ƙ��BNsZ$l}DH�b����>Kb�}YG�C7��J��b�I�o�?�y���U���mae�6�xI��s�b�+�=ޢ}���6M{�j�^r��q=B��=�US�jm��LY��6����ĈI�F��}JՁbT����&&����G$��E�+S�����fן���Mz�B�40�/_����I^���������.����)p��PG�2f�QFP1�(!���������=ȻnJ@���~��*�59�x	�Vc������9SuV�hT'rL�ƊM_n]`��u������}D4�}B���|�'Dv����������ě���O�
�X ��$+q��:�Z(�qM�Y�Z�/�;��g�L+�e�z�*����7�<6���
3���.^st�C�.e�w)�i�ki�X�]w�9�:������sANe�,W�o�������ړj3�����Is�9?:4h]�����2$X]��Ie~*7����_q'�'��TF^t��.B���M��Mt�{n��)��̕Y�����8X��Ae��а?���&��?���l�� 2,4��r ��l�ίƐ5��ِ���?�רg"hL�WmV\L�~k}�@���~�i��F�:��	�J7d�%�`����g�dR)E�_��S�gZ��i�V��c�.��=�4����:�ut��s!v�4��:bm�W�o����j�IE}��s]�f���(.m���[Vɸ���"�8��&����i���(���H��f5��b�~���z!`�ul0�^��5�Yh�z�h�;��YU��!�I����~w���Z�,F�g2�ux�W�)H���3���q��?�� �[�2���������>*o�w{��_������QC��J��q�~����<�a��G�za��qz"Ozy)���x������𥉉B;[uHG��;+� aС�$�*r�r��+;�"�24n�������i6�yj�����yA�(��3/�m�~V�������?~��о+��Q��7�z"�̰jlA��yo;5?�x��`↸Fr���_��`����REn{�V��F�U(Ey;Idjh]���֋(x#|��x���_��~Mnʹ��u�)/q��_�K�������I�����WvD5�J���8[م��Te�S�w�NQ�H���xVW�JG��(C�ۼ���tUO9�g�-����vU��q�����k��a��e}���6���Ӥt1R@�ѿ7�/�Y.)/��_+��6�e�����k柤��J�.?3��y���?7��)u��� $����Lf�٬ﭻ�DF��������]��Kd����鳮uA/��[����~"���|QE�V�܏��4�㷓���ދ�A�6�)�}��V��־�<��V�G��nT"ql�,ͧe9�.�N�	cD��@��
T$fv��u����hs�16`�p:��!�/�P�9H :���X$t���V�q]�3L\��W���MU�2γ@��\�_�T���+�	E ����S4񎞵06M�|G���y{�'Gs��`�h��E�[���3/Z�;�""��^Ĥ��:�5��ė|ֺ����-PM~��D'x"��t�颳�|`�:-�9vu��k;�)7?ICF�G���'
�#�A��_��@4��	[ ,t�G�٪v.��E�%�mm��c��ڐ�5�kg)r�R31y����i�Y��(�h�ϥ�T�P�i�&�EkŲ�.�/?��%ܪ���̹ǿ�����!�3�ǲ�,�JA��~��ݯ_�ɡ=��~z1�n��-���b˸?t�o��N��N���1Rp���+��_Bۃ���pb��1�����)�u�Pλ�=�F8�ۚ��Ȥz�xms[�0���C���X�d���w)X�%A��#��,���ͫ����*�����,i�f8T��y<��=v��,m�d	߅��(�z>f�#K�o�$��M�H4K6�ذ؆X��p��lF�W������~��x�V�<6A"�����(0⒪�����7��`��|ds_K���6�<���0 �`�>�u��h��y1�ԭľ�e0����Ck����-ң�Bj�۶?�����
���[��y�����B߫H�0,i��a[!z��1~`�Ύ����z0��>�T��t 9�3h�����俠�7�E)H����4�۲���z���5X���I�$Z�b��0g��RMߏ&��_ߔ�"���&J�%���vm�JUO�|XC�L�����.M~2(�V�L
~���T����z��8��ϝ�h�is��[�,���A�)�����&�/#��B�լ�2�V4�흏��!7B�Q�=@iK�
6�>:��x�3���X)�=�U��"q��ј�&!���ʿ`'�'��f�֥�R�c�]3��qvi8�]ָpɁ��V��V�Z��E�Ʊ�iT���?kL8JtPK����lwL�3��LR��lw�nUWqXD��M�,.��B��+w�p���(xp䰋
��Ђ��UYFG���tQ�+���?�̿kp �ԞB�F��a�K�hp�ƃ��	��zh�fI~=}�����B�,��ѯ)|�b�U��T�e_q���~M��:��Zb��Mu8�n�[�*nb�lyc`�FΞ-�q}����H��i��\t�ݱS-k~����Ēn(T�b��?[ՉZ���KN��"����S �;�]�q%m���:|n~H���~�XI��HP�{ԮD��P��nXdܩ��Yi�=8�y6n�+���2	�g)�[уh)~���ۯ��&r���0�(��m5򓬪�$^a�T�:2��&x[��|��(8�j���T�81i1����v�iNBN�Z���?:i��su�y(��\�]M�H'e
WKq�~eI$�u5�y7�� �5�_��n�^Wu?�����+xz�[�E@;Q����y��8��ہBzrR������~	�� �"�`�p60u���w]W��`Ѭ�T��X��X�l���8JP��zv^�!=����@"Y��m���j
��T�H�>�P���H�&��v/��K;!o��pJ��)�t�*8N៌nρX��hK�	��i�_:��
�%v�e�	.��ٟX��)zpj��w��$?�`T�o�.�B�U�p�!�4��`�X�̀֎Q��F�J~1���Z &������nĴ&��t���fEl�%�"ŘT����3!��(���Q�@%܀��̶JRu�~��g���}Gc��"`DF�¤�_�sl��(����>����m�������4v���>��=Qd��B+N�q�-�	=��8�K^�_�C�0��t�V�_��=%E{�02���i����f��d��Q�) �[��0�<��	�ٺ�l-RN�9��(�4���9P�05
��+ԡ��r\��E�<�d�S���CI��#��e>�z�o�N�[aL IG���/4�4|f�� R�*�k� ��u���G�j�˶��Ec��ڟ|	64�����b���k��ת���q����/91 ٝ��F�
�~�)�y�:�]/��W�ŴT׽�������oB��?%ٚ����M��@�@Y�������=�cfOt��3?9��&���NX: ��h+���j�@OؓT���-iM2bTZſ�S��f���r�>�MH)@����&�$�/��S�%@k�J��hZ����k̟�D|��2��`��|È' �-����t3�ʺ��@Kjg�<t&��5��[zK7gs^ː>|tQ�6��E6�Kx������<�3��1�sB�u/���"�XU�O��UDd_l����IC���T�y��Ǌ;>(U�9��H�0�4�˰!��ގ[VCb#����c��ʑf�If(�R�E�Wn0�*��Se�n�������G�x�f~6����@nW�
�$��:����g�G��7k:ե��a�y37���]��]dla��2;W��.9�.J4�ICL]���vd���X�N[U!����yC���yit�|��X�̈�0~���<j�]9��L�W��Hf����	p���%N��G{f�u�p�.�+۔�9̠� /�@��	���䛡��*�GWK�5������^
�W��v�;����o'E��2��z�D}JC�v2w/K�UGGi��e��6���(����-GΨu�hbS8-t+v)���a�,��>b�ך�I���?��g��oN��ck�sj�S�Z���Og�	��j D�^��ikl.����(�	��s;�]��lo9�
��	1���&�S���9+ӭ@+c��N�������n��ҟ،������6͓��|w|xir�OU��)���`G�ܹ�΍>�c�]���B�b;P�$�|Ա@G!�EI��(����#L��`vG�#v���*�j�TX��4�
�)'U^� ��k�\���z\~}`�T�lԃ��g���-z���\��P~��%q/��N�E{~t���ND=L�!��&J�D�ZI��>�[瞆-m�{]2*k��j�.��|�!S=5�O����A��\�48t.�*�UN�7A�R��%qk���(G��1���.KP�-V�1V$i���i�ߏZ�ZQ]�Ú�w�(7U'��c�L��̺|2�����T���{���ޣo�\�~ήړO�ʣ�;��u ��Ea	��ڲ5\�Ь�OXf�w߷���P�#�'�"���#��?�����)�ٽ�g������4�3!w^'�G���M7�+�b�m|t���%�V
B_�'�<�w^�g�~đ9�j<}�_q�t#��˹��$����pdj>�n6��zu�D��\�&�N�E�w�!"�wOii�_h�4�|kI1b���M�)�p呴�h;wu�@�زI���i�7�7	�.`e��u_/_{!��[&��21w�lk�2Η���`��v�-��3Nhѧ>�[8���,r��7��P攰��V�GN�T=ì����K�8�Ϧ���D�Ps([�"��,ү�����s��� (�Ŭ�l8�Z#� �Ūh>�Ha 4Y�Ų2mf�n��g��i��kϖ�^��_7_��zS���C��I��;���ʺ!���Ѳ��_-�N�g��>�NLO��OR���p����E�ˈ�M@ثI���:�:WN�yEwGC{ܸS������f`i藶�	IcgJ[Ӓ~KԦ�u��r��XE.�(���0Ǎb�mq~��� h���"|a����8J���.���(g�QlHA<���g5�t��X�'��s}z9oU�'Y�n�x�h�Z�9��"��1�RW�oE�=gJ��o���a�Lљ�j�ȯpl#qB#��7�^�t��^��Yiv�U_���
v����_Kh���� E^��JR�6'�>�h�M��9uH��s������Qs��Wp��]3lx=�g��g���FS�Αg�o�Y��&�����gt� ⩖?g�6O}�O��X/�E�|E\���¦�,�$�C��[��IhC*���9r���c"��!p-�6X_�ozt��� �x߰W�����#�]�B7CA��8>^ӯ�����^ ��. ��r��ZӬBUp�rg������5a�	Sx���4�WH� �U|�!�}2��	�5P���rN?p�R(y�
Fir[*�~M����.�n+ p][ƃ1���Q@��E����N �U���bڕ����_�x���[���8ezI&�ʲ�z�M���X�ȪY"Q�־x�d�����m��_|�i�_f�?��_Q<�c$9q�Ws#�R�BV���}�΍&��O抠UuM&�^Ei��"�l��D��
2}�%��5��|�.bm	%1,�$c���4X�9�6,rӁ׈{!�ڂ�` ���[�"�b>�`���ɒ'	���A�\���&��@�J��ý?fO�Q�y�����>Gա�F��>ZP�#i-�Gz��,^��V5�2�P���be�.��!�iՙl��M��Zx��f�P�hSV{:U�a�:4��b<J<�X\tz��S�t@��Ө:l��b�|��t��������yh�.�E���{sgjɚ=w�j�}Z��$-��?��Z�B�AM�.�Ft����A#�J�tQ�6��t��!5˂�"ԗK�Ug��'%
*�3O�e�����YU�*�AR|�'Ɉ���V%����Ƈ�[�[(�_u�S�t�����l*�+616�ƴ�Rt>�>����l\�m�D�Dݤv�������=��j�ܱT������D�NW���L�4k\ޘ0y�[@\/����������]���D�o�*_��Ⱥ��2F?fv��K�zlM>r.Q�����n��Z���cޯ'�N�ص�U��F�%8f,�6,��y�AhB&��%�prќ������bO�4� u���#���G�*$-�h�ϔD[w��pJ����?���q��L��Wj�o���L[�?o)�\����#�3f�p8��2cϐ�4�%���s�,&T�"��ykq�<�9p�)�1�w��T}�&�� �����-�� ���!���λ��}G����c<�{���ń����oxV2�Ҟ�0d�����>Z6�xZ!6'��u������K�N�>�S�E؊�BJ�C���JQ|p�'�'���Zm���|�Ӑg{�L�s��m<�ەM�CAR|���k,��������#����7��˩����w'�PW�����wl�9���ɦ;iUd'DY��U����s��x�C@�>��������8���}J|�3��+o�^��RC���՚�ɋ���l�Eh�M��O4�Ć�O�#���}`b��J��o�(��wٓ"Bp�H�A���:����܉;�X�/�i�ه=wL�Z?���x���3#WG�?X$�ΰ��D�&+kzl��R���M��i=�=��(�];^�LK��iۚSJ�� � �N�=���זwݐ�������x)˥$��� ��H��B��D2�iNo�"a����jh�#.%�ܧ��6r�H�[�sg��,^)��BG5��~������\��|��b0L���Ab r��5�EAT�E}d�{��=l�i{�7���i+�m���U�sb�N'���� �	� ��(ҁk�'�X�&Z�z�%��%�z�9Oɻ]��(���Ⓦ&}t�BhS-�^߆�\�:!��yŻ>���$<{DM5R�R��O�]�1���-����7$[H���k�v�˘NA޽�-/z��$�B��&g��6�d@�^/W��` ��)�0��û�z�i2~U�MDI��q�yqoii.C��:����l���ݤs�K�N4+~zV;q�g��U��C��N����/��B�<�wջ�z�'H���d�V����p���}� �44�����6X���7�$L3C) �e�\�����Z;~��`���U�tx6���>�0d����4��d������&l�ڞz��o�(��%�������JR�J�7~d9R�-���*���wO_�C�D|:ۺ)���C���L�J���Ifǧ��M��Ũ�����qX�i2B��ї���0�CKxn�dT[ْ�7��\d����w����ڶŎt�����Y�"ӂ>=��j�O?�L��Pl@�
�zQ�^�O�]"ٶ�	oX	�ygi���>�B�3@���E���g�^�"Ym�����g�w�m�U,F���Z�g��$I��3T�N^`a��!�Oψ
�E�,�+�5��dP�3��k�����B9l�('H�����å��
|�Dq� ud�BbM+�"{����Xo�-�1v�r�mX��}g/�\�trP����|�V�GH<�o���e��Q���ՇF��"S�푂(��{���7��;��i�G����fH��%,E���q9z ��9_,���gY�<�rC�O��H�_�:�=��Ç���%���@�wwS�^j�&�䧡�F,�D����v��}%'h�?�8@g������T�rf�Y���S06��:
��}�� �NW�c@���˵=���+�ikn��6���I?���i��P�h�.�t�P�W����F9�E����Jp\���n��2~�����߳ċ
�x2s���'u�)�8�=�Ih�f,�P	+�c�8#��B`�h�̼kg�B�-T@�K^�Z�}�����o�i�m|Iץ�&���|F}ct���m|w:��H�%�5��1�@�f�C"j���ך9w:
p8R�w3����?�<54�ڐd�hx�c�� y��d7,s�5N`�*p�{!?��|!�������y9zz./���&���ϕD�䞽��vi7� �NN��K BH{�$y󛵘WQ'f������T�=��&,n�Ȥ{x~�R�g0e(��I i�3�F�)WS��f��F� ���|`?)!�[(K���){��_�j`�dP.�E���QD��_��q ��!��\�`[d�{�L&C3�9/������b���l�9
l"Jd~�FmG���㘐��YE��-b1{j�a�Q�"���f`�[e����)�2�5k�������b�p�CY��H�4���滷d���ɥ࡟	�����u'9}V��];�/��KX��*��iOV�u�#���2u�%�YZ�ð(�P��s��=?h��2� ��v8![��H�mN���[�?Í8�w�<஬=�C-8�~�L��o{D��C�V7�,q�!�oʹ�fd���w���pؗ;� ݁U� ��p� �n�YBGe~���r}*��؎�{���KN��a��o}��6�S\�Gt�v ��� ��г�f�+]���x.���rLHstN�>���,[45�Jڶ�3ǟZ>u�s&U�C�^����]���G=���'�E�t��v�m����ny6��?:º
Ը������Z$R3D��H�kA,�c�֏���� ~}��i���WIF���3�s*Q�<�^�i(�V?']SW7�\����������qS,*VyB+M���*w�13S���� ��2i��GZ2��"1��S�6��QO�K�E1�-%�C�~����������X���������\��m�U�#D޴�d��z7b�32ݔT���7�r� Qj��Za�k���&H����4%ǭ��tܗ��-꘶m'�z�i A;�L7�����ԛ���Ь����=�WЩAH�����y߼��L�\����9�c�ga�O!B��;n���$��b��7M��hk��(��V����&{�#����)���'g[C�(h��ŧ�Z"� @s��l����z�U�Ȥa�w�"F}�qͬ��"�d���̑��l
O�b�OU<��U��/U��Q���8��Y�Ϝv,i{��6A��>�󒁘�+F�*V��
��8���A8p��3����3Zyw
4�,m|���Zت�>�.X�gB�h��~���h#x�%M��\�&g����3L�_���������s9�����-'>��*�5���"Ȃ_KR:QQ��`��?Ld���B�<b}n߯�VDA� U�~eux�{��]�#܀/�Nm��煮�]��]�����
K9�z��H9�+��̏�
�W��6l��juqy���JS@��n 4�ho���L��YɸQ���\��X�b/]���H<g�y��1��������P�hb�7@CM%�[�I� �g*�>?����˦Tb5�[���7XE%�Q��[�A�a�2ЧŲ *��;��,�6��Ecq���4�"�ݱ��eϲF�����^�~�܏��4�l���V,�P߽+EY�_4QG�4��Uͮ��HQ�4��Ƌ�V�m�</�����ɜ-�3|�GȤ���P¤���U���u8�s�_1�!�	�������
T�F��B���:�H�S
�:�5�����Z�AH��41I%E��N
��6�偗Iz �r�9�)\��x��ߪV���Ȋo��n4�v�7�OJC��b����!��KTa)0aN��`�t~��E:���%Bm��\��&q��̨��n���I�����W�ǌ�^�׏AOj�z�`/�D2��r��zl����;,���5�-�\o+ځ��(k̛��r{�F�sb-�#1����֑���7�D����8#��VhW���4!�`�p��0�d�
o�x*=�O>20j���]?��ƃ(��=o�������m�F����Ց*?�)�H���sg�>)f!8��V2W��J���`K��.A�u	�~�"�PW��g�T-Y���"1u9	�Ν�٩�;Ϫ��y�_�gv��v�`F^��o��<��3�̛�x�ڗ�]�y��Pc����D/��(��g�J�F�S�dV�[:L]�� ��}i���k�ʣ����3��l���$��� ����6*���v?o�������5��U��Q�z�M��ֹ������x�
?��Хpl4������Uj�/�r���dd��Q�M���Ok���P\�����1t�Syo�¬y{���YQ�^��C�hSTs����X�Ґ�暨bE�t�NI�����[B긥��9�xVQ��q��H��n�"�m��R?W�)n-��tǕ.�㿰�o7�S���k�G�1X�b��ė�ug�k�90tF+�ˬ��{���N���lZu��=���:����[���J�u
�������Fi5�q0$V���n	1�5�(T��z2FA��h�j�A�Dg �6�^�,���]�靧^��g�����g~�>NJG^��nA��ɢ��U|�V(z����}�7J}F�`��1H��U�DJ�|����A������O��8Q7]Y�=�n�n�l_ޠ�p<��wt�Jf9yOJ�����W�.�e��4�� 8��
�+�~��<����j��aV���u�Ԓ�f���}�>�f-��X�I5�0�g�K����.	y鸩��Ϛ�aJ�S�]�[N4�M��1��yz�QI��qP��k�uǗDJ($�sv�h{{ҟ���������R[-�27�o�4�8t�>��*��]�Gn�l)=[�.H"�=�4A"\�e��W]�4�����|+1���UtvV�ɝ� ��~��i�ω:�h���p�e�9m�<���ß�٥�B3���r
�G�&fM�ؑ�_+l�Ə�Η��Sd�N���v�B� ��ow�q��;�id�Hb�>]iA�h����O·�AZ(gCK61n R��wht��+Q���8/3��5��gb!����42j]��Z.�`�t�էF�����)1��+'�G�B�&���X���;`X�=5�(����5����[Sb%�#��1�������H�����aWf�2�k���C�G��3X��5�A���-@/_��!XBv��z����IJ֋x�Ҏ�/��;U6A���쑳���;��lj ݦ�3X�^Z2�x�HXB�B\���=�_^����?A�ă�;[t�ֽ�&�V)س@�]�}�%g�I��nn���Ӽ���`fIp��98���M���ȧA��2`ant�c ��r�	{G:��Y��I�挒�tR��Fl�ct�<|Ug�v����;=D�\ƲP�����t�
i����k���@���4�u|�|��@Se�$�<�<C�KI�����4t�B���<���PG����&b��$?{&L�}m,f�Aq�ݖ��K�:�"Y.�dk�b�?�D2/�����1S��破�A�ߩVwθ���Р����� 3qLDε*|%x_�Z C��$��6�a��?��0Wy���洟���5fX��KZ�����]sa�4Z^��5��3���\��4�6�a���� ߸ؔh+un`��z��\t�M��Fֲ�+�����1y!�	d�f�w)������ZY���Q�ϙ<���v�/=��Mv��f�ْ�~P)kr��m�W`J��.�ձ�l-�'��+c��O�W���jQ8�De�C~�� F������
v���S��氟�뱜��t5�]���A����~���`��o(����^M�[���JF�!���ֵ�̫H�i#�q� {|�@Q�o���'�O'd���)�_�(I����!q8د���J�w�N3 1�z���	~����Ty�luV$!�ntd�vl�&�����Kµ�/�y (�}��(R�G�jr$�	B�������5lX�Tc)Ͻf�fzZ�`
���Ij�j� ��mϓG=�8>j�ʯJ@��>��K�P]���"g�4�?*��)�S\S�~2	A��N>� ��3zv�oWǩ��C��>����!�}��Xn1�o � ��*�4!"�&�e�C�rH�X0�C�nB���1Ѹ���~{�/� ���&��3�� �Gd���o1M��c���1�E#�3E��iY���f8��f��Io�%ߏ��*���d|�b����� ��>���^8�S���PG�0_�ⲟ��X���U}+���z��xc�j����$�u�:���d9�.����$��h ��ieo��4�1GTQ���Dֱ��%"_j������+������+���bZk^�(���\�۰���Y'
�BK��T�d��[��MZ�Zw����bC��'�,����i�f��%��SQ�9��f��]O��*�gp&뛦��W�;��?�F��O�}m�l6�ߪ���ZT���g�=?� ȵ�t�?��gK�3��G"@�
$>�}�Eo ��-y�������w*1-�5�e#�Dl�(����Rǘh��T�s�&����ض�}<��1Vv\:�_�I���%�a��U��~�Y�F�����A����t�[˞��q���>�-�{�[�K̨�:1=��@^�]���.��F9^ϴ۵ �0�)L�f�t�@N7MS{����\�y���;b�����%?L'��eI�bB��QL��o�)Z��,&�
4;�1Z�(hD?
[3*}f"Ͼ�_uT!�ة�����8K�op j4������ғ>а�7�ʺ(1�O�?��yvn˳�uy��d�OQ
��gW�gJ�kv�-��tY��r�J][Q?F�s�w��2���'�Z�
L��G)
k����9��O��LWo$��6�;�n����}����,����W������2��R|�lW���]ļW��>��({x�L�t[��,�,��ԓ^��Yg��ɽ�7�c�	Q�����B`���4h�b�;����������%g1v\��-㿽�c%Ub���6(�k�����#hВ�\3��N^�s5�"�����bw�H� g���o1�V�,ѓ>���z%CǦ,BN��`��&�u�z<�-ƣ�������@t_�l���п8��.��/�34��$*� ��{@)z�T�?FB��]���ِ�^�4�evH�[|4Nm��wJ^��o[�|�8��G�����vuV=  ��U幛s����y������wxˇ"�@�N?#�tZ+M��hT\ŀ�d��H��o9$N��;�i�Qf�S����B���ôz�,��|fJF߽R�CV]]�{�]�5��y�M�#�S�;�����F\�Rp���%H�ֱ�[�^���&�����?rt��Q��8�:ګ1Q1�K�����[0>�e�.p\�r�R���]0ON��)U� %�xw5��Pܔ:���ǌ�� �܂��i��Wv̱Q"��v`��fK�7�ً
���1X�<����H������a�b��R-�}����gH����D��5�a�����咈�M��}��GҠ�HB�#5{�4�B������
w�d�0`�@7�[�\��|�4���Ȥ�K��,Z)�	6ע�� wn��?�}�*�	�z!��f��>S��+h<K���$N����v m��ji��Ҁ�_-"ke���'7�z�T\Igv�h��0 玥Z)��F7�ij.і���x ̒�"�E��p/!�&H�&���c}��'#��E^ݹ�#��fbdC�5�}�M���R}�S�1�&x��q��������S��а-|�R�D;*7߮���l�'���NFѵ\ �$����l�9;\פS�&.��dX̨@��^�?�v`v���Pv?��O�U:�-���{������+[��W��$�uܒ�+]H�y�u��i�X����?���;#q>��{�\���|���lZ���	�a�)����5À ��N�<Y��;%*9��m��"���)\O6�pfu��\�H\�aI.��\jK��=Y�g�H@���u���=��b�j�ԍ�d[%0�)eK{�Ƽ�����e0����0˦��a? jI*O�FE��ҁ������),�p`��,/m�Xw❰Ce�����CR��]��~��	����4ġR[6O�ي����ʙ�p6��-�R�ښ�n�ʐ�C��G�on�c��������q�P�R���p�oKk%@"��m�P��
��n� ������O�lJ��%f��N�n�"�Yp3��UT�*b�> ���_���#�)��W��]�TD�O/�D�9�3��,?�ҋ��F�k��Ql?���A3|�ȝ��q�d@�;�yzl������U��[nb�R�	h��n�m���#��¨ޏs�{��	����a�Phv�ô��+�M�x�Lb��4�#���)dM���gj�Z|}*�cz�R�Wʢ�[�_I �sr����f�Ӄ�AV4?E&�s�*��8�}�&d	��ɗ�[q��x�������@<'�2�G��|������|
�RP��p�=s��.�Eԯ���[�{qJ`c8��AtE��&��N�~���ݩ��Z�� d)<C��`
��YU?�s��P�0<�u?�W�_t}g��Xa��P��$��#[��H��ѺBɧ�-�: �R0��J�sx�`�70ɭ�R�{��i��3�;W��
�b����1�Y��AF�F�tK�\%B�um/C%�(�����^?w>���(r��%���m*�s@Y +M���������
Y`�8ʋ�F�����Z��6�Đ�c�gC����;��{��v���Q:ɯ[�$�n ���8eZT���'���Fw�xq���&$�8q�nbL*B�:�^V�,a�/.��ˊ$l��O�m�|�SY�O��&AE��1cU�<���f]�/S��QU^�$��=��S¹4�'۴U�bZf;q���_��y����[�PK������˾���ߏ�t˼���}D�&Ul�'���6��P"H����J��Q�-��G�L�{h#.Zd�޶�P��Q�(A��x:�EH	|��
o�aZ��q��r6���4�a�f�[z���Z�7�m�`�]&S	�[qk
�=Ih1ڑ�1�5UA�0?_?����KEX�twҲb�A"�1k+��d��{Ty��EO�<%�Y��<6N�a�:cG�4��ڹA�)X��t��Jhx�k��꽾�<�>���%7�>Q]����̒�rm�O�},U�KIH�����|L<�!��>d��8Z�����[�Я��:��Q�ŏ	��hj��x�-{Ug�[n^%ÍUΟ�NKal��@<o���-7Ri�6c�����?��ʹ�/;�"_`:U�_�Q�O!�n�u�I���� |�|�� �1�(SEJ_Ip��7\�GSa��`u���A��'~r�>Q~.�p�`���y��AO��?������7�&����[��X� ��TC�I��kb��d��5?e/��r�32��l2��Þ~|�7Xru��n �>WP/�Ob@HH��X��j�$�m�}{�x��L�1��,e�zH�l�=s<6Y_�w{b�65�X����*>Q/_�]Kɲ��#5���ڋ^�;��j�|�%Ϋ���u��©�Y�`� �E9��b��aƐ>z��n*fc��@�V�WS��(��\��U Xi1w���x}!THO�v�x��|��8�ƪ��E�a�3
K�M6)WQԿ;�Y��x=�Gd���z�����<�}�Q8Е��R�,�A�Q��GV���k@��>�v��qo@e(k�������v)ҿ{��fo؍¡eT=�ug�͊z��WG��"0�n�s��:��E���2y��ɻD��w�à���+"KCX�f��~���HAHܮ4������$5��υ8�@1�J�ҕ�I��8JZC���M���=�`��,�4�D���={��޽�2MQs����~�����d@���sT7Ye�����������&��4�6j=�I��vrڡ~����g�d���]x|-3�,�~��T��h�/Z!��֗��8�-�(L�_� b�%�8.w:�o�M��-������s�j�#����
3�������c�]Մ�]_�����ҩ� ���Yi"�:���t����Y������#���q���S�m��Zy*`Ƽщ�����g
�n�Zw��	���!�G��S��?!z��kIV���蘸l����7�s����n�'O)B\��*Ґ(�3�i��|��ݒ6 ��H$�$1�����#f�O�o��N�g�G�C��ʯ�)������l�׷a뛥|Ƃk��ٚJ0|
}.������1�v������U`�)V��qK�ӗJ]�JK��i�}�,���j���O�O{�θ��+�|�]& �������x]-��B�F��Mh��n�Z��ь�ky���Q
|� �T`u���'�;��2�1�V�c��&\;}Ȉ��E7|"��CU�/uz5Z=���Ȳצ�"3�@}ͬ^�z��qr9@˶��L�-�����wǼ��A�<it��E��"M6gu�����;.���|�V���C����rq3��F%ԉ�&��sw�vd��e�E�LS��P����P����e�l&:�x���isF��~�pe)O�7m����%����x辤�5�{���8�����-5���8�Ϧ��;BՈ�|�(�K� {��:�*{\����
��>)	��C��H ��U��U��!d���H=�&+-���Kն��hp�G��sƩł�	���f:��h�F⺈U_��X���SSnv\d������Oo�0l�ڒ}緩�s1���j`(8y�K����Ϩq��!x
��ܱ�A��ЕEk7(�lJE�ʾ�Bs�G���Gx c��N�̠��zٗ6?Ė�5s��da���%�����F�:I��G)~�[%H͵��ۉ������t�� F��o#;7�
�p;rt1�f�s�q�;�gڰ���> 1�]?oV�{�A>)�;��(�Y�����K��Ms�R�]B�d+�c���\d�즨NjB���|BSf�Y����?��x��bXRj�D�K���!��0(��ፖ,u�x�؅�� rrel�Ww_ex���4s\�{�S�>1����5�M�����m!6�O�#3
�ch�Q�e���~\Fk������\7�z��R|�����5�ۺ�w�^"^�8�C]��q{�Mf��.wd�����\�,��e�n��%��8�79:��J&Ziޠ}O�U��	��vRhV� TI���껄M����a@��<�~����с�6|��y{޼DM��`;�$�P�	-���H��;�+i��Y�d;H԰�[��(q�"��->_�Z��C^�Ysp���0�x�j�7��a9V}��rH���O�ԙG�ݏ���,6������	,�;��+,]�-Í(@&W����9�ߟ������G��\��n�]�p��Z�:IKxm���}�輤��/]��i�ka��9�� 5گ1��$W�����a~$��}�mHOt��`�<"�?sS�o�fR�60z���m=��D�E��7��S��8���P��ϫ�_�On^z�|�H�(IA�c��"G��ww��$al��+���;��\��	�s{imͳ��� � �&�N~����_�7�d�������!ʲ��e��|�?�P�	�R��i���53���.9�P������쓒a'�6�3�yf�O�~��tk���� O�iބ�5�����������	����F��8�pn9(�yb�[i�""�ߩ��#�<^\r0�9±�����#$M��H����I>)+"�8^��.U�҆��'z'�FAi�/Xt�`��J=��ً���-�t�M�^̚�y;`��U(���ݚ՘�!ͻ����l�p(
,�;����_�J;dG�s���Qj�p���0�JZ�y��ذ�P
�� ��uO;_�k!X;���4�KW���
Qr��t�l͍�=�\�f��d;�?Ԇ�v�Fg�+�%0����q-���6�tc2}�Q�&���(#����'?W�z�80a֤����?�U�}Ŧ`yQ�㼱. �Tj�{��A����|fM~�n���*���'��� N�!�hJY��X4�?h���ˉ��oV��$�A�y�v����;s��c�ktB؟im_)��M�����KMx���=���.���T��>l#(��B� i�@��j_^����n�RI��� =�?&��Q>;����~�U1��~�Nv���B���}k��69�)��hkw=3��Z���B��^�w8c,q*�>�$F�{<�_��d�d?ls4��U��	�6��x��-�\�D�yN��>.�g��#�P��n�����|����ù��"~I�i&��a�S�9�VL�5��N�x��sA`�trE�4�Z��������!#,��aSܦ�e[-�-�K�+企�%����[�T��Y��*���*���PMF�,�HW��E�H�L?D'`p:��Y�'��A,a Z�?.p�?z���
.:��"O����pHp9cN?�a�I9n��s����o�w����3W�؏�A�ڷ�� MF,��&�16�����{�ꑶ����� ��d� @��:��M�&���jcJM5������Z�*��"\7�Sz��$g|n˜�jۘA��"x�O��AM�E�ܠ��)T�]�����dWH7J<��14G��^3"�[����3
�ʓ�tS�d� e��ӂ��������q8��HdC=� �����*8DI�i�����}[5v�d�6�,�U�N���Wm��B���+�0N����|r}l�=1�'�砜x���Ed(
��`�κ��p1W�#��N�����>���o5�IX����m �\YN-ɂ�H&���Bk��� ����R
�����K�e/ ʧ��0�0���Ϥ��S*G%r<�$��
.�7L�Y�G#�T�#�.��k�ݚzr�,�����Ǔ����'n_�]&��w@��|k���+��tu�����ٍ�s�e?���t�r�����(ur���K��3�u��5�c�k ;��Z(���4]��0�hgVJ�=-O᱐�x*�U��x3P�6�M�22>�P�=|\?� �4يwV`9�����^�����'ŀ�T焛W���9]m�Ҙe�t��-�p���M�X�\��\��p8\#�"�N�|G�@�XW�R5�#M���'"��Vd�D;L�G�����X�^[�VtZ[4����:�������8SzJ�X��J6��|����:�V�5�"�Z-�7f{���a���Q�nf���L��������u�t2jd�ǻI�d=�e�y��7ĺT�v�`�'�^~�)]��[˵y���6��7b���֋����=`��9�,X��v�|k��!��E,�����\��z�tr��­�f6帗#������-�ܷ`w㬫Y�f>|i�r1��iv�������,�K�r}�p;�Mu���G��ԁ���"���?���+;f$�k���3�4<v>�����͝������b�H�I�_H7m_O�����_2�f�ˆ��#�~�������K�S�C�ҋAM	ssę\����!=�%��b= ۇ�!5��" e��a���]�y�]� u�'3�Am��$.�ZƎ�9��M��6+����;q0HRbj%8�{��h��=^�·����E9���b�o*��(
�Q�~xw<�N��a_Gغ�Q+! $�"���~~�"�Z;�;��r���R}4��Z̓be��XyL' ��Wlh�mU�WK�kFCŞa��u�%����NއuJ�2�ծU4���-u��^::�笲�K�߭Q^�bu쳍�҇?zRZA�S#q��癘��o�o]"~q�+��Ɖ�|o�S|l��soCN�:�ASj�8S�	����#le1\&�w��
�y��Iw�4ֵ�XG�ǗyMx��7����}�d��	3d00���Ar�$�r�rL>���P/"�z�Xl�Sx�Z]k#Pi��~�mP�9�V���p8����u�kGu�XWR���x�'[A���"$Qw��/�d���W����=��2>M+��liR ��(��0�M�~i�!#E#���������^�n"��9·��������Eg�x��kH��̒Ua�5��, �_�V��
A<����%�GJމY�t��ucř�n��B
�/����#�2m,r��%4&���ʳ����~%r���_�v��� ���;oǅ�8`\�M��<�&a6f��V:�X��=zs�
�����,�oye�5��+;�?p�n��e���0�
F��2V|���.¬f7��)���맍gڼj-6�:�d����Z��j[ Xh��_��7�����5���KJ�>�}�T���0�!�����;6���H|Rʟ�X������Yz�y{�C_`� �~��I�{��|�ʻ�%�$�ʫ�qY���C�Q[�d_�x�!
�� a����2���\�T7-j�/�\�<VDr)�%"$K�T>`Y���_�
�c����s�څݕ`�f�]��oS�p���~u6u��l�v������)�X0^�t�	����ߴ�#�U:|�5~f�",-�ƪQ/B@oh=�#����Fž@���VGA�%��t!L�ݷ��ũ����%ն�(Gɝgp�ŖNNT��^�J[9�h�)��7E~E����� �^�Q�+��^ȍ�~�9dV=ԚJ�q+fq�7)x��k�!rj?���'���`|�^�]������"Ή�2|6H&3�>��6�r��8GS���&�����f�F�-�yl<�5�xFUl ����%��)�̉D�1�8����{��t�6k�������o�}�,)x�/����'hV0_*���	0�A�F%�8�?:uW���j�m���Li�8�W��C�%�R��_�W��aǬR1������iG�S ��7~��1FAq��H=[��Hj����p�4i"�l�瞄9�}���*Ɍp:�����WѮ���؈ὴ�|�/�Ղ�ANF^�L��@6ii�M?��i]���Rk�0�t
o�z�5��!�s�v��#��l���
�R�4���ٰS�Q�(��'2*��M�Z�3?,�1����Ȧ���dfN�֠F�� ��v2%1�.}z��S(��v��5R�*����;Ht�;���\�xC&�kKKܪ���?�g��7����$����),MhM�^���|�i>�wHcHD���W�!i�ԁ��AY�j0����H��h�miՍ(�˵�:�8N�a�i�A�5�1 �\��-*"|����v���o6��D�L�G�hn�.6�]ڃEI��,����H�o+˰l�T�����{%O-����Q�T�Զ��{�Ī1=��9p�L.�wM�/z.�\<��!�:�\�iu���-�W�SCT[?B
�')ޛ{p@�4�������
�<��"�Z��X��gL�@۾a�d#Ef�'���Q�V�N�{�)Ba�tx�ϥ&�Ag*fqg�y�e����YbC-��rݖ�
���.k2�B̆(w���{B�Fi��b`�S-����p^��6W`�/�{��� ���{)��<���c~�.r5��&u���F�5Vg
rR�[�#��t�����ݷ�!�B���{K���qa��*0r�m�rϮ̣$���%��`,E��鵔�2�<�d����c�L	�u��^�R���vX!�mκ/~q$��4����=���G:T�y�&:��-O+T��p[��/5�=�wd.I
�����^�pKf�=c,5ݒi%�	�E$��1��kS%I��q��ǆ4��֎�>`�H ��uՔV)c�E���`��Mm֜�����[�W�A�A�'Qf>Z@<����/�/aEh�l�)HT� �լA&�%<�h6��)�+@��]n���-�ʂ)?�«|��Ҵ	�q���-wR(/���I��L�acOq<XC�;^ ��띵��d����(�(0�C}E��A��"��G2h�ar_7>�$p��RBP�'�)���;J�i��Y�M���~8���5�w
���s��ͮ��[�����Ƌ+�J��kS���0����	#
S<u猅1�}���~��yP�$�O��1Շ��#���zR�R��)
f�Q��ݙD/�G[XZn��.x�N#�P����΄a�@�=�*�PmK\�EѠ�&�@(�Z��:l��'P)�4�푨�|'|���P���GH��i��
�a��~"���jɘt��zڵW��&v����9��/S=��������J�&�
�ҐV�C��+~B�X��[�����`�,�`�W�񶥮n]����,�A�!s�n���1$� һ��[ �����q�nZ�^M륽�,�Z�)w�kj�:�u��I~��5��[oap:¿zJ8ԙ󻶅o��+�VB%k�Ә����	��thU�'�q�x�9��TiX�����]Y��[�l�wH�V.���w.ܭgT�:a��U��D1~?�VJ�-�n�_��N2�y�ڻ>0LE;clݵ����ڝYNOM�`������O����F���f���J<�JY�<�Yr�"/�sN��~��i���sw�6f$���J	4C.�(��sRk�=�S�^^�U���<-6��)Z�P��{���~l�An���̛os+��툩����K�屒=�F�0�/�������}�'v/�~դ�,�c>6n27^ub"V����}蔟���UZ�EcЇ��cʈjo�C�P��ؚ�5�kr��x$���LU��f̞����8�;]�a�����K��v�]�DG?��\?�N��2{G���v���Y�.# %�Y���K�mN�Mr�up�u0G��)��[܅�����Ns�o��ZO�� h��	�*�.�B��{���" ��6��/@�ƍb��%}��?vO_��`H_Q0N
�H�R������;�X�P~���%Ѧ=~� C�)ic4�r-��R'�0'!��sV]�����᪂U����h�T�W/�G�mҷ<���{�EJ��) j�b����
Y�'��,��P'��}�~�2>�*��J�c;q�)22*�f�ϤdQp$���twƕ����:C����gL�ekt��*@B>�ofW�g&�$RǓ�>�6סTJCO�W�*��sq�YGz]���3��O����[k���M1��di��G��M!��r�ßS"Z�7�!:y'�+���x�V�N�5��'@Up�JE�4���<n����}��{�$O����ߢ��O�;��83J֬��r�w��y�;j�5��~9u	�d1̱��/�x���9�S!�^�죯���q���q�`4�oF��T���� �xk����TD.xd@�gϸ��+=� ��]&)8� ~��%=|/�3>$x��6�0I�+{~�6Z��7hmBH����+2��h0)�Fx�*��e[KU�̉�4�Y����3�t>d�6f�;��2�.�ٺ�P��P��[�GBka��y�zLxg�yh��Z���	��E�Z��j1m�EV�z,Y�Bϖ|��͋Pm�۷�XuyvŘŁ.
�E���4VPY�DD�l�T�x=�;��4oSD��sq|�J�0���͓S�*��@LѾI�AN����c�93^S%g��%�54�n�J��	xS�m�o�2|�u��/5�W	��8�2�]H��C;_0�k�0���3pF�{�2��z�89��X�"��j��Eg��^l�3�x���l���(2Rx��xٲo�� �<��&�zl�BȞB���� �� L�THP��T��<�@���z�	�0�����MkN��A޼J`�x���s
)���z���=�2��	â�,��y3'����RT�C�h��!�@O�vek}�!��(F�E����u��N�Z�I�I�t^`��<hhi�}7�I'z�]Q�zf�d=0���L��Ǔ6�(�)R<7@EsVr%��`O�L�<*&V�����9��|�Zdx�&��'���3|5�ώ>���r�Y���3C��߁f�0-����Lكbж�����,�h=�7�/ _6.�3�X?Y��� �F�LT�V�}��e��������@dY�m�$��2�(w��	pQś���k�\��B��/�L�P7z.��I{Gb_b�R-J����`צ����?��vf�a�gl���:k�"S�n�h頷�PվD�����������

i�c|�חF�[����QB�a���kk�[{�q��3��"\Y�Y�{~Lj��@H�����2�sv]��N�A�+�F��`8�~�F~�D#�Į�x#�^�=\8y�#^K4�A.e~�cu�4���$m�W�F�S1��"�BӉ#�a��R\LzW�(8b���6#�ٳ���B1к�%�L�f�{r�� 3p������j(UH���'Ƀ ����9�uDa�. �;u�����&�F���<�^�sՀ%ݿ�+n�oV�+�.j�M�\��,�g�-*���&��N�]���A�]�We[��D��s��ɲ�Ub���^%�r�\DGYr��&�7W��V2��
1�^~h @�g7���d�?G�n�6�!��δ�+����I�%\Vɀ������%�	�l����d�5�`��.� �>=4vQ �(9
��A������٤T��w7&����~�Tܝf �BI�/����{�+�"�B���K�Qq�ֳx��?�"��fY3¢�e����S�w�7���q����	���1��qg�t������ɿ�.
Z���O��8tP;�ߣMD-��B\��6���S1����Ŷ�c&��bU��^ǌ_�Bg���`�f�!W��}oF����c���uJ�PhP���jwK�p|���F�;�3)�|�ϊ�\���`/G��$�Ł�6ꙟ�دu.��H�[�ܵ�_��3�t<���&�(��_l�E�5}��bʍ�E�ږL��-�QX�TRBa�ahv�?��Y�ӊ�A�"�#[>�S���ik�YmL=Y5Q�;�E��=�?Ye6�T|Lz�([ڃ:D1�?�B4����	���<�$�-#�����}�Z��ЅK��N���x�;��W%B.\0y�i�5
Ut��P��L5Ю�-�R�;�7��/�U>�g������>���Oϕ�ܗ��]��q�yu���?֫�fI��鑐¦��"u]h����3I�F�1\C1s��������o�e�YB�?h�f��X(xe^V,��]�9-�/չ���s?��QGb_���^qI�eM!�pL��f�`Q��\	��'i��?�yHXy�i�g�YJmG�m�ӟ��[Q5\��3_�
nc0��V~6�f�L'�ۊ/���i�0xf3柸(t��<w�E���%HY�F�.������ᗈ��XN7w�]�	�ו+	�Q���o7�J��D1���D���z������(�?k!��p�搦���{��e�l�YBC=��)	Ĭ�jJ�e5~��3K�K���N��eV�M����׿v#A��*\�o�	�cP�p&�Ff=8�&q#�Gв2��,��J$K\W>.��ק2,
���=FL�$�Z�����`oE}G�է �Bi~�Z�O!Q��,�h���-x�u�w�7�Qq^��ƻ��Yiάآ���x�����J�<c)��r��f6�*ج�ӀmsB*��usP��F�S*n3Ɏ/�d�>f=G8�1�'�����Gix�O�AQ�uF��d�u�kQ 6Z�hA�t��`�������U��^�pe�9���2{L|��$+y��%hߘPty�Ц���>Ŕ9���E0��(��<�N9;����7����!�ERd����aP�Qv�Q��N����^u1�oRO i�5��؄��ǘ��Kvl�|H𡑠f�D��p8�|���,>b���Fg����};�`�v������rzl%�?[_�#��q�B M	F�G����S�iE;�ߧO�+�V���h�1H�W�m]�y�1���!�(3�A8�mC	���
l�A���"t�Iɪd��g���_�0ބ->墾ק��l!�47K��}	��i����vQ[�V[�[�( ��e��w�>yӧ��.����e���E8/5ϧ\*����^��R�j����쨗�Ý�-M2hy���ud�����B}�8̌=贼�5��k!��rv$矒8;���
Ul��'E`�L��&p(��j�LcDo3��Hs"i��p0H�3���ֈy0a�LQP��IK>���j��$Z����ȝP�o�I����:/S�	pF"�L���=�b&b'��]�'�G��oyZy��y�m�����G�,�������&�W&����*k��ϩqw�w8?�$�,���;�
��f�8[Pk;����o����O��#v`ݣ:�,�R4��|��Dfx:�s��k~"��m3�@`N"��3�x��D-���+;��o�B#�p����'V9z_��"�q1�9w ��R��%�q������w������k�-H��ad������u��Jպ��l`�S�)�"��t>�C�3S���n�@��q �\�Rl�������G�B�����Yn��L�=x����>B�C�2G�J�A�8�9J�����Y�~}�0ZĢ�
�U�$���u��d���WX0�`+�����Px+��Qx�S�|0���}���h�6.J�I�m�@�����X/=M~O��6f���²���]t��LO�N���Cr^�t�p�F3����}��,�z�4
��HM�#P���Q-��z����4F���.A�ogy�)?˫Z�Ҹ�����s$n�(P�a�|�t�*�x�-_�Lv�9�Ykm���������E��]����ȇ+�¦��W�x���*'�χI����c:1pL���GՋ2e�O$c�Bq����Ĝ:s�Z��^���u tB0�ʶWR�ԵM@�L^��Y~�������#Xo(rR#��d����n-�;`�k-�^��M\�_q�oA�[8�|��n��}�@��&���;���)hF:XX�8?OAS�S���
�J��.S� �M|�p� �je��Y8������:+TkJ�5��y�[��H��Y�b u�
�N�&��(���lw��4�F���@oBN<��^�W�@���ʮ�0*�}�!�#�!���I�u�[�>�,#�!$$�.Y��zÅȵx�5��mw"���mE^=�μ��~`�9�0�52��I��`�k)�U(������(�:~�G����R�|�ݹ�8֖���|�ڃ\1�,��
�D�;��=��cm�)��0w�9�H7�Ёm	r=���	����x���C��o��䇳
ϭJB�g�`������DNܠ$�y�v�Z��ǖ��i�ѩ�Q�4��|��f~^q3/���e/b5�s������=����r���W2�#>q���PA�E�@l�݇eEr�\n˳Rw�����aQ�����a#�\� }Z�c7�\CF�q����<IY��]Q�	�,�l�r(d�Rͥ/��鰚��:�*��Fz��^���-&��(�y�>���'��y��5q֝�j��I�\G:BI��
8��mg ��ץ��&���A��q�,t����t��m��B����Հ�2<0()?�V3��ݨ׼A�D�;߲w�k�m)�(���0%|l!]�ӣ�|{��;ct^��\��6�'W�E�W�Z�<7�x`�֪�J��QX6,����ލ~
����|��0�es�(���Y��Vъi[r	]���yz]��*5]n��*�r�Su�Q&�E�J>��a�YAI'��@o v(��Zv����:���ϋP�����,[j�A��� z�U|�=x����!���g� �OD���+����r.E8�C^��y��6���W�o�/��
mns5�sݑ�L�i�ygg��+���N�+��Ϋ����WL3�Y()��?��w�>��%���|P�kOq����?�$����
#5K�n�n�Ue����[`����=M*�>ö�֍���@���j�Ä��#����6�gJ0�J`�����3.7||:��cJw �R/$8� �`��y��$j�Xg>j���><�0������H��*`$�<K��e��~��Y�R7r9O�|��'�����\t�͟8�#�`���hXn%��#����=���v�z������ȼ�.!E�~��S/[U���qC~ |+bxD�M�@�wA�P�C�n:�i �5+���d2"F*�t�I0�:lW�Z��v��q�A|��X֞��eg}5_��D��	A@���.D^~9��6��\Qz�-��2NX\ ���t��Q�[(��2A��������أ�-�í�&���1�WeTd���B�&��|b��LҢ8�G�����Je�M��0z�=NXWw�����/#D<�;�۔���q��뜪��;?���_�?a46~�^��҈�w[D���k�ؑ+"�oH)_L+G�L~e�n��&�������.Td��j$���e}�Vc8�I�h	��f�(�ұ��R/5:�U7���P�iib�Hq�Y�α�?\73\Qk�K��WrV��7?#"]�S-ϟ}���Q�����$�Ln�N?���D(����=(/Fm�`��̆�iq=R��]����W��m��	�Ҷ��n��E`���t2���wH�gŹdTub�C�V�Xܕ����ц�&��Z���V���l���y@�Y�	������Ѽ�j/��m�B}�6Bz�����l��*�r���0c8{��uB��`�I2:�,g�Y�V�и�s~3���/�8L�q?�%T�蛮(j_t��I޾4n��A�D������w0�]�Z�]�S�T�]r�fp����뷯����GJ�����}�q�Ԏ]����ڴh��Req�&!�<q:�R&���x�U�N����\�m�H���c� �����P���s�����4�k��t�_��lyI���5�����A�	W�}�Ljw��l��VU��H�uy��W�(n�!��^�[5P�R�� g���ޮ���^@�ʁ�+�8��"�C�Ԛ������]� ��+����0}]78�}�	��3�c�S��@u���HV�U��.�����?y]4S�_lW16�����s�I��C���~��7��4���f@�CIY��Fy�)ǡ��1F
��ezZ+7Pr.�ݐ)�������*2�ѥ�|m���DV�>�)H��G֯���S1vW����i�51��uDq2>9�g��9A*�%��a!�߷,� }� �<�H��M��r�%p��c�ojX�n��C?���L7k����S?~�8���c����h 5�s s��i����ĥ#t��N.���q`��ܫ7Tc�֟����^�fZ�ݏL�LZ%�_��h����P��=�p�������*>>��T"Ɔ�9EY��I��7���t3�>^ٳ�mw����K@��T��g�u�r9uIe�c�łXH)����G@ԩ%0��Ͷ,�WP�'����̭8��Z�t�1��f�Gdܵբ�'�N��p�K���Q���Pܝ��M�iL9!k\t�!r`��CO�Uw�H'�� �L+RZZPD��BL�&�%�R ��N�T������B�3>!{���5;N�똑y�S��m]d]ǯjO�:}�֬��ri�0>���j`/��pC����g Z\Xz�5	|��m��Y0owNm�$С�>y�4j�x[���%K8:B��nb��w�1'� /��⿉��Ę.g��J\�]��N}���$\rD� N�;��6����r�.ֽ��H�DAָ�%�rbRi��釭S�gt��$�xXǓD�a5��"b5O�#�Y�}����j��L��1c$
��`�_;\�x.oL���2i'�{�i�����������Nz�D�=2N�B�w��+��.�d�C�A�:��oY��-i�@�[�hD�hO�2zzF���7�F/=��; �٪d�6e^=��MR�����6'gk���|��$��l{BK�WʮC�(��WF���E?��X7r��u��d�Wx��e��Q� �����8�Rwz�s�@�^s�^��5�gUB^�$>���;�%zh)�����k3U� `(��-���Ǻ�*	.�p6p���3�Zf���y^��(��/֬|�mf�8��p����|����	L��/�i�d�pz�tBd��`�[��Q���>o�eD1��v��;��t���;˒�+h�Lv
!l�/e�g
�ׄZ���5�UN�����tp���ȓb�)��IR�9`�敷��f�E���N_a�ǐܯ��z���fS)f����W��o�^b�By��4E���}�c�M��O�ӬD����;أ�'��gb�:��A2[ �Y�#���S�,�>�f�-p�Lƕ*J��5՞�ѯ+y ���� �Jn�|����zx����myx	R�*����p&&���^���GɈe�R*�%��z_)�s(����/�"ٙ�ϰ�ڞ�K��/)�����x��ȟ|���!���	�j�t�C�Y�s_h�J��w�/���(�h��(6�P�0�L�ԋ�7)(�0 �n�8�s�6��+�Z	�<&{�a$�s?Pb;�V6�aD�S
'%���,%�sCa�Zo,����\�`���=/xjj�v�q�d:�2��A&l?�j�2�1t��F:������,?? ;�躓��޾�C��p*��g`�~��]FޢWxaؕ�t�!�2���b�dFq�����p�y25�V�9�}��'ڟd��XpcY�xk����k_��� ���%���V�K�RHf=�wա�R�5��W>�$A�_n�z����x�����%���*r/�+������ؐ�:=r~��)M��U�'BJn趎�-͆�As~���&ȎR�"(fl�XW�7~~��2r,��t���PST�(�(�C�gs��=;���wť�֜�
n*f��?g���vc��ɱ�)�أ\�t"�'f(u`�_Z���_�'D��� ������┦�����a=%�w��4�N�z��4G��d�E!�V�f� ��� ^gzN[⼤U�>3+q�nF�HNج���"�1M�{������J.�.��_u�*���9ǀ(�6��[0��gi�xi��G�Y;��U�S��O7f����֬i�G�fs���h�̂�"cd �[����!��
��Xr�-���@Ì�Ol�zأ�`�Gف�t�����;��aL����ڣ�����
������B7m2�ޱ�ӳ�m�����Ͳq_p�q��jZVo:VmO���q��{�/8I�~u���S��4K	{��R��9��9jW�aӅ���hď شp�~�/���3h�e�Y>�O7���f^y����a~�o���G���|[���co)oE��ћi%z�Ա��d���*�tb�f*C����)�%B��L�xT|$g�sI�#���'�~�m�,��������ҧ�k���%X��r�w�S��;�9ˮ�f	d��9:�҉���ٲN�G=)]�����u�H�U�qga���T��o�V��Bi�M�&_r`[C?6��R7!m���{6��g���l�Ua4��ܢ���~��v�:�ʊ����a��)|4z�/��o��g#�?˯��C���N(l<��rCb���K�}뺅Pfsy��]�,���_�w뚓d�� ��S<6rx��8����Fړ{l.xi;�ҥz�9B��q#C�6�0�xΔ)��M+xo��8����L^ϥ�z������/ɧߖ&i���RC�ͤ��U�S=�B�5��i��~>h���o�Z*��a��4��HlR�&wY���V$�7��|������Y�����q�x���.��N����Mu��l�X�m��P��Ά���R���E̳9��C�<mw��Ug����#�DB����ɓ�=5�>^r�U`�m�=k�Ӈв�xy�i�A�]��b��f��/sn���v�yi���_鎬S�s��ΥU��,
�Ѿ�58T̹џʶ?�3ޥAJ���,��Dot@��^СA�H�%�E��v9Q)�<��/�<>C���K��5�ٴ���-��� l�qD'Q��
\v�(Ȕ	��c���K��[�jx�N���D7 �h��d�OHVL�<Sl�yѧr|t!&�^V�������G���c�z)��;B8���/��,#(a��$�E�%헃{)��̌'F��L�:�~�6�h���7��Z���oIa�+���H���d�2>��$b��7"g�'���V8��]~����ʕ�<�z��sT6@�}y����
����s2F�J� �d��|�)�����2
�[�p�]h��$����8~��]D���n]�p"����z�KE�.^�b��KҶ���^�bIr�G���U�a��p�^�k�)G�*��{�YF.	�Ȭb�Z;�
�}�O|�pfΒ���dЌfS�����@��oB
�p�G�r4ئj"�`~N��#�7#������<��{��q)"D�A��7�PTu�Q_���.\Mu�����%Wj[�X�����J��t�k��BJ4�S�}��Ig"pL�>i��1%�S�4��;�`���2�b�R��zb;��2#5�_�u�?r��'��"̩��l�;#ܮ�-2�[�(x�ͤ�p�������v`͝ꚨ���󃱿�_��Q�{��Z�yV&x�|�}��@�4v���
��4�� Weδ�M�?�&�T	�@nn�/��0���SD�p@_�����M_H����m�Ol��~m/���_n���H� O���1���+��!��F>^:j��c.sW��Ѱw�6g���Qk�`z�;\���n,6�����X\ҖM$�By�s���1��K�y�~�Z�#� ��MjA^1)���NS+W�'3�I`��@����� F�*X|>7�dW�C�n�[��-1�D���mBs��W�H����5�J���휟r��9��-<.nS?��['+w�uoRE�`WMD�+ä�x�³2��t�����/^��b���Y�L��E�f�����9-��A�LxPW��[X��Rء��%�$h��$���1�[L����^O��� �t���M��jhf[�sfR���	��c��P�Ĺ �:O�	�$a��ș �f���Mw���Q�)X)�R%_jX��*f�5�>�� �y5�b������=�$.�R;�`V:�J2'/K�E&yo�Tjy �u@u),�99u�v��o;C�� �:�j>[���SŹka�����(�>���bϱ� �R�4e��]kT��+�|&���"H��n�e��O�Oc_*�S�-D����ܭ8�����x���aXmÁh���^ţB���ؖ�[\�!죡��DeY���C\�P>���q����0V�e��ku1�V�����ѩs* �ss��Z�\%�	r��[P����-؄Hh��jUPa�ˤ ��j�A*@A��;\�e�N�	{��L8I㓃:��\!�e-���b@$`�Tw��������<�FMymw�����ș�vą����4σךS�4��}T�2��FsTF�"b�A�����k�R�ۄ��Q
+�@������3k��S��.)�{�,�w��zDZrr";Q����l~�gT'�T���r��|�$L"L���I��G31i��V#��W�V.�P�@[����r�%C\��уA�-{�=c��E��E�5��7���s����:�,b,��C�"��)X��(��c8�/4��L}�_�p'C�"@խ`G*�O}���Z5Q�L�)z�����/px��Hhվ�=�k$�pU>H�A[����jW�ޑ���t6��Ǿ	aO��[�5cٳ�d!&X��k?�����8�_G��(��u��S���it��X�ʪR3�D1䇹���:;ޏe6��\��BPd_[��D�Iς�%<"!�������lZC�r5����:�:�0%~y�8�T@B0 ?Y}@��Hz�#׼����T�hO��?m�}aH8�V�Q�>���pK<7w���]Gw�Srvs�v&	��+���3��w����X�9��s���k�
�(%n�!l�E��;�B*��U�� |���be���<��8��ɏ�"�-K�~���$��٢Ba�-|k���^:q��="�2��l���-�EJϭeX��'���]�G*�3��O�%��R�˷С�2:��Q�&b�O)Դ���FM��h�Ʊ�J�@Y��a�@d�g�C��S#*�-\:�_Y�ASY�����3k�.�yx�ۻ*����
 /M�� ��?w���k�ƶg�>ퟜ�6�Y�Y��r�����mQF�)s�ҿ�hNb��b戰qTr�Ƨ�~i��mH�X�:�!
��)�A��	>�N�h�`t�4o��V�_����f��U�?�P�SL,@�F*<��_��[αn
���a�|�=���)�F����Hz,
�!�^HEn}��l_�6�w���@��`}���� F=���'=	�њ .��[}� ��g��M �HB|���H@�驄���_�7^�`�o���I��qѯ]��v��^��a
U������3 �~qD��*[E[��}���&����}�׭��(�r�U�P�Ji�9e����0UkpC�O�@8D]�9�s�'K��@
k�{]���`�L��/������__�=�"��U1�W|Ҙ������D-�����w5y������@= �Ey��rPS!lV__����mqs�mx2�|rj�g��4�3ҍD���?��¿E�)��4Ȉ*m��t���[y�*y�'M�T!�i�4��B�F*��C䎅�z�$�C��Hu����֐Ҡ?�m����q�Zj���fW��ג��Mo{������v&�Ǥ�c��1�_qY��FMiY�Naz�'�~,��ѷI8f��(T��:�y2L��0J�V`^m2	kY�� DJ�_�X�;F�zl&��7�^X9�.�tvy� �{"q�s�U���.��&i�<U�'�_�ut��~*�����%Wof�=@���u)G�֝����φ�!�Iv�y�%�`�`&�ɘ���%�7Ev�p��ًFC�+|wq���k�+�N�I��0��������【\��\b��L\�L�Nj>Up.X��DuQdJ�3��8��&��������j���d���@
:�!��uh06��_���]���੺�ʯ���������\�eM�W�2X�\z�ۑ�}�P��.��M�E~v���Kgkӝ�turT^�>N�e'�.!�wzo�}6d�����=�}+'9V���w�3�K�uI����!�me�#U���6�p��;��-Y�;,�7ihPe����n�֣/����Cu�s��jS�Ѩ�D��,	j�]b�:p�zN>�.30�/����:c�C��l�m'�:4X��K� �O��Ȟ���S-~�[?68�Q�'�)Y;9�VN�ZA
0گ VO�_#F-ȿ���4�qB�>�	k�>�W�h�����}&���(��l�ǒ�fm���lO�i5(s����^2��}�$U����MP
oj'��) ����U�y^��W�6�EX�a�|���)� ���5��&A��S���S��*��8nh��}Gg�SH\@������