��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&�O�}>Yo���>s��d�������a<4s�^ae���r��(e�ſ����h��ҍ~yP�3��T��ڃ�ך^Rڿ��2��Eu�Z�lfL����[K����c.�����x�H���3�0����*�dm�M%�')��"������GM�`�"X�Ḅ?a�}5Ha4��� S�^/�Ru�R�b���q<S��T�w�Rfs -�ﴇ1-� 
,���G�z�"�a/��?��
�@M���p1K�&�3�,���q<��j&#�9���(�� ��}�{�Zn��f�}��B��<���06s�T��=_�"Dz�]�s(��O� �I�����R�3��I�E�pOȜ@�$��s����L��`�� �*zKS!W��	(��MP�Տc�kvs���_�oS@mi�"\����%g���k�S�%�Q��A/�"�ij�s����q��@�r�(�1dz���w�톁��=�\���?� �Z����Ł�Bz=��.����.���O���eZ��W to�;1��X}����||vu��`������F���3.Um�	��Lo���">���F�p'�HK�@Lai���6'��=�ci�����}���Ț�)�� �� ��=�=i����EA��$;�y����q7�?�p������(�n�~�.�v��0�n���j�"��5�n���q���(.���urqUٌ��T��]�Eֿ�74a���9u+�P`��� ��1��{ ��3��q�/���Q���d8ۏ�,��^W |�����\z�3FgQrd &&H�6���E�:ř�	���b��v^��?�"���p�aq����bx��n�8��i�i޳�_,-��+�~�4�.M�`�9T�r�
:v���Q�hr�ܟ@�l�Wsh\9�Ƅ�$�z(����t{:V�RG[�x\��1~���|�t�Z�zZ����jD��k�Ӓ�q�(�l�P��o?I׎��2O��I���m�B:���Uh��o$�l*�u��@�pRCF�Zɧ$~����m�r'�0],���AT��� ��k�(s�u� "Q�>9��ZLh�F�Q�t_�g���7*���D�F�\����^��D�F��<{p��c��C��]F�n߃D8���)�Yɵ�ak �*-XP�30�<����Wͧ�[��΀}m�)���_��S��$���@:Y�S���*#�u��3���ķH�y|�s�U�ʻ�ك��O���4�4kO��/���p�r��ǬW�i�������X�K]��,^W���M&t���� i����B����M�X��zW�s~��dm�iM4]�2�mV��L�1^WԨ 1�����\�#4�>�rC�d@���H��-�V�_�M�x7t=>d�&���_C��I<pqpS�)����_��TK��4v@*ʜ�n�%��̇n��1�g.�k��˂lW��М&�W��3|O1#@��93���8������Z��0����b�]RgO��|��ܳ ��l%��΀�a���\~��v'{��A1����W���<��!��}�f��D\��R!W�ED�A�����ij�b(fi�/�\+?Ύ�-��RaH%)�7�	���փ��o����U���L�BgQl�_>��W�8�3�f�,�_��۩����(�a�eV7��<F��*�ݳ��"��Ŀ�m�������8��;#�#��d�SZ���S�Y3���.���z�J��	��QÉd[�B�[X�P02Z^DjJ!�(�����I�lV��\7���8"Qt�0%|+�w�:@�a)J0����bmV&��O�8(���H��C�滛�	*�4�N�2& �6�yU���q�`V|�*�%#�q���4(�_�ߧ�Y�ͪ����5�Y��(>��̬�#\y��K5At���wW�Z��vfd�R�A!�;����M�I����%����T#�ǡ���P���Ʃ6��a����@�M�������941rH�[sQ��ķH��F�qtӬN59zN	�f��䩘�@��A�k���TX�L�k��x(�T�B�PK4O��P7�����W�E��

�ZM�d'�C>80�A�j'����|�,��I��x������)��3�CO6��Y�����ɛN�i�@h\DZc����!:�X�O���v���(�D|W�����8q�IdH�ҭ�z���v��Q��ӱw�)�y!���������J:�I?�9&��X��I}�&L�
����%�?������b嘏�Q[�I�n
/8�� ��Y�J�Ri�����e��y&1d��~���l�%��� �
�U�{-����� Vނ[�]#�+B72�	��d"�F��a�4�6T_���9P@��p,�D����Bc�D�fG���{I�H7p��8��dY�
�`ы��I�h_�@����k�>��9!��V�g��2�������,�zu_K��V�ψ`�[\��V.X��i�2��&
�?M	Tz�Q�y����)��OzDrS�y�uT�_�E2��k#-�-zV1b���H�@:�h#�v_��n `V�� � e\)��hᖆ�ѸH�:M(.5�}L�����������A�H������?����{�-�֡aSX���ьZ����}�;3���L���c�#+k�"��+�Y���o��X��k'}0�+��Ys1��V�ҍM�~�E*���q��O���rת�- �v��-��M\N���g����Arf�MS<"�{��sN�@�{.4G^����ǒ[Fj-̅��p��ͣ7g��� M�Wߜ�%�W��e�J�9w�Be�!���s0�׭t� D�����������'#���"��x���p��ٕ$�l(OFL���M�:ċWZ�Q�Rc12�	��ˁ�l���&D�Z V0Io�yڎU1�L�aF���`A�LAZ8��0$�O��_�d�f������QA�t��O@��l��~	N\���/�H̬`��i����WN&(�oj���l0$���<���V'M��L�/��B�U��.� 4�<&kh�f$���΋�']�$G��\)����lg4���+���hzx����m��Vv=���+>��Dn��j����^�`~���"*�u�B&,
�S�	� �x��<�}/<$H���T&���]�K��)If�D�~at:vټ�0|����B�څ��2ǭ���րPq��F��e�ú'�����NjN�g0R������]C�W�$��%*�����f��������T�����n�fp�*魝?[���3kT���ryt$�c�s�tI�G��HHE:}/��]ta��a�0�����և����,�� ���o �|��*n%Q��9EC^0��:��<�Y�e���������gbiq������Mt&�w����EgB70�tId�K�RLiVẃ�HF�nm{.�a�Q�x���ΫK��GA�2�^�NB2-�m�����t�]��t�\��r�W֑�bQ�2�[,k>(����]�tV�/=P&r[$9�<��[���/y��|����tu�z�\l)��Ar0]pZA����>5�0g)�����!V�(���)����J��
�oM��7�i�o�G�'�i9��r0��!ɢ훅_t�ʹQ��5�]�gF�[�E��ψ��D
�n�0!ԕ���~�Ԫ|/8(�7�8I��}L��1q�:�������۹�Y����2��?��z�����vD30�X�I>����z��S#���A}t��y�_���6��/h�J����J��2��]d_�.��޸��G`��p��8��0���"��(7\i�Ⰵ���hT��n��-~4�ٞ�����oW-��P�sb�qOI%]�r3���sC���ؘ�k �%]1��G����wк�>����!ĩ����=�DU0OLp_�9��52��#����N�q�N��H�"��O��T����'�wl��|~4��r�|�-˶o�!��{������U�/��J~!�* $����3����--y�7�ؓ<U�٠�|,���;�g����{>�����0�����&���`����d�*��9�jJ�Q�Sb��b�S�bU����2��#��Y�.��NE����ڴe��`"�d ��e��ޟ/�F(���d���3x�C��T�"0K������x�gS2�V涯7���ƕE�Y-hޝqkc1-�^>��+c*��h���8��Y�41:���6�}ON�-Z�?_��5E4S��	l�����H���͘��Wæg2B�ǷYκ���lMb��s��xڬM|1�ԣg`�yW�a��b��zZ��2t@��U��/Jde֣{�y�B{���[����y����~"xD����l��[A�{����/t����~�� K�mgyf�����ھ"g��rLWP�����Sa.����OG`����x��[�U��a�T6R �L�m��/Z㹈�"��rӲAϼ"|����$-��E�C��*G�.ѓ�H%`���@��W��>׍�.ϧr�#����Adp��B�����=���Aֱ5xr�^(�h�6NK(2.�m��m�2��Z�1�cu��_��~`��pi1_F73�)�+V�流�)%�w�)PX�_f�on��x衠�x�M��R<�b�?���?�s��mȀ#��:^�돻v��M��F'�{������q�Ɨ�q�إw���+˗`'q7�L�̀�Ĉ��\�2����f�ޟ*�C?��N��*��-N���R��ةX��`� ��/��zsc�~��87�G�2�9�͗���*̢�u0�9��Տ���q2��A�f�� Հ���*��Z���%��2��PB[/rJ�h1�Y-�i�0ps����.<�����	۴r��c$g���eӱ����ώ�F�5���fs�e#�a}���*�K��}(@X7�U��o7f�ߚo�,�15~�p�i���k?�6 ��I�>�d�uEv���%M"6��F�� ����̍5,�ﯫ��m����Gp	�7
��ӑ@L�/-[��aV�g`J Bh�_���(�B���߬��>\�~�5��J�V=�Z�&ݨ�7Q�w��$����$���9��,�?��(5;!��T��*}C�}[&nP�\eo�����
���Gʉ+3�V7��
�2�낣�@�*���ڰ�(���=���u�K�Q� m�pr7r���	��z9�=�|T3�C�[s��?��FG��CZ�3���Sg����Axº���̂�0�O�qBE�q��d��\<��r*���v��ڕ�9N��������2I�3$D��� t%�1>�d���<���=��������� ���9�o�`��|�������?_�`>I-��wi���X��\ ����ʎ�7UI�����ʆ~����(�ǟ�,)3���N�#�#��U��^�;z6�����Iiɳ����/�!�n�#�T��^�a����N������l�A�Y@���v��R�N��V�d��L�^ݳ��g�#�s=fcD<6�\��[��H���)��?y=�ii��FMNbߗ0�l��O&_)YK�+n=����sw�EY
-��]ښ{��@┸P�e��`�_n9��1^��6GK���F��;x�7�='�rg�&qO�@{- ��3󜃥O�������P��i�eM�j �}S髞{��B�Ϳ�MA'���[&�N��*5��ol5�d������)����v��r��;�j��5:��Hʟj?��1�a���d�N_���5_����D�1*���m ����,�ů�f�F����߿�	/��@���"�;f��[��et����6�}n�(j� �0���6� ��k\��\���e(휛[�([�3�_���9��1J�$j�ǟ���G��T�g�z{���T��G'ّ��J��CEU���s��6��7�N�C�Å1/F��&ƿ\�@���Q3�����yH���+�3RQ~�Jb�K�r����8@U]w>�ZA�yS�fg%�P�-(�!��;�/�Vع���ȰӇ���j���j?HA|r%uR̃���3?,>�T��+䜅qN4��xOp�ȿ�%^�!BE�^�9-l�`te�{e�6_��uG�o̹�����l��V[?�S"8���Tk���L�ʡ�=���+ϱV�U��F�e�e��d�����o6�ûdcP��.�A�=�3��Bi����3K�A�w�p�%c\o�I)�K������+��?ĵ�Ƈ�q���|��w'��U��I]�\�S���""�鲬Wu�/����0���~��5��Bݰ�pqq]�AgS�'̦c&'�Av��m���a
�H�}֥�h
�u_*���[Ӕ�~��*�]�n.R;�4�6Zz�����Q��v��&4�Y����i�����mϣ���'���a:q�$I����+X?�T�F�:4�����J�D������ÿq-��0 nF��.��|�R0��kW� =�R=�+�Í#��e�KsTV�C��������..�r�u����q�'eS���b��§���E�	�T��L\�aq�d+���]�V�>��$A$���9ǎ+.��0��bW�&�_9{���?��m��V2�.fǌ}� ���hv���z��d%�2���G1�?pפ�c�ןUn)U�1@��"��a���z�26he��!4� >�a�dpc��5 ���jR�O�ˡ[������	Z���̐�O��\f�oBڳ|�lj�z�7����Q��֔�dS�_ɢ2$@�<yi����v`+0�5�O�`�g��i!��>R x�� �����G:
�m�sz
�l�ݫ@Jec��c��xJj�y��F�RS���b��c�����4�u�[{�G��5�6�z�y�������wu�{�''2�j�L#4��׊�H��v�˼�^�4-���>�����8-	Qs���<I� l�*!mqB)�7�E]L�`.�XJB�+*��������aM&0{ށgn/;���^�4h �Y�G�Uwu`�S���ŨJ�ȬیG��u��օj�R&`������@!�X��XO%�x=Y��f�}k�����A�=�����=0F���C�����_�,~�O��� I,����#��49A��&A�xp�����_j���y���|���+h;�����ձ�W$41�-�����~\P��K��Pi�&"|�[\J~v�N���)�@�@�z�+JA�������γ !�|�|�8B�J�b�����-	���tD��˟�2�6+�z�.���{��vԳf�����5����ñ��R�Hj�BX�,}
Zx�g��8��iډ�2���H��w�k�f/Vsz��;lR�^��<�x%Q�a�H����g��͟S6P_6���BE?�HF�	���,V�x���B�l[)p�%�?�gf���bux�� �<���觪x�ͻ�vs�����lu�_�K�BvW��� ����Y�>�D�\�t;^cS�{)K�L:"+P}R�fȾ�J%���%U�8$����78��Hs㡟�i&�hyN�=�y�b�oabO�[���$��4�x�_#�{�SM�
�)ہ����J�P��#�_2�����V�j����^��	
UDgPǚ���@^~�bu����dL�b�R�5l�u�����`�E�3���յt>-�n�7�G�h��2��+^�*�$��q5��k@�Z!ժ����j�+�B7�dBB�|��nڍg�Es��RU�850w�����vw;DeH��3��2�6�NE	{�q��u��WE�+��tc8YP�輓�s�������f����S�dM�>z�;~�"pPL"eP�P�r�J�S�D�g�&��N�H��L�}�"g�2�L0Ǆn��DQsf��ɡ��tXx|�i�Ͷ�l1��]3ԥde;�v��^a����g��!4�-Fn�n��ȄK��䟞p,ؠ�i<|�_A6Q��1�e7�j�7�>�r;�����{>�鞏��lF-��F�S49h�"���G����"pN%���U�Ӟ�Fۂּ�`��F�I�r�fe��3I-��3�i���V�'��O�U��u8��.�]y}vC����M�|�UFM�ʗ��GgOc��@�LI4T{jI72
Q�T�I�q�Q6~k~��1�@��;H?��×4��!�AJ�T֍�ҍa��_���C�+���/>s���ȸ	��
y{n7V`W�:��<�+��e~{���ґ�?q&��t������Γ�>��@�k��RL�[o�!rQѯK������e���n=\~����9�se�|�m������n
�%�`	5�7U��Z�� }��*��5g�x�Q#���Ar#�W���HJ�����3��T2WzQY$�a�/�S�1iҰ�VM��� ��Y2��.�3�V�L�S?�V\�F����	�?y��m�~9=�����V�;�ǳ�lT���t�a��D�Q��ﱨ��Y��[��J&��B'�SM�ҽʤf"	Ǧ9�ˊ�!�Z�:�=*����z(��2���	-�)��Q�y�;Ѓ��}�z�>O/�֤�R�eRDx�w6�;�^һ����9H�3�o�%K�g�/��2Uo���S�߰��y�M��R��^��tV�},�쀍[�Z	0���^[΀N�Ш��F��*���L�%������qf���N��:�d���Z��,*�9pg��!����X���_�˱�;*L������rdkܧj/��ƴ
f�!���"Y�w}�b��� ��T�6�vi�-`x��!�C��\M2�~8(U���|koϩ����.M[c�Fd�m�䣒̽��n�W'�Q�}��>ޖl�_�AX�̺��,(�ۼ%���1K>G�R����c�[f�Lʖl�S�Br�p�r�c���ʞ`�`J ��T��բ��D'QÖk����x�T�$�I�?�l��&#���L,O����K���Ͽ�A�3��T��kC���M�����0�hE�^�#��y�o1�
�	�ew�,�d�?|5�U����O�&��צωB1�XTrƯ��ʼ���R�Ը�o�)~�0*$��~���s�?��W&���k8嫛,��}�
�@��[�3���Sk��bi��[��,�F�"~��2�ud��F�h��sx�(���N����7��9/0o8@�"*�~�ۍ��!z���,���ѯ~��j �Ey�g�S��?�5+�s(�K�H|���(�j�2�]�'� ����>g����%��HJ��F�06s3	�cl�DV�f��Ud� 	w�k��H�g���ю��y�#Uߘ�}w�'��`ϖ�O�	��''^���V�Q�YW�FA�
H����)5Zj��{��$3L�A�6��Mճ`G�S�l�o+��@�~n��U��Ƴ��^zc�
�J;m�-H�y�n��`�����J	��?4Io~j`��{����������X���n�U ��U���\�������ƇM0����C�ٛT�x�^"s���0ϰ���&�|�e`�'���4(崜�eg���1�)�<�,���{���n�`�]�Y2w��,|ŀ��;�P
� �����o@�$�<"t�_:P/9Y� 7ȝoON:=���!B�	
o��XX�l?V����
���SQ���j�!T��+�wH�� �/Ͼ���<��+��E�b���X7�9�Ry�N�WN�)����0�&<�K����/CN���������v��In��1��?g�,ٌ)��4���0�m�#�T����e3��&5+�C%�.D�yA��#G(�F�x�u�V!2"R�+��'aP4�A�s@e�H1	��XC��{8U��e!�>-�7�n�f��U�\
�0�&��3��.���遞�v,��6s�N
Ҡ����+_r8K%�A�+,�9���~�!�%��.��"��4T�ͭ����h�aƀ+>��¨��[#@YL���?v�����]�`���iLEX�ty�n!�$�C�? ��	��J�q���͠u̾�J��Jez�.�e�\��YDd��h�P�ˎc���-��5D*7�h���p .!�P����Qǜl�9�%�f��Zmm�v�ZK�T�B� ���7�.����*�a�)^h�6R�nfh3�;�4�-���W��iE��!tg"6�8�J�|C�6�� �i���F_(d��#0�>������O�5���J �^[��:���E��x��.$�Jk��n9�0��U4,L:>?j��1Z����(®><|�)��P��L w���I�*��8D��!����	�5��K}��{�rq��1����N���wd����,��7޶�D�j�zc�0���0L�_?pa{���Do�X��+�Џ�<C!�l~{=7~+�M-#��y?�1�q_5fC���5a�{�k�r��-y�g��Xe
r�Ar5bڬ;���L�.=�5��ơA���S����8�=7Y:���7n�Q��5��oN;e� ���!V�ZTu-�ݘ�%,�t6Eh���k Ĥ��&os.�-a+�FV�.���鞛!�6���5܎w]���|WS�m��n�f��kh����-�X��n#^f������8'Y�H��<'+�����,��xg���@H!�D����
���lג��] ��Gw���J���P�E̡�B� 	�@��)w�6�OO���=�R^�rծ�� �+�&���7��.����vcI`���KFj�#wh��� 5�*(^�ɮ��8��_�k��6�	�z����k''fS��Pjt��]L��Qb�QZt��X:���h�t'v.R-~S�1@]2��'���ψx�㬍\�E-���0bA��z�ž��"����Ps=k�8��n������[t2�m�L;�0����q6V�)*�HA1���	�7ˣ4:����`�3����;֝����
X���1^əۈ��åE����&4J�c��H����]�u+ed��Q&g�c�x_��$h*,�ey�4�E2��i&j��F�x��_�Y�s��%u���Eq�Ģk�R|�8bn�ך+TH����2>�R0X;�)����GX��ۮ �x�����d]u3��U�Ș�H�f�7�� t��(��8r�ڼ���X���Nl�P-��Wob6!��{����x�Rw$<��A �&r�[�H��u�Oa�.�听�j�%O�W)m�%�e5�H�L7X�7������B �&�^�$�ەXD���v*O���4q1�dguj�hjG��x|�ӊ����+�$���lO��I�f�δ1�$�'�J6PV��	����Gg��N��i��3-.֘����V��k�K8˾:F��Zn��3y����#���qa�v+z�n��MiҺ�	�o� �}"xO��;	�O>�c��E���]�Ĉi.����.5��3�iB�_��
[�����#<�0l�6�PA�%�����U�L-�`�@옙��aa�:�#C�e��9��!\��i�}�_)����<� ��
y�x�5�tYQ�U�.�?���΁�?�S�\���r�~v�$w��g�-�T��<;��h��H�%jO~�L��e�k����g
ak�M��n�����3I�/&i���^�Z�~�� +�.H۬zD̦.'��&!5�B�?@v���AvMC��h;5A��z�Oo	����������g���g���C���އ�Ky�8"�bI3�?�e��柟,K"��Sa���.��O�w2����A1�}�d�)�58 : ������P�v�Ȣ嫎� ����ۃ�-[qw|�k���!���4T�(���y6���^�'j�H�p���e[���)�Ldw"�J�T�s���j`��m�lM���R|<@=�P��lk���jw"�la���E�ۭ$����a��<���
E��X��r��"x�Z1j�����f�\���9��L��B�M��?�U�c[�p�v���_�c|���ef��@���h����8�_cU .k`��Tx�7��r�oi�MW[�a=çJF��Vu90$��W4�:T�7S72_�(.�!|��d�I�/���D��j⳿W":a�A�F6A�"�U���f^߅$®,� |�jOD�M�Dz`4�R1�A��yRA��Y���E���<��L�&?�7O��,�d�Y�j��	��,�Z�j��j�<��4�p�sq���dqҡꙊi�w)~�Yn�_�9o��d�8x�7��vL@�$��" 9����עw>-52�zD�C�7�����x��m5��]��}8�r�����)�4�����C�%"n�^q�cz�f�N�+K4J�Ϝx����&?U�D*)�9*�GIio�}��~u_&W�M�5��X�����C�f�I[ǐ;���ݜ�]C�=�U� A	xU�= m��t=�v�n�
�r��eY��!W�]~�hLӺ���켌�)�Cm��J᪻M;Lc.�֖x����;���u	,��=4�\���u���
��2���(j��S4SA�O���4>sX@E�6����D��[p�Q��q�p��g�ae��W<4�8B[u�J=h	"lnY�e|>:
 ����H|�=��G�%_�..��n#r������0����M�0��;z����:7������}>��+��X_�*�t�5zi�U^�Y-�H�J� ��Y��0D+D���Uu�j�B��A9R��a�Y������Cn�PUph:���*��I�%�l��H@L��MC!��P?;&j�~/8wez���I��6Gm7�$҄�/Z̊;�B����7����;vc�&܇�&>K��*� �I�/8�
WQ�~-��[�R��16ʚx��c�l15�õ�2_���EyV:���I��
�
�c��ɠ��`h�Ntʥ3����Ó��șK�����Xw�:�N�\���B� k�ia, �r2~lg�n-�@
�[ �K�(���,⵰����){��f�u����.T�*JenՅH��!E��&g�?���ޏ_W�f�g�J�G%�	k�j�����H)Y��pJ��U�nv���r:|�%���i!�Ӧ�7���+aRq
�K����sy̐A�tb�@�0��!1@��X�%x�>pE|y1=�O`v7����M��b�tY!߲>_�SiTK?����Y��_�~�S�'�	��35:�(uڝ߮��[b��)�׺M��y|�����`�W��:.��bح����?6� �/���r6
E$_��	��mn� �Ȳi��6'�Gq|Y}~j�0yYƽ�T���L�d3)�ɏ�duZ+lF3���l�@��|�w��d;�A�S�� [7��vqX�E��4A��82!$3�5@�8�"GQ�n��cqr���A�)�Â�k�JmO}�ZJ��Ŋtt��.?WU���3���Eᢾ֦��c1w,Vw8�� ��� E&�raey|��6���f}nC�P�a���&߳���XrWԬ��N�m��� X\T`�����!yID�RX�����mT��˹��;~�~h63���j�Z0k����)��F=��-�6��t��?wɴ�d_ۤ�N����Y�L��[T�h#ȥ�eC"0Nn`��PBc�N뿍��F=O�|l��CY�%�D$	ض�< �M�oW��o�k�����s�!�Y0�����J�RM�#�f�P*���m���%Ep���[K���ѿO�`M.����x�q٦?�栉��-0r��l��\dgJp%�A�oZ�/6	XHg`'���5�Rr{����.�ج��%k�j�DX��0�L�EC�ڄ�\�#��G��f1E��w����4��H���ĆV.]�����j"��iF����n*�Y����ˮ�1Pܥ=\��wS�'=L�QV1���E�p�E��n8n0��jh��l��&�ά8�z�M6C�M>���1����F�\|�Z*��Ѭ�/���H2T�����`q�[y��6��ϮŮ(�ǯ�x�����u���;lB�ґ�<��rҡB��x��KI(�`8�y�\�˾�-�V�`�ڧ*4�)�D�2�&q6���,$ق��ôs�A3��-{�W8#��f���p�B��9���B����Q����9rv�A֑��g�9�1�^��<*�v��b	�4�a/�)4��w�R0&�5�M8h�Gv�pbu�FL��s�|���%���܊k� N;�Z�\m�T�0�3Tq+���}:r qIT˶؉���'�����>�v��`���qvp@}2�� ��^��Q����A�&x
��e�t�ɚ����M���AyC\�u���٩��Ϧ-t!�I��x\d�"�ݢ»p�ZOp�Y���IΉ��|xj����@'����a�p��4|�P}-��3;yeQ�mN|� �Jf���L)%����?ȕ>��Y�H��K���Gɫ˱^]�/[EH��-��+ %��F�y�D�*�g@����ƌ!D,ɮ�I���t�!j�>�O���|6���"�H��F�n�9b(�w��5�Ow)O
�H������KEȒ.p�?A@#\��S����H��x�F� ��(���Ѷ�қ+�N��� �sj|/:eGF�qa����{x�� * ���`t�j���$6���i�k��(䏹ǣ�ҏ�Qq���Q;'L�W�8ЎI��J�O�i@D���j/s��0�����3'K���"�E)��x�z�{2(��OH�04r#�#��`�n��;��QEPt�z	�@�7�� G�u��[?/���K^$�a�lׁ�iƺV\��Q��^�Ѵ�10��r��&�`�I�v�>�(Exx�/��;t;5`�}�x;XK�۵��N-YgG���3S�,�W@��q�^����XE^��ѳ�����Yɑ��^Io�# "L�&���ո�5�9,��0���h�`�X��U#A��_ �!ԺȈk�%=^� ���k�Y��K�~��4�'�s�0w�=[��.Ώ�)
G8��mJ�a$τ���7=�F�:�B�1��5����Ƞ�J-�hd����K�>�����p�k��p�X�%Wi3*5��ʉ��Ä)��V���EU���kax��m�Mp��
S(h*��ctA�A`K����V.8���uP��~��X]p ��=���/����6Gv���P�K�U9��D]������g���$���~Vۢ���������&���iط@OtĆ4�b>