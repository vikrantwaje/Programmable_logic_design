��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�������~`�?j#���Oz(�ybת�:X;Q��
Ȝ��V����U���8�D�8��,
[92��y��������Q��aq@1�2p����5��,�g�a���b	 ���5��G��r>��T�CF2cΎ���/�wb�!�~��R������� �1,]�z��q[ }F(V)r�P��X�~nP{o��\��L�o�'���8' r+0\>(z��;k����C�� �u���PE��x',�ٜTW$�WV~Ĝp"�=�F�M��)�]k1�3������g : ����?����+x�_	6)�6�YAw)��!��b�M��7+�L�m_p9�w�BtՃ
"�`�Jr>W;v�ǳ��,��}�#��9�ɜיn��Z��;j�G�$��;k+����jS���3¦��f�������fuAWk�Y�A�uj184�3ev-���j�Z�|}���T��"*��&1c�X;J\��@����Lq��,�i,�_%��[���>�³��n8�;�V����=PTN6!y5����+"[\�%�̗�5m��lT�Yp;�,t��Vxƹ��,�S��y2��v'w�a?�Ә������5;�}hq�=����lE�U���H1��FFs���{]����p������u���o�v�zAT��@	��"��g�DY�g;A��I'�Gj4j��	9�?}�L�\^��H�Ks�n�q����/gd�^d�-�]�ۼ���/|�z�-�[�����C|��G���eL�k��,�#�Ы�Ռe��<T<��V��zP�|�7CO�wBm_qϻ#��{&��V�N��<���Q+��vUJ�ŀ�^�Z�>�j;\���V�+kZ�J�M �.󰷐\815��/7�q�`Ʌ�V˰h2S���VCeW�A�4l�s������	�p�I#`��'�`���L��`�@a=]6 (�X�1^=��sr���a)�P@T�]�L֋��$��}j8DE�׹1U,�V��X���љ�x��_q�JPB��)�p$Կ7�r���܋ѯ5�OQ�gF��5�n>��Qy 2�Њ�^C5�+n|�I�̢��٨�L]3�RTC��k�u98C)�q�A�~�U��x:��D�6�A�4y��m�m=��p!��X�W΀��ݶe���c;�R\�����O�Az�m6�tܚK����:U%��n�\���ʼ��Vz��[�p`L�9A�SR�fdxg>�;��7RV��bon�%�T�ț+���%Y�8�~�5A��iv�w��2��4��~s^O��ľK���Xw�'��W�<�ü����*&�M����Vao��#ɑ�%[�*�(�k�7�\rŷ)i�wK�>M�@K_O��K��Eò����S-y�
]�ul3Qc>[�GI3�(g�����2e��x\����%�|z�~t��RÇ���H��cҤ3&�y�q�����
җ��B��Z/ T(������^�����m%���<� o����@UB�������<k>�C콩�X#�@�_K,R��H<"�zf0*k�TH~?�c[_&�
JJ�z����_1�Id�O�.p��ɋ�(�k,�&���n�Z�L�� �����V8�"̒H:A���MNT)�@	K��?���0�����F�������W�X0�s��M��R���� ]hr�0h�S�}�6���Ϋ��Gz� �S�w=}+O5\-��*��N�Y�L����bI������(�ٓ�
��|df<���e��p���=��qVE�(#Uma~�V����e�.���%�W�%�,��N�Z}ps�
�}�Snǉ]���h
���L��"O�0!©	gxՉ-�;%�K/�#@�e`0���>3Y��A���M�Z���3j�˃u�жf���e�����Zg�
C�����6kW�2�o�Ww*֪�^��Mguv=�
�i�g ·8{� x��T�9=e�k:!ppv��}Җl���x����$�"�FR���W��vtMu�V�}��w�ϩK�$0V�����͊Zb8��f-�!�(� �D�U#^���o����8x���vǺ�;걹��#���"�Lf�c��ǔC�x0c����'����U/�
���a*u�h��w��EZO��KIrHǖ�`�C�`E��W0r��L{G�W�^���r��/Gn:����z�x�la����<pˍ)No{= I�(���=�6��M|���������T�g$��<U*��P�S7��0���=׃�eaF�q0��^[��`�'�0$,߆��ѬJ��_�#۫�	WD&�^�4�"L��j�^�D(�s����/��g��qB��h�X�53)�,^��F�.�d���n�S%*�H�`O�c�g�����~-��6<�a�?`���r�=�p�l%��9�Πn.��ܹ"�n�%�k�W�yf!�)x��\�)�Q�DJ����p>Fll�0���W3��we��,�ܘD�u56<Q�sAsb��xN�22&-G8�;���J�ϯͥ�
��ztJ�Y�3�B��s9��^�d��Xljx�ۓA��"/��)�IpQ�.����'�&+���u1*�G�۾��K��s3���v���?�,LJ�1UD�P�+��G��ZO[&�秢kZ޸y����_�#���=iMXj�@�;��gG\�@�B�#�
�AP������i��j]��4����
������2~dU���Z���ͺ���
o�̺*��G���Y4��Sy�)`j�u�}��t:%jO�jxRq6MNQ�H���&��x!��%�4��#A*�0��6vi4z��86,&����:�h���D͑n]� ���(gs����>�P'i����i�7�.���t�L�_�B��˼f���I����,�s�J�y5�KPxm0헶�%�-�発.�ɘ�G�az�����
�ާ{(�7��B�j�κ��o��97O��{���~�.[e8����s6`���x����崙�'(\ǫ���"��LH��D2/Z����*�V��.����s��?$���t���>}�sU���Yd���u(��� /���f��~*W���B���M��|������8�xUo�!�1D�t7�����Q/V�!߾���K�+�N���Ɓ�x"��c3s�����'5�q�36��be��_f�3�M�:
iKmz��G��+�:��ұ<Q�߃$$Q��sy c�~y�C;
�rU�7В�}�X�.-�@���e_����t�h#a᩾��B��%�	p�Y�	��]򌔋���[)���~)��Ԍ:�G�^R|4�Vё��8=��O�#�4�I;������׌*�z@�dl�,h�Rރ��"T�8���N؞m˙z�?���*� �߆k�)0���p5��P�j��]X6:hM�%Y#CCQ	0U(D2Ly�b[��#@��/�;.�^�p���q<u���4�8�u��(߽5�}�W/���G�l�礓���<5����թ�v��]��B�<��=�m���	��t�=؃b�)����'�u(<%3T=�\SH)����[e]��Ҽ%U�w?p8 X���W"���F!ܻ1/PDk6��
7���Ӂr�d,H|�Fđ�J��$��]�Y�IA�ĺ#g��^Ak�|�{�3��Ɂ���Z��sX��"� �w}"X!�+3���S����bd�38��o3��(v�<{4�Ouf���Q[X���G���T��;e�D'�]��۫�F����a�P9��,�[�m�0m��<�?�aq��9a�C
���_�R=�!��Iu��
')������~G�N�5��͟�^&�JVZ��چV�]Ȓ�Vm������gV�� I�,?�<dy+�7鼕ia�B���d��N�jp�6��~gf�e��4���-�Z��b��m�6��uH����u��:?�y�.�i����m��N<�o�W"�u)�޿Eѻ�h�qއ�ŚH��ՎGT��Q]�R#j�v��/Ì����f�����p��5������2EȀWG[�PnKP�4T.K�C,hJ���]��\e���� �^���#ިe�[~�)8�R�g�%6ɥ��FSЭ	����/s��9�f��#E��!
��p�[)+���b�h���d�<7O��BB!+��=�F�g�)��=\o��ęT�GR�RKF�h%�4%���W���`�{��%q)�f�3��':N��ZI��ZT>�b����;�v1V����J���W~"�'�w�� ��f�$$�{���/�nX�#,f��"!"R��tz��]���D������ͧ$ث���(4ﺋJ���?౪ ׌�f=(j�p��X����v�m!�!�\�a�������I��.�"������?��§l�)ɟ�\�� H��=��^���;�y�s?��c��J!��ïdĽaI��	.�d�L\�@HQ�d�Z�rO�6+o���P�A�</��u)(WÕ}�Њ��	TC�����a��3���V{��
Jې���_��'�z�C���ZG�f�@7Ι�0n�� h�����K#�KQ��o�,hf,�>hj�����p2.[��}�I{Z��D�������	��J��V0E�3�A4��)����w]�����2����
2$�W&-ԇ��곇��������{t�֒B��jO���L^en�6Y��ʉ,�F6�\U3s�b�H�1(���x�L��G��A�Z�����A�e�Q���O�1Α�Nd��g.�V,I���V,�4*�3��W7���\%�C���t"�b	"���&"#�t$Ϟ�%�z����Ⱥ��0g��^R�2z�`L�|��(t�߷�O�i�����0��u*�p{���H�6�S�T���ៗ�A@'�x�x����'�L��Ѧ�����9;f�,����z����zY����Bzo��%�m��[~y�$���������Z�x�xn?��~��.�EpNKq�itT��9b��!�h�#X/�?v�i+$��d9UڦNB�����]mH����_�z��=�ʃ�ֹٖ��ܢ(6�
���Ζ��D�6;w�J��}壨�.s��(���L�aM�ѵ��M��a;��KU���;C���p�gZ��&������kRET�{�u'^]���=x�!y�4t	A|��4	{��ـ1S'���fR�pw�����8�*�M��͗ex���[J�LŎ��5J�x�Q����V~����P~�jʋ���w�v͒L2�E�0J�R8�\tB
;��2�8�� ���ơ�S���h?q���W����i�b�R&����-r�B��T ��+�?I�d�{��PM�M jd���DJ�8 �K���Ɇ���hި8��u���<�q7?궜�����Cp/����V�WvS��1�u�S�AS$ĸ��R%#T���lRuϥDS�Nⓟ��7��Wn���*,�����=�&��� g�⹩y2f"MՕ�C}���i��zы�$Q��@���8�OtjyF �n�)n�\��Ll�R9 ��vF3(W#�����U��cX�
�>	���Ǹ��t2�[��/V{w_:DЏ��q��~�+��$��h���|��۞^�$�����q�XF�1�W����*uǔ�b`� ����+pm>�ʁ>��18y�kvs{�9�6>D���1�Nw�ZV)Hÿϓ�[.b-�$�&�>	������
.�-�p�z�=�g�֧c^U	����i
��rM�˿��@r`s��}4�kͮ �k9<�H1vnÈz�E�7[c��P7�<*�Xw�(i�]�@��q茛����/�d~�� .�o2�����~��d� R�� +����ƚ?�ёL�kJ�������������Nu|o��B3�X�1ф�s �����6Z���}�L�|tV-G������ڠ��Ʀ/�܈�,<��v��D��00m�p�����W�p�8苠�HyO�i�,��J!��0�H�Z�!,�k��4��6w�_���@Tﯲ��A�]�T<h�d�X�uJ�ġl����ܻx�b�x�~@�E��gbC94�kX.��&�y+��da�p�uu��P0�������,H�����{}��o�/P'��7�m��I��?���PqV���I���a�ğew�C���Ĳ �����&�Q��9ZQ��\r��_//���;Z��0�:��E����?{jƗ�]����']s�}�X�
Z<��R
�لM�5����}"eE�S/�y2��C��d1�Rm��I�����D�9��GH#I�rU�FcR3T4g�����i�nx�YY���3�-|�{"��(�=���g�A̩H�OGn�X��!+Q��Ձ=Cf�fqiy۪
1$�	�H���t��t;2Rȣ�й0sG4
���Sii�Y���@\��;J��E��)��t�LO���҅ၶ������[N>ʳ����gG� l� �u��h�;��v����𾶳�ĺ*�,:+�W	�Y'���[��a+�LwJ6e�����wkq;&tD̗ j�H7Т�R@���dƞGA��X�������^}�J��\n�_,� ��z��A�aK,N�6�R��&�~��w�Z�xX�2�y�1~m�a(�&%��[d[ԏ�� ғ�� ���_K)�lp�s T�n[�s�7��I��Ag��UN���1(Z��i{�b6�4ň�x�/g|H�K��ð���[�D�?�#1�?��k�Y��?L�vKP�q��֡<�I����\]��Yhl�~��e�_\��_�ոz�p`mN��X.��	���xD,Th��2P��Y�B�����]_{J��U����&����JӶ5�.x'���A�GϬ���U2�0ǋ��)��6b�1O7�i�<�Ӆ"K�!Wh��L'��c��J���ϴ&�ǋ^���f��F�T����V�9`�sI?7���[��Vwdm��4'�d>p�m!m�5��K�=�8��QȺ��%�#|�ϑc�ѣkC0�}�E�~��9�kĀ�>g��S�+'a�|<	W .�&�6�uD���t�m���N���\
��ڼ�O��l�MᴫFڷ�T�Iz�����~D�vwg��	�e�Ѐ�.�/fQ��"_�	:|��IU(	�����$�'�˨���wU2�tM1(��M�57����	��ҲmPB����~a��6�C0����J�@���#%`����tƫF�Rn�mr�o��!a��A�F�ܪ7��I9 ��8O�-M.��E�e-%(H�&�<ًA��_r��w�/�X��'��#[��A���餍�pw��<��Rl�ŬJx	�y=/�=Qy�IΈ:��E8y���a�$��!���k���R�ȟ`bh;�-�D&�f$!^����%F f�
�D���y� �������)�hZs�W:�ȆM4���n��w��s&R�@��}t�9\�Om��h��v�p����4V��gM�6��O�lb&�g�+�XRx}2da;/y�ޘ GC�)� �x��|L[74f�
ࠕ���t�龳#O�����J�T��:��1m�Ƃ�#�_M�#m��jH�L�F� ]y=N9��A��,�x��qY��
�	6����Z��[�Wҹ��W�P}v�Ҝ�E���;�2�`��}r��Ď������s�O���2/��]���ͽU�����9��Lk&/�����[K��l&Yσ��)�=����ۀ���𦧡��1��ur��u���"�G�q���îV�;�?�1?~vXv�a�;M$������}�U֑�U�)p��v1
 ��+��hu�=�_�P�AFQ��-]����I���4Ǒ[�^�I�-[gU�����gV�z��N�v7N���Rtx���"&P���u�1-z%4Ü�H�Ott���p,s�W����}K̽�c��I���NW�<|�>Ե��&���%��\�	��x{ F	����-W�~)�sXP$�}�q��i�&B��o+ޏz�w���D�u/��<����ܯt�dQ��w�sOEU9�.�jD����z��h�"p'�k��d�V8	���"8x�R�x� �Y���,( �!�e9�k�O[lޖ���V/!������S^�8���W`�^	�u��o��J��|���o����v�	�JA�G��`��Q��O����R��A�r�>�`Z��U���#��CO"|���1{\T�M��)MO��1�8Qg��'ۑ8Z����GB�}j�I6)20��h����ge5��ܯ�?̭:n�5�T�b����v%�Pr�h����9I��
�>w�6у���q���c�������8�>Jj?ȑ��%[�]����4�f �G+�|0��m��7��T�7�V!�^Šp.ݜ�NC3K��1�*yU/��\ϧ�7'���#�����k��|�U���s���Œ�H��������<��7S�!��n�oϿ�-�Rk6W�f��#��dh��]�ˮ�u�f��M|;K3ي�Y���-,S�& s��귡�9[=Bc�R[��aPt�feFQ�8z�J^��8��~�r�	W�"�r2U F�gx^/UWb^��\N�X�$V�Ų	�zZa�Ψۤ,�͵Btjl�U4��	���(�+��q�{�� -�Ƹ�؅�N�e�����-���m�Ug�|����N��'M0��, B¾�f_��.t'��arj6���u`��:5|2P�����M.��J`W���Rh|�!?8%��G�C�Ō�=�O ��4e�����;gP��4����威�(�pC�y͡4���wwN'�UI]nJ�`W�	�e���?�@:� �E(�3�1§�4�]XS�T%j��Z��Ay6�vqFE���F���藹��O��FƗ~���O��������ݜ�\s�w�[��hY����$w�6���i�r�J>�3H�����@�tL���7�m�F c�A)��;t]vJߪAك&����/(ڴq����@B�ƣ���L���ܻqn�� ��)��	�2��oPa�䦣����<E>�����[��� 9�\����	�x!�{��^>�5�t�y0˗yNA*���_h�
�P�!��f�N2a[�d:O��U2�ʊ��E���l���BE��O��,d5q+�L������
P^ڸ���=\K
1�i�J+�����_uu��\�
�����C�l��e�6_�~�~+�0ĉ�2<9���4�����Eģ���͂���|]_���л�d�Ad�(% �������i6�75����ޤl2N��(������	*����̃N�M%��S2T5^6�q8�skVj�3�'�`�N�s�i3&�AN�lJ�v�����Psǽ�@A=>$ilG�m��2���Aup��Y �P��h������!�!u���&k-��O�=�+`6�]�Bݭq���ѕ@v�_*[�JȤ�-9B���i۞G��k{'u�o$�C������4�c�,Y0����Y)h����HB	���O˭�n�L�g��W�N:����c�^�b��X�j"����lHEf�V�ۻ�)��<��T�4�;*U93RF��wsXz�E�{𸕤�'����Hj�!���d��D���%dz�"�1#���Š45��on����5�1���R�shm\trz�-�Y�-Y��XA㒧k��GNs_��2�=��B^rv'_�!�X�Ӻ�<��_��6Aq�b���T��"ʣ����Q{{{��,�S1(1�yx��i�X�BZ�xȧ*S`��-��t� K%�C��z�4�0���&�w���p���(�1e��d@^��z[�{����0��MZV�.>�D�A��Z���wF�l�bPn��d@�/�H���3o��Ͱ���3��J��\eG�pޠ�қx�u�r[0��/v،�{$K!��@�^��WNO�d3�V���.��A�*��QH�(2�U���R�\P�ר1����Z�0B�U��(d}�=HێԷ���2�9����L�� '`�gsB0@�Ј	����O�����G)1�f:QD�0ks`�ك�����}����јð���g�QA�F{<�NP�60�k�����T*��{�|��_|���ׂ����Ή�r,U�^�*k�)1%v����>��V���`P��O�S�uM�B�?8��v�K&��D�sIԉ��Թ���!e��U�V���2APF	�?�Ol�VL�m!QNU�V�H�ȎR���Qpt�(\��|�%7|�z��� 1]*�˽�RA,T~r��>�T�.�:�Yd�_M��L�����6i�T�r}`�Ww�"j15�x���r���u뫉�<����ئ�'"iBm��ܟ��"}�>�>WF˙�l)B���Dm�Q�tmdo9l�7�v�6� ���A&��VL�P���}Jl]�Հ�,	��v������p�?�i����N�=.0۩A��oD�f�V��fQ_��.`Y��9R�7!q+}\����%���"~��Q�e4���ړQ�r�����| �s*@AJx�+������{t�Iw�� �V��Y��c���;���� �X*��hu����"�N�׀P�-8�~ݪ�*�>��c�ҍ ��L��X"���BAМ��rv&�. ��6Ā��[��؉��ɮ����!�����w�2������8_k��|Gi�g3NL��S���u�����8�W�ߴj�!Uɩ�)�Q���ָ?l������o@	�����^.�ITN1�S��p7(,]M<�����_�`ݸ]���Uo��rUa�1�9�fL��}>W����Tߝ�C1U��&�]�tZ����֎~+?S�4���nڅ��9ib�<�R�W���v�mR�B�|^�1_�j����{�z��0ҥ��1d딘~�p��j�6*]�R��$;�}�A^���ձ`���N�g�'�J;q�|,؍؋G�k��-[[+��]|�����8b��
��;�D;����Xz*Y�.3&#v*�F�d|�&TH����^�����,y� S��b�:L�ɠ(/�-
�>e���I.����`5������Pl��~B�ߊ��N���X��+|����"�2X�לDf4.�3V���.��6z�Q[�VU�1�+���C��nL����_�1�A�џ\i�v�Cd:�=����WÊ����ȏP�k���my�B�@B~���~V�E`��?��QE���q��c��9_�O)'�2k��8���wq)�9l=�i�Y3g����eI��Zi�db���CM�"��R�$0��E5ʘx��(|�L��=��p�r�l�R�p#���qfb�Ԓ��q0���G�R�R��-��׆}�ɚ� �Wg9�Ln��/���͍~M�qf�N��W ;:���U�x�;A��ǎ���d<��P���3��cL	0�7[��4�3���H�#��L+��Wp�%�]��ba��Ȣ���댭x�KJ'{��a�)f��'
�M	t�fQ5-2Ph�x�ˍ�����x��'����X�����h3���h��(�6C��)
���X&�Q��RM�i�?Vn�u���*[g��v�r���CC�Y��HT-�s)��� xh& ��.4�n�����a��nN��֣C�j���V��uI��M 3�~�{o|^!o�ôk^eP�b��O[��e�G�����&vt!�X�q{,�Q���L��x
ތDS�Ͽ󠥘��)������|���>i*�|���6pV
�V"��啄�ۖ6E��4C�8s�@O�8`�>/�OՎ/��~Y�����կәO��!0��Ps���3MVf�n�)� ��z_�����������A#_QҾ�/b�)�3'�
%�v�һ���]���%��J|Aֶ'..wd?A�jM�7I�U0QUMS���^�f�	,�J��Ͽ��3�uS��TV���KAy��12_���7���7S�,\4[&�3�����U�a���e����Aڬ��8� %x^e1+�+0���zf'�)Mԋ�Ʉ@��w\�����֔St1�'2A�޽Mu�߳y��<呟��]|p)�s��4E�Pۖ�g�$:�v�K'���~"��#wRE�B�Lf�"��������l���`�e���o���C$�$.|8�(�IN�.v-�!r��_o����<K�.�N����p�PЪT�uv���>�jii�d�
�?�[ڀaa2=pi��1޺���Ăch�,�p�\2a���R`^�	��Sy�̢��f��J�j�}��!�2��t����!$���������ٯgᬿ�998aB��ϵ�eލ����$g��D(9ξXDkdyn�]�e��5���n�V��X�))ό�.Ł|������~\f�nG�ۚ����Q:�TwƴH�G7dE��n<Qcrob�����%0����L�\	OY�t�T`��I�Q�b�ܭ���eh��ƓF�^8ū�y �=�GK�2/���Cqa��_�3�p����4���[����Y�fc�*ݜM��`/�d��~�ⷃbF�x�S#F�%����[�w��\����6տ���o�N!}פ�Q��)��$���SE[;�WDe}`�E�4�h�,V��ٔΗyg��=�r_�7wF��O����/˥��`N�-��rqq��6�1zkCh��36�H�yu��ٮ<��C+�%�K0{i�bo�+< ���~�e8>����`ȳi�WCS�;ʁA/�F�KT����2�/R�^g�e^{��S��s�����5a�=o��A��e���@�y�&�4d�`�G�ܮ�ْdAJ���1����[2�N>��.|���S�<�wI�:C�IUi�����"7�ER\�Z��첏��p�n��9K'���Y���Zs��"m����\���5oj��P8$�OJ��Wa*� "�ޖ�'r�=�v�R�Г#�}u�N�4�[���i���R����Q�	s��v(L�C
`'��Mz���h�j���k�.VN��`�R9��2�RE��>��M���di�&0᠛[w���FYS4޻���nY�Ț�Q��>�R1�>�s$>m�O���D�,�w�P����(B�&>0��a�ӯ
ɜA���k`{ڃ�}��L}�������:̂����c>�=h�z��ڃ�ڰN�͉�o����.f��O/*t�2"ag�n��r���\�&9*U�����˛_�Г>'o�1�:@~e���X������ ���8�:�+�S�C�5�D��m>vɹx���\�e�A��0�`�=�@���k��hi<La-ES�%x7 j��Q���2cAi]FIJz������ ��/Ǐ|�F>�X(�˕'��8Q¥�L�ۭD�=�%��9�%M��:T�;dT��eT���eh�+o�??^��I�z�6�}�֤�Ӧu��YC�Z��%�8B�b���f_3�X!"�;֭�ByE,˱"y0��[������(��RI[sG�F&=��Л��)V�ΏC��7F;�R�&v�/��g��u*
����[���$Fp���,b2Z�`vU�k!�D�������~Y�+mtnf�%a�lo�[�j6�:'�<H��y�r\ƟD��C�e���5���Y���;�f� 
�ű��M����>������͜��we�N��l�S��\[���:Z��jq�<��L��<��i�v6��p:n�<޾=����h�#i��9�v�Yh+8���G���ܲ=#��!4\��4�ί��^CZ� J1ޡxP�{�2�k�����J�'��~�@/ӂ?m_�gbu ҇=�����K+P�?s���i�<�(��%�R�zo	�Z/�֘�m���4��g�k.q�!��i���9��6������v��8ư5�Ql]fQ��g�_}�m���W����G����E<I	���c(�r(Q�^�f�W,e��
�Qjw^*j���U��O�	V2�D �;~F�,��/�����D��/v~�e��Y,c�Tw��F�$���/@�Ԓ��k�w���M�/1��OźR�WGҀ��K�s^ �՘����eiΦ�[`���J9+IN:W�)�hXOTW�Dϧ�'�5���L�
���>�����F���O(�{�lWݺ�W���	C	f_��+����gBɺK��\����:�b�0���G��D[��ú�1���޲}hf��օQV��O�Zd 2�ю�+��J�.�7�*�Z�"�Diz61h�!�>�ߟ�ZfC	���S��U���©��JDز��*|T�ߡSzyz�f�1�`4���GU+~y?T��$�>�8$��	�P�����J�>�/6ro�Bކ�������f.\�"d������G� 5�e1���Ș���5�#�}_��H��mP��{�GR��	�-ϥ�r���>���:i�F�8C�Ȳ�4�
����.L��|-1�N(�������b'�\�}��٥��?$�0���6)u���#�¥�t����J��stbH��p��TFt?� S�|�b�8�Rg);�}��`a�h�U��9��7X�� N�L�A���I�*m4��`m�4�N��[)8Y�d��^|Q�}����J����� �žE�"��E*Y�
i�;f(�i�w�����Oُ*�]��bi���Tt���$�ɍ*W�g:��"KD�-e�AR X���c�>rg�<!f7Î���П
���c�`+��B�1��[���s~�m�I�f�'�YV��xRQ��Ĵ�)]ޥMm �)Ԅ���]��;����Jb�cU�}��-	S2�$�&���W����@�������ó\�(w�I������gv�'`�)�V�(�g�3�F�c�n=����I��v���#"�q�*��3붗�h���`�}���v������j��|�@)�����\��Z���3�'-k����+�$�|�@�|���@'�����n��������娸�@pj�&(Z.)j��'�t����� �z����6F6>�K���
�1���s�Qm�x�Ń%�,[V��>� �p���jyhCO�vw��Ņ�__ܒ��F�����}v��mu��g�B;�� '���˪�K4U��2<�#g4TԹ��#,3Y�E��zXnvp��y�ߏgx�X7ߧ����M̈�i1�F�	�q?��U���i��?�w���=�.ԺJ>U�M�*�<U���G!��ܨ��S���J�������ގ9f�uGZ�L`lN�4m���;��ʗ�s��呚'2��1����Τb��)����<I�}�qk�hz�V�(�f6��X�u��.N�ݷ�&�3An"3[�n�̣��;������q�H���i��'j$�\�ԭ������MU�Ls
\��w_\�ƘK��Ҟ~!�`�{(�0w��^�#���g�A1��p����?7�<-��6�]��s��>�Q�v���h�MJ�y��f�Y?^���1f�\U�#�E���Xh�� �ɫ���<>(�_�d51����Hv�d�@
P>��������aE���◑h���c��R�B�����Ə���ފ�κ��4Q1����u@�YP�I��?��v�e�pC���9f��&�R=�Eނ�G��z	�&{ah��hzJ�(���f,�qn��vw���Ap[�T�I�N���j��>e��e�fa��a1�h	ra�����Ɵ�M�M\��{	�C��'��GRm��Z^�kK.7+���ޏM�{�t��>Zł�ڔ���zٲ�Uu��/ۤ%�%��*�~���c=�a����CA��-�#8�Ҥ�B���}v�'9����߿v D#,C�����E�VHT�f3�4 )Jyv�����:�Z��x�7em�m�cF� ��{.� ���=�9���j��T���CI�a�֩����<!����S�9J&�Ձ
_�\`�9�[E�D�u�9����_�"κ"����y��{��t������ǒNOU�P������E�����ڢ���Q��@6�,~#�C�Fb AՁlXw���*H�4���Bl�A�nj>χ<ס�֠����\���V��~	-=$p���%s[$z�� 5���G-��o%�E���\S�X�O�t`��\�2����Ou����r"����SI��^E5<M4�=�K⇺R�!��0DD�lo��~�ן�!쥎H�F�J������i���	t�`�� �
�O��b�AW�[=���R�-vMnD�������I/
�e|�Y�L����,�T� F�a��y����g��a�~"�����t�7�
���է��Hdo��_��ā;\�)��"�6� �Կ=Q��S� <�ɱe1��K;H�f������F�_����Y�~I]��w��;\�6����e^�'R�;f�
Qn�s��G��3���y�Z6��H�М)ZZKX�>��~�^Mt`t�ן�M��5'�<�U�\6���#��d�{{���&��Ad�^5
�hn�>qt��w*�?o��){���!_]$5Z����qj��8�C��H�Q�v�v��O���nۣ�D@�^�j�/�)��7#����}�X�_$a���Z'Tpڣ��o؛{b�l�W`�>��=����g��DD�v���ɗ���'Վ�	� B �N�����H������K�!�Oǁ�����&�<��Չ��U���}�A�	�����:�6OAݦ�';�u2��U��t�׸�ϧڼ �T��ϛ�G�wR�1�^BsvU�G������P�m�z��92z�h�%/����u�}r���3d���F?��&=�vz�*�^Q5�p���(��o�im
�h��s�#�~�$� :������a�+
�7�T�Q���v{� lƌC���$�:�e���"��Y��L��9�r�ps�_��p�?�L��FOk��F�8\}�s��Տ]&��y�4��V�E��ʛ)��X���I����U��)#¿�;ׇB`e٩Ч	�ȚD�]�W^>ȥpg��6�E+�\���hu~�u�l�p�J3����iAj�Y�x;��z�𿍿�^?������3������в���3}�5�++��� 3�`1'UY������t��^��3A
:���b
 �F�O��_�@5���a�
�1̂� ��ɤ߰1���-�� �,����ґ�� ��b�s�.�T��w�'2"�>�d%��_��XS�z��3�z��#�B��Sr��YbV�����g�����Xo3�?�zTC���`t��U5��ۉ{t�I���;�k2}|��.�A�@�a���%���	r��eѳ��!YU�\����8�.*�Gi���q�Q�]���.�Q)~Y.Q��v�[�B���4M��$b��1~AKf�څk�0#�4��&��{���S�:K9+�ڒT���G {���t����7
l�1��0bY&�ĝ
��*8��3^p�:7x�._�*�'Y�G.�9�Fl��evy�h����'uU'U ����꿖����2�`́�[%\;�Se��xF�r�>pq��>�m?�,�p���-���膚 ~�쌉��Т�x]P����: O�T� ?�}K��*�J�A)�\**�byqc�v�倧 �+4=�F�k*��P�#��k
�w@�f�g �3���<m���d݀��'��q�f~��3J���������Ii��wN�g�>�5�S�b֯���B��SxyJ��}��&��0�
�0�n��!�Y�8?yD�:_����lr�^X�NK��L�u��T6XJ�bg=�q�R�Qޭm��3����$A�����+�<ڈ����(s��h0|��tt�(�X	8�-��Wy�p��P����L�'���.��B�8Y��j�De���C7�}mw���l������!�Q��R�b�0�P�D�J�I���m\E�e�!�H^GrG��mהI�����Q�W�	��d�֭�5v\-���l Ў���w���:T�KR�h�@��·��,����"P�,eϸqrس�/��Gw�Z&YpT��/�(��G|�J@y�3��X�����6��)�c�2-�2ǻq4�������������1�Q�o^z�4�W����=����m*���c,˷�;W��2�dA ��JȺ�pi~�8V�[hlf��J����������B����#'zE�B����H2�o@c4�W۷��Mt�%^沈?���T�����b2��^ҫ�������/��e��55�$q��JR���3Rr[O����eWݧ�r����p���h*�Lh��ux�H��&Xs��2g��AAT<1K�^�3�����%(w���;N��쳻~�R�U���7I6���2��!�7`qC\���w��H��˅G�B���m=���"DՀ����feOZ���?eYع[�n_����9���3��#��<z8����	ZٍӦVb	3jap`�?�(!}�i7��$��b������W�ـ���t��P9���_���ч���n�;8o���OT�˂n4P�i�,x�v��Ͳ���;�~T���=�_D�V�?���o)}��sy���>�\�=P!uz�p�ﯔf��yG�!g0m�����������o{�V�g�7��	�y���`M�G ���f�vV���u�]�J�@���z���oy�b�p�᪩���s[��6�'q�j3_I�.�]��~���H�������٢ō|R��KZO�7/�P~�Q�� �e	��y��[���_IM�аy\���Pb)m�$�>��Q�Gs>5z��Ƃe�)AP��{���u�q����@}��j��0;�^���\d_�&� �y��ڔ�Oo�.Q�U�\&M �4n{hX~��eV�g*d�ű�m�$��v�M�2���G�=jJ�=��	%����3;� ���ٿL�=���(H��jр�H���
�n	��&���DAhvP�h�8o�4���r�O�{����Y��]ã��o��J�<~|��F���YD�x�� �<����0�δ�}�3�[��x}Q�ڧ:����w���=�&��}nʗz������:sH�"����%ly� �Z���k�F��Y1���9���f�]�q��� < |俱W��>?��P^Ex�X� [��)��g�uM$/�4V܂m�����i��)�/S?U�=���ēt"@�R5�7o68�
�f^�L���1���G�+�Qgq�T���0�=����s��v���\���l����N:
�#Qe�S4�������,C�7S��R҆�������N���òS'r����4����c>����%�k��7�W��t)�{�SV�z�2D_�4�Oz����a"~j��~����3��}�z{����<R�I�bx����e �=I���@��t�Wj�vܵ�'3�:��vt�#�Ҋ�������A��N��T��jg��rJ���3���c�� ���,H�r$��f�Dǰ3a@��3[���Ȑ����b06����7u �e�� ��c	��sT�6n��H�2<R�x�"�_`?V �t�v])���P���d���	 z8�Wn&��A�OG@�"j7��b)�d�Լ�.2	$���4��_���ۛ����.�8�Ʋ�$0�ݕN���.�F۱����\\���6�ދk����1���k � FF��q���ئ9�`�����Ѯ����ȳL�ф���to{�ֈ��K���+`�O��İ���΁U]B��ӟ?����m$P�rE��s������0~C���!��`c�'�/��[�E�h��Y醦��������ΎD+V9V]���uGItjf�.�����Cy�#�}�HUsP��v<R��u'_'뫿0H��m�E�be��:�����:���¥7OG9Z���Mo�hKָ�x�D�
z��"� %��Sո�Ke�����;ȭz8,������ـ�o�.j�1I�� �7���U^m%�ܱ��G�$):�3mG�H&��a������$�f�ufu��UX�$��@M-�3���j�A���c%r��tMХ|�>��L�X�)D��I��}-p�fX���DG�]�p�����Cƚ���X+
�Mj9B�ne`r]�-@k[V����QU<p
��פ��A��EǷP=儿9�'�29�݋���71����۰4�����c�ߕa�?��|8���}�~������Y5=wɐo���5cy2� �x�pbJ�[?+f�e��Bh'X������t�����Sy_m��pe�t	K�
p�H�gxm ����G�[��q�G�i�/;�mP�X���:X�[�F}�[Z�¯�	ʝ�0���%\�'�L7���nMC��B���k�D��L.�	�n��T���K��Ə����(�F�0��9��k8	�W���_`��ywsjRVa���	�h�W�5��Rז�[#���|��+��&�a� ~�v
�������H�ݠ�U'���e
�v��m�j��U2~��d�b��}ɔ�a�����C�|�$�:�V� ��B����:N��*�@��x�Ӆ쎚"��g刕�ȠP�d�v5������ʴ"��w�	�ڒ��l+(-I�|���������h��4m1������Q�K��jޝrS�3�J�2tt髶�0?�����(?qv~w'e^B�
Ҷщ�$���9[B/�ԡS��w��Ms����&�w�L�Q�tx�.�����<��;�Z17ݣ���=�h#�J0-g�L�8�|c�Mc2P�VѪ����3/��E�=���
��V�L"�ʣ[��&�w�����Ù���+���H~u/����ė��rO������e*ƻ��S)9��p�о��ʥ��}P��$���H)!�#����Pp�N3P��� 2�T��wQ$�5S���@�?�[H����tW�
�M�wL���z��B���њN40�ُ'e����q���M��z�~��3h����떬�f��DՇ��%�y� �M�>L�3;�b=f�c�"�<�!i�I0r�/0�εr[3�k�DG�W®�]1�o�%e�����0U�bf�xq �x㜊���&��A0��3�\e*aG�����<GZą��w��V�RU�|���k@rG�`�ΖR�I�X)��]ft�nV�cp��):���)"_4����U��菺�oډL� ��J=C�A��| V�*(�x�X��Զ�֔��.��z.��AK����p(��V�9)�N8�׿s
�o���(��D�2D	("B��ђ�Syi�*&m��h�����S���(Q����Z�̲�<}�%@���E_*��B����,�g}��͸!�A*6-Щ/�z� )��"/� $N�= ��O1��#-GUd.��;��c�aS�,��AD��-T�[
c�r�'
z9I(롴�̿�>���%ק����+�s�bO���+�1��*�q/�JN��nA�cb��"����������ty0=\�#��J&��rrcex�"�2₢Ĕ�/�C�_��2&K�c.����q5R`�evb�Y���KO)%�G���x� �S�_�Z-@/�S��z�9���H|��Oi��x�%��� ��z�M�cJ�hi��Nd��'S���E�I2s��vPu8g��S�\0�Н�+���I�E����=��j�ˁ�Z��p~������S�;>^�
���ni����(�R�&���`�A�mb�"�;�����g���@'L�~�&	�G�Y֮��W=�dyL��ϊSL�R}wG�b�;m���Q)� ����P$���O��{<rx�hK+����a!��[����,�lc� �����]�4�0�&1�"�alN��Mӡ�^�(󯃢�ߵ�ؗ6����2�A�)��:uE�t[ǝ[�O��L�<�)���F�������G�<��Կ�"��ӈ�Y�����'��U���G�q7���������@������Rt҅@|i��+��|&z�b�E��Zӂ2� ?R�Ds�8��=��"�Ê���U�ǂ��g��4�ͮܯ��@�����J�>vG�7X(w�F���rey� u^��*l�'�$<t�M�w���נ�#��QavbE�VBVw��
�'�I#���?���9�?�x���j��_��:$p�d��u��Uδ8U��ON���=N���M�&���яEzpLl��L��	@��!¶��H|�KF<�(3,�e�ɽ�l���Ɣ�x��ݣ�@��,w�N��<�:8��o�{/����YD�<6�Ib�}����ء�+l娨
�+�!�1kH^T��p�v�|u���������,�FL�����F�����Z%����1^Be�{Ͻ�a!:��,�XY%�3�Wr���~���B���*Q�ұN ��`��0'�]����$��v*�c����\L���,��r�v;�K���L|�L�j��v�H�U�ĩ�*��|.��m7v��4�Ĩ���q�
NFi9w�S���E*]���w� �ĝр+h���!�������g(�hu&dLߌ�T��;�]!jPM�8U��!)?�G�p�*�b�N
V]�����-HX�MOσ�!>�����*|�����ۼ��DnC=��cɂ�o�;���ewN������K�-d����4�sm�#�Q�EZ�W�ɢbr֕I83b�vLep#L+s�ת77�ȖP=��Vd�"���쾰/R)��(7��L_.�eۻ�1˱7k<��Q���G�#*ow�@\H�-�8+!D�.5���=� ��,?�R�JtGE�X�RUqbT��ly�~����7���w�ZT�y���"	�[/���3k�&���4-�a0�՗c�G���_���/�YN�wiϘ\ZS��/�BF��?O�5�w����?w'5:f|Llj�vp#�λ��On�� ,��cH-�LY��ը����2\���̙q�n��؛Ԛ0�sn��/u ��'2����Y��	��X���+��X�J���5��f7��� ��f��� �6�+�W�yr������PFѫ�'o��|��3\)���aH,Gx�+8�vՙ��BYG��0aa�e_���[��U.M��\�aڊOg��A;:�ʒ%:���0#�w�pˆ3$[��@H`	���*�c��<����2��mp�8=�av�Ӣ��p#7E�1�FEp]$�c�#�� ��lS`���F���(fx>1˹FH��&�t�Oq�I��7��yNa�;�%�u����eÚ���VP�5�
t��|�Kk��J?'�ԇ���ã;���>R�Cj��V���i���V�V��"��}{�l�E��̩�޿�])!Y#�{��K�N��K�u�w�<�w���t�Q��*ƚ?S/R�#� �I!9w����#�,v;���yE�U�����*e�n�y2���غr/�&G4�Oo���D��B�"&T��N�A)�&p}�Y
��b�`C=T��zq��<~3)���~�����ֵ\�S����$f��>����%���;\^.t����$$�U���~�ϴm3�7W��D����������U����z�����?ڕ� �m��g�F��8$�^������
B�0Z�<nad�0���Ս�R�����o����/G���(�o�x0����D?i���B�26�i�`��.���k�d���2�A
<�[�*��D��_CQ��31�u�.�ԵYɢx�8�e1���wM�	�1�`����G�qFc���7c?����|��$'�����Y��m$GS�-�a���/��i+��W0�F4h�������#���rpQ�V�V�=Sh; ��pT2J	;P�r]M��T	^7�.s����G�C�<�qz�$���#Y�ݭ�@���.�]�K��u�h�B@r�����y2m�n��pi[�.���7�L��E����|��K$;R��]
�Gg��ғ�]���}$�д����G�ǅ{���<�n�r�um��?�-@`HP���aU�����m�]�Y��&�֝�@I�#���e�m�g��)�� ~��qɅ�H����,[{%(`��D-x�+b�;�!�.�Xs�+�ȗv�yH|5�Z�h�u�^o�ۣ������)+m��gF}�Ϳ�YGG�����{��Y �>��Zr��k��f����b�>�c a�tF��,�Ec����Or`k1}}�ڦ1��Ѝ��� }I�`<���}��f=�1�z�UA)�:qW��|���G6VH8�AĈC2@� ���:�5��N�-�t���/i;ca8Kv,Ya�H7�e��� � �D�1|�Y
I������-v�jMCD�iXF�X�J�D���N�4�5��.���"�G[��o���Ko�\b
�zGv�;$K-�w%�= �R��n���1�3�K���	�'U�3y2���M���V�xȱPOz�P�p$��(�pX���.y�Yk`��9Z��ֽ�j�>.����bn�sN���ܑ(�2BS��t[�Ze�u,00�G"0��qdeo�Q�A�S���J}�����'��|#f5qN|	}:�ԕ
�) ������g�VϘJ��ϫ��Y�B��t�e�.����*�J����yU�dv*/,x]K�	����b�� �B�t+�$2�ܾ����iK������D?�1���(��Q(D����h9�a�m	{��;v�:����U�7��D])�4Ư%�%�Wq�ZT���"ZeFW�\sF�	>�t��%�z��.����vj�m�W�E�N�������B1u}d�:�~<�����uI#2+{��F���0�O�ݼ==ɼ`�t�ɕ��@�|�%Ao��Gf�%$�MQiAvc�n�Y��.?���?�\��zy����O���)d��9�Sp⹭hw����b�%wC���^����΋�0�Bz�\aڨ %T�:����]���@yA�F� 	nOC>���h��ߤ%G`��b�0Á�~�ְ�N�Ha��c�$غ����@���:�������������ۻ���J/�T~�'�/�|A� x�a���3%^Ḽ�!^BN��R����"@?�FK?�����J@w��SP��	�Y5��\IH�I������V�.��3��a�À�\�����wU͍�5��l�{�]���^�O����=�C ����>&>��mgMD"J8M;�]�[�1�N�����&�93o�sk��|���6��ќ��gg��*��jg0���Z!t���O�h�(J��R��'L�|V��qYn��r�U|Կ�n��p�
9%
�:������{N�8�e��̭����,����3�v���0S(��ѽ��h_��.�-�0���"��]"C�,
l�R��+��y��\�,r�#�UBĮ�W}2���nۖ8ArKٺ��C��{�rA��+�&��$�����c�J�m�4rN?�쉆J�k��
Q��%��>L����u���'�8�N�\�=_�d�mpl| �L͉�.h�/n�2��+B,n�P|�;�w�͊��9��mE��:Sn8�s :��B�(�i���,(�<��i��U;/��ߑ�>��,�^7�	�ge�½6<���|,�Hs���6�/���}R�p�=�]��Wf�s�T�1#����*V�#��0�ʬB��L`�,6�f�+�%�|��X�iԌ����P]m����7�x~9�ج�^��� ��ֵo�.�/�l�ˤN����c. �̾�ߠ/o �#~����'�>區հRc�M_��%K�%�przk�*.�����-�e`�I�����=����")?��`Y ��M���&9��Π|B� D�?a�t/���I�~	B9Dop`'6�4�:��|n{v��P�'����rߏ��s���{智O�k���������L�K[�����jf�#kN՚����\��� >`F\e��V��";{ɶ����j̴��x(Y󞎎%�LY5#��N�0y[9v[Z6�d��(��Q���ek/!,�v�zh�fuX<3a��t-��!�y���@9#�N ��Π�����n�j*(nI��q�uQ$ԃ  ���S)m']K	 P`i��l�>����Tf�3Գ~��x��[��>��M��(���G�97�s+L-����~s������5�n�3��0���!��[#|�k ��.�;�V�T�C �|��/���2c�8cQ�ʹÐ�`�r}��HNFs���Ygϫ�_̈́	�Ddk����w�h���4�aQ�4[=Ϟ����Z��������5��g�J���Ɍ�k���ԃ����� ��1�F�}��ڼ~X�֝Y��*hK���mn����bsJ �P&;�G����SXjx1r�jl��W�����BH@�c�kx!������k�2������t�VXj�叱���ne��	�L��UG����Kaj���o�M.��r[�H�dVF���\���~
�m�����=;���3� ��z���%_L���)J��+�Q��)_��L�M�HK&��ٙ�� K6����=b�L�	��$� l�$����Gmr]��;W��+�
�i����kA[�<��A������5����G�b"�B�\��B���ޫ�� `QGŽu�+��$�<���91�K�ϻ�=
���zR91�0��ؔ�t�G�"�h?�(��6ر�մ$�[�D5��`�A!�ӻ��Z�1߇��#��m}=�����H��~z����K��Zb�@�g!�~�@�e��zm�e�E�gk�g�^Ap��}�»|�D���%��bP?�t�#�.����GP��&��IFZHa���#��������˾?�NejR����|(��� �Ba�"�3��C��b���ս���vYFg�� d���am& �.�ŔC�`/�U�2߆�kG����e5@~)�K/�G���d�z��C���e��� ��6�w�Y����,2�o`���+��@lʔ1}���hqc�P�/ν�s���S�jc>�g����1C�F�鍘���T�� :�b1zpQ	P�qw^��w>��U�?����ْ��*ٳ�ӈ��q�����/�m�81�WI�MM�����;ȗ�܋�`H�~
�v���­� �+���^wm���/8���ʄj���O/�M�w%��+��z��dM)��-�Ew��Fo�q�g(#���2�/;�A�x� �#���j���.l?�ݱjXʝg��!Y�����r��\$�[t�s7F��-����&;�#A�I
x�ׄ�	�h��@��[�>^�Ҟ~�'K�3T����&,��*�0���ڏE6�k�~������H{�!�tۖ���.���������g�)�L��Ʒ�F�0��߸�`���]�G�t��F���R�q"w�P��I`hT�� �l�vrrt��������w0Ї��g��H8t��ѬFW��ӯh��1�X��5����$IB��nu���6j©bIxA�b6CDB�x���/[������� �M�>�1cI;���(�ӳS��w_��m�2�4J0V6v�On��FS��~e������Bb�P�1s�"��Dd�n��p7�J�y���x��s'��(t�67'�Y��!QM�����R�n��Z�ES�R�E���&qpJ#�3;rY�����^�Kf������C�M��al	�s�#�hpn$P�,R3�g�v�U��;�ͻ��l<�t�m�o�Z����h� %����2���R�>h¨�!,$a3��;r���Ëi0P� �P�2
ְ�T�}��HTV
����k&��t�-���3M�9�"w�>�@���ݺ��,�/~q�Z��u�*�o%5Jǳj�H�.�Z�j�~oA:<�v����;c-ckу&���B� 7�4m� Z�P�����C�ë�tWY�j�2���+�`JOI�H��L�q�i<��6<����b`�&7B0X1���q�%��A�4��3�$m��>3
�rRA����O%���~���b)�S�@��Ŗ�j�^����+�l41�09]%+��"��rx3�:$�^)-~o����w��ay�w�8-A����}E�z�U�jrTq��%Z����; I%�����E���y �f\�6���9o�S������X ����Q�v����B��K0����.��IaEʓDhVCln?�|��u���*�1+^�躲�@��2r�F�[�����7}~��-:̟�Hm�;��c(�_���ƾH�M^�O��|Z�=��$č$pd��;/�Z�9>*ݔ��+�Fr�@`��u$���h�j��X�4��C�˙��۹3��z�`x������3N�h�JO��}>
�ε�(����	���dA���
�(�D���nկ,on�vG�n��ְ0ܙ�����Vb	�z����7v��Y`���=�]_dd^�Ku�ر�<���h�'9�Z��ZOۻ&�߲�d~��{)DO�����`$�����^�MJj&g��3z+U�%����V�CQ��Pju��r���c=�p�ޚ�+ׯ�xjs(�B�93 .%�Gn��#D&;C��ty@;�@�%#�Z�*�p1�[���&�a�nl���%��mx
'�j}F���5��u�C���g�x��=%N;Hd�r�^tI{�L��~�Z���,�V����PUL-B�<���5�޺�&���G�'',��[��ɕ�8J$���DB�/�V:�xoe��iI�4��_^kOeR�tyS�ZG��� �f(QB�52�q����{���I�j��e���\O���B�E�F�R��|lewד�<pQ}��K� �cP[����$r���U��D�m�zq_�߯*�i_���3{�ƹ� ��������iז�RH5;ZՄt[���T��'����Yg���؝���+0�v�Z�[	�0�-�F�~LZ��V�|ac�&��P,��c��v���2� �+�z���Z���	�׃����c�$����0��;[�	^#02������f�Y��'6K���U@��A=yA���R�4�2S�K·�ʢ�����Y/�~��Z�|ۅ1@��rg�eĘr?���4��ƾBXҿ7��袭ZSuц�з&���7A-�X눮5l�faA�KQ� m n�n�����(�&/W,-^y��\��l�r���5uܼ�|t4��`f�1W���p���Ye?�0hD-O�d��z�L��<�v^?��~�\��i4��N�������Z12Ǹ�Z�f4����g��P7�P�t��`�x0�"��v�TA�HPH]��c�l$��?�^�
�ёi�f��3b�i�@�/%h��iF�p�F�[$�g=Sb;)�S1I���j��58�e�6�߿Ŋ���<��^��
r ��Uz!�+�8�V��A�+�*4�Ӕ���*�]�=�?%��<�K�w��v�� ����8��^1p����V4g-��Ϡ��TV��ef�2���� PJ�;F�˽�B� �f�ֶ��:O}&T��~jn�_��HL֏b��>7��S��L�PS�NX��ѕ�5�$
0Xq)��֙�a���2���I��`c���ւ� {JZXp�o�V;u��@���r���{���;6�U�"'c�i������B�K���Z�(��*�޼
���I��1
��g+����A�@Ǖ��}�_��|`]�$έ�nͺp��d��y�0&s����������I"��;��%�s�Lf�Uh�n�9��`uWR���)�z��p�,�Y��EV�n0
Y"H�:�MR7R���@�KU�1q�@9���ʜ�Xa��vS�ڠ��~8���e2}d��U,�"��Ȧb��Ms�~ ��|�#|�hD]����L�|�4�C��^2�����8���@Buk�S��)r���*�	9lrj��K`[�úm~'Ș��镼+(H��	���x;P�-�"[C��:a
�h�
���(���g3J\� /�un�n�~�Nnp�\'��לl��<�@�B�w�I&'���CP� �5��[�k}��6����Q�t�c9���:Z�Z�;�5�>�b#4�;o�Jgף�)��4j� �����5E��m'������m蒝�����D�2��5^�s� �4�Q2��=pL�zp����["@�����>����G��=`OpH���:�;�Զ_�%;j]	���G���`Z�&ar����Z��q�Z�mD��}G\e�*�:{�h���|�-,J�1}�6*we����j�GA&ln¨z8�(困:�u��3��*����9� �`�O7y�7W�T`2ȼ*4�?ύ+����_�|�>`����ݯ����^r�#y/�}��6�k�)%�K5w���iq��o��'M�κ�I$����V�րvŔ���vB8�R�QǮ16V/?�6�3�� �w�Fɔ�2�M8��Qe��Q`K�s���ͧF�Ŵ��S����#lk�}5�m��1��Rxg 	X�c�Dc���+�]wvБdB��Uk.FB����Y�2���:��P�UOC�.S��2O+q��!�54���#`�#>����f,x����{�|z���Ҕw�! ��G����|g�����Wx����a�{�ޚv~�c�i�MZ7q�#@� r5���m�9�7cs׾��s-i����"�e�օzj�H❘��++��o��ZO��{�f����S�i(�(N���L@��?׿��2A��0Yd(4�w���|6�,eM" nxi8��y�ͅ��Hs�ʫ�}K�f�g~�~�6��riyq���q��mo�@X����$b�_-`^A��D7�Q�ا��4 ��A�	) �,�mG������v^ԋm��1̕��
�f��ѷ��Hc�ڐ�>�c���'E��%�g==a<�x$����q�kOD���b�9U}%ĳ�s��v׽��X��A�E�c�^��N�/eL��)3�w��}�p�#��2)a�$$(2�§������AL�����z���a7w���EP�K��NP�v�P<@�5����\�l8�?+�p�c��1��3�w�1Ƚ3��4����Y)Ůn�ݪL���ؽ��vLw�����dc�a������x2$��Y[�1
�,8x;^1s�|��h!_��6Z��R�R�J�vrt��2q�&h��4�	J>Rg�f9�~�rr�x6poܭ��(��o�I.E�/��H�)����D�ӗ[`\��s��Q�Q���4=vJ�E��r�&@>��nBfJ:�Cֶ^�U��WO1k�V��+��.
]r�Mx�H�f��~M��Y=��@�F�'�n��7_�<CDg�i�$qز����Nf�d�|.���}��O.���4Z0�
�֗�n�Y�=Լ�Z�#�6��:3��&�|�j�wmZY�WW<��u�%i���ϟ�?]N� ��;�[K�6��"R�>�m��z�j�
d1s�2_>!p)}k'��_iSy0��/��)���9�P})��$!2 ��E0�e��[2��F#��E	��N�ϩ��񎱵����J����	]�,&����W��'Gge2,e�H2��O����v�9�1h�Q$_�-�99�s����%V�!C��Lz��O�l����s� �q�,>,pm0~.֕�?��j��%}���;YV;%|;�-Q��X!2ح�D��3�:�}�;zS[�oQ�b������b���O(�tw��!��6�#F�2\��T���툃Zy!��C_�{�^��d�OV%/�*x$\#�m�y��5������;G����&h!��̳�TN�j��t��Y3��I�~A�W� ��+-=ިbX���*"�Ja����b2�s���Ij�5���U��If1.�<�7%vGb�����e#�zP��(/ٗ>(���o�[K�ķ�]�z�drQ�^!��#��r�dD%&�C������Ui�(I8�F׈r��>�6_tʡ�lI~�l@oqG���~�6!bVͪ�W!S��.��������AJ���~��U�*X���H:�``4�^/��Qg&���6 t�h!�@�V����2�Oz���}O��������ѵ K�opH��qU��JRZO��Q��r�u�;�8� ��q�b���3��^����-�L�J�~ ֈ{�3R -U2o@�^M��$Wq�^�Xf�Ui�>�i���׉��NA��w�U+���̗��e��\5K�ipuDK���3�K����<���j�����;�**T!�
�s7�p���Kf&-� �`�c+� D����|�6���0�Ph>�����T�2�+��������'m�W�F}��St�uWѢQ����~��_����X�7+��T�1(0 Gq)Э���%%�%BK�h�?��,{ ���d��`��2靊A�vvW��.�mO�r��}<�<��1�ѥ$O32����t��]�&u�[�A���8e���� k��;سXa9`������Y|��WA��AR;��:[���"�	c�7�j��� v���w�s{_�^޴�m���=�| SÄU��%���c� ���v\Ha��P�91�*d�S��	��}��?�0�SĮ���f�g�\�=��?2 GwsrNL����} ��4�����8ZFK3�.���dr��ę�����{w��Ed{�Iy�s��h��u?p�*������S���:k��r�n�<ȸ[���D�u�a��Tq -�r,���,����N�Ta��>� �z3��')������~0�{���'�8]1'�ՙ�ӥm��^%ۀP����7.�ᚨo�����ƻ��&���6�㕳v��Ll�J@��.D�aZ�dU"n@A|�y������f)���*BtZ+JK>�m�c�?����o�|�0��Kr���FN�v3.���g�C2/c�1-�]��y���������������e�Ч�@5
�@mkp[e��.=g���sd��b!-�� ��8oK��sm
/
���68�%�PQ����w��k�Qpە���Ika���e:�{������N���.�mN�-����Y�]4�J�0qW��5� g�Zk�l�ŀV	�Xr�Uw!�ҭ��zR��Z���vk����*I{d����)g΄��t�H�/Lz�H���dj�ZC3bY�#����I═�8![(r�%��ݿ�$O��{�~uB��n;��[&+�5ڒ��W�����KnV
��Kf�-EBv�x�V0��a��(6���d���t����GU��A����)zu���̬ɜJ��a�/��F��1�|X��9[�iYY[��� ��o�׷T�oh��� ���Q"�ȹ�<L	��np�5�P/��n�n�r"�q1��5jܗ�����sZ�C��W<�!13�i+���W�Uҽ7��-�*�AH<+X,`�i�H�o������k���N��n��	,����T������S��3W�y ���h%�-s�S��j��4ڟ_�-��T������%�d�ۄ��\Ѵ�a)V;�f���7X;��"�:��z���O,Әv,���G���|d�����`#z ��*���^��V/��ҭ�\�٠z�q1�1H�-�������X>@�ʎ�v�A����L�KQ��h"n V�j��wH8�x��5��T����ɖo"���&���q�~�t��	TP?�9 ��<Z�������-F�\A�>-����A��m =��+C	�A]�huPVT�0�v��VIB��>�-x6-T��X�z���X'�z2a���5��D�9.ɽ����K��Q�����/�)BLO� �͝5n��L��ߟ`�<V8�77V�栬)�M��c��+��K)���0��Va�x���!{i�%�5,o��ѹ���$P+dϽ���d�I�dLLNP�DM��,?�NҚn�K	�?������(4�Hn-E�1�ո���B���=��0P��_���y�A�^-�wìWzk@Cf�O\��O ��?��|�<&��&�?\���t��K6�G|����5S��	�	5�U;^���5mC'M�B��z*�`z�r��H}n��`��y�~��>��;nt*�����9>$8^���"j@fHK��"�=�����Vk$���3�
,����[~���;������37r�Q;cg�\	o_Nc+�5o�[�j�����n�^�����$]aa�[(�EѲ����d}n&�D�N&�q���!D;��ob���s �����?�ߋ��-�1�i)c5��P���Z�I,f��mo�6K�G�Ď�b��ت��y�f������W�!����p�05O����^�J����N��v�0�P�gj��.|����F��9s{s�1bi+�+���n���Z�@)���9?wv��^m_�d���S��Q�R�9�҉����z��<���	\���t e�R�hY�I�`�7�)��xȲ�����Lw4E�^�nX����t��u�`��Fϊ���1����\����>14��f��i��T�j��0*!Q4�����>��3<�fp�dE���ܔȿ�6���$�I�W@���f�#5"Tn��?�������!՛�KE���r6U Z�i4���:s�h*v�H�R�7� �)md��p��L�X�s,�;t[Q�c�������m6>��rs���t��b�@�Е7AL;^	5��IPᬁ5��?�
֕��Y�^���F��3&,X�7�����$�M|����aJ��X0�rl�^pZ���eT�ti��������lR���8Pr3dd�t�߇s9g߸#VQe�ZtD�͹<�p�S�����J|J�����J i��� JH�Y<���^o���PC��E˧���A�}MU��ku���L-�G�����e`$�bӦ�(jo3��=3�j�JzpQ�ſ��H-�@zR��\)�����iޚ'=��Jն�Σ�>����L	�RG9'�B3>��sn���Rv_ɛM�%K|c���|�c�B���D�tOo��Qc��hi���0�T��ߕ�m$ts��I�\�:�xpE�{jT�St�0�U-|C�,�DN�S�2x;�oɺ�������R!"��)�Ε�-[_Y�k�tE#4�̎T1 "�m�"�A!d�o����s�ظ�y�؟�7����BG�P���!�wGǽ�*�u�|g�|��=@e��hkVi���A���!Pך;�_[�о�7S�-)���xǟ$�c������7ϼV�`ML��xI`?�76#����C-K��:E"��Xr-����w9��K�@O�I��8�����_z���7�SQ۴��?�j��4t�u��/�&�E��>s+1�]۝:����C�Hqw��=��d@�H4�	�q���m��L�!�.���vs:~c4@���4�u����,jf>9"�UNHc4���غ���e3�sVy�R
�e�X�:-�Q�O�����W&F��8�7j�.Sr6/.0�K�� �����PYr��|��i$s8�e���S:�ڟ��������֑s�L_���02��fe]���P^�̶׎���%�� �<hD�V�[?��s���M_�ew�nzs4�=?���1Fg�`b��1׏y�$�n(�Ś��� �*�;/��#��K�5����8'6�1��aJ�s-�zm,`�Z�'?;�J����`��_D����Fu���H���g횛���z�� �p��e��>|�B����->f�4=i�Z]�>������6����e����K�~x�ӦtY�ܴ�qT���bń�_�����;�	<eH���[�ɝ�1~"�X������Q��q��)7�Gv��$uC���-�1�
�m�kQ��mG�)��{b��Bpo]����>*���_�	� iŢ�H��:v�^�^C�[����@��TǦ՘��Xz}�c�ĩ`<@�e-:�T5��R�E.���з$�D�R�Z���@B)oh)��X 7`3�ʘ�_S��M(�ysk�A�=ʼ���2k�F9��@RՄQ�9٬3z�%�O<Q��k�X�H����v����� ��;mB��%�;� ��`� R0�U�"^�-~���9�,���SX��ΆE#%m<-�J��V�L�@�Yyn9n��r!��m��td=!�M�?��1L�+�t;��q&HjV��â�5>d,~���v�^5�Zya�=dC��@�dF%{9r�WĎ/��,���{@��S�G��Ma�������.J��_�d�N4�G������oGR�D�I������V�R�H�i�<�Z4�����5m�6��k*gp�5��]���(>H�y)jH������RH���0�	Gv)s�9g팍~���$�
Z)�*�=�����w����ز��T�n�?,ǧ�ͳeJ���yU#�Q܉��X6�b�'�@$�E�h`ت�Z��ʈ�J��r �mn?������Щ6�[��A<�q��%)M�;���-��4*���nOq�DQn~d����m�@�v���J�G�����<�MKH#Eln3@��W��-'��7�����X$΁� ���v���0lۉ&h�o����-n�����վ�AO�G|�0I�u�%���w�QY��B�5a}����\1��<���y�&���)�d'�2�0yE�ۼf����f>�QX+�%P�r�}� i8`+��i*A���-W�P�u��&NpBur���W�
��Kι����+�)�u����SJb[Z5��p���{.N$���"W����e�U�R_���o��lp*fx�i�T9��ε������B���c�Z86���
9�(��;���
�Ok�C��M2��_W�,j��i-������v,��]*p:1;b!-b�q�BD������9s�:�%͢����y�1�9~���y�N1����e�E��{-�
�@�Դ��*d����=�Da�N�a-�
�9��(`U��GU�F�1i�bM�A�}��!D-:Ⱥm����P�)G=�C�sYUbӽ�_e��ǽT��M�%��%�M�ګ6�	���0%�����&C�Gfu��8p-ES��O��c�d�]H��Q0�d�5�����m�+>��û����y}�ƃ��JU��b�����-�[�	��_?�J��=H~,��^#i�2lڣ��!��yH�eg��Yg`m����ˮ+�Z06HFB�����U{ӑ<F���W�͚~��*eW5��R �1fD���W��`8%HŒ�����E���E�A��nB��r`6i�A���|�~%f�%�c�Yf�R�i�D���KPF\k���ϗ�bl_��ǥ�րGo^y%h�����^>�D�Y0�z�{�5'zk�Q�8�f��j�@r�P��B���d������;��e�[��Y�Z��"j�����}���s�ZLqncF�x��QR@�V���ꩳ��M��p�2���l���[���,V�%���#��=�1#A9<P��<JV�J0�Tr�^5}"a��L�h6/\2����f�m#$ܐ�5���k��ho*�|?M��v�R$Mj���\��ɑ�=�n�}3����W����h�����а��'�A�r���Tq�D=y
;��55P;ήb]{Ob8�_?w!� �xⒼl�ˀ���e�P4&}b�t���GBq�s��D���!4`��x+bT>�т?%�V���/�^+�-��w>z������ dFJ��D?�*|�-�^9:o�<�ZG����<̼�1�]�鼝��2{k�xY�	��I���EF�*xu��}(uό�`e=p�m�rj�k�k)>����Go�'Hd��%�=ן�l��s'W34��B0�vB�i9�1�$Y�[U���z,���4�9>�-�D� {+9��Q9/�-$o�+����E�#�x)��`��|�!u�v��b�����ѠGiEL�}~_-K�7�p�$�w�����N��ֲ#��%^�k�����9���a�ʑpj�t���Y����2"�p����w�����,�3 J�WO-�_��6^M|�˶AS����Qe��^K9�Ar��K����v���(�F�h��;|������Z���,9Yړͻ*���?t�/NEL�T4��G9�Cj�J���Œ ~�݆�|�+м@(��n�߈� �y]2��в�J�G�8����>�d�Co�SCN��
�G�{��~�#�&���`�pu0��R�7<�(�]��e��r�?Q���øa�5��Ce���g����"�J�IV���If|a��5�-�+��J�����,�!�%���w=:�0j��ԛ2�B��|X�mf�&c��� �����ݶW!�F���(�w+ư��ZL��yM�gߦ��k�Wz�RZ4��+eg�\�2�����qE9��J�A�Ͻڻ4[i��z���X�x�CZD��i��Ďb�)����	�&��@ͣ���7��P?q��A�_����t�d��_���E�}�<C�j��h=z�4���?��~���`��E�� 1z�Y[���d�EL���3���T���I+�:�O����e8��<���7"�m�W�����U�ji8`�}�Yf�;'��<�D��^�s�:�{����f�����<@ w������]&Y^$�;�V��;��|4��&��)�f�h�k�ܡRU��u�B�X��g)�I=��nèA��h��g)���(:vKХ%+�%��^vi�_1�[���	I;��7;d��\ {�0�P��p�"t����Q�A =4ڃQ6���xI���8���$n�Hl�c{h!X��0��kl�1�5U9W-C��ł4�\:��'���e��/�s�8^����t�D�C�@���G��֜���r�.��y ���D��P,���N��n^W�� ��p��L���=�P��,��^b�1�&	�넗�����I����k���'�2c�-$ 1t:mf�:�6q	��$�2�E�x���fN���IZ��H�-�@?`����2�G�L@|�(�CJ|#֮݌T�;:X��8B�� �n��}�r
S��9Rm�*1�v�j�� qoy>w���O!�Qo%6����tb��_�@�ma����o��������-H��te�X���Au[�=��ׂ�z (w���ꎤA���"�=x�<cv'����=��`@Z£0r{���
�UX���i�x @�MF��K��D~��]U9чv䲣�\��?K�	B
�@j3p&ʈM����!�=vm$ Ska5{6BY��⎳D'8�E����0Ă�M�&������`�n�뜃�%g�WBAU�7U�"�T���;B���h�����6T ������@H
���o�!�_�,�kˇs��3�ef��;��=^�����t}�<n��r\գEU]v�5��6�ad�I��}��r�F�g*���BD#	X�U]iG�<5dX)��.l�f�d������@ƹ��N}hf�#�8k��Kn�Էؠ1vOpnv�����W)�s�0�+9�*��Z�n�Ov�A�q�e6��Z1�fY�}�}�zn�yZ��g�E4|��HH[����a�g�Ѧ�l2a�e��,�׀G�����n)X^�\o����k��pN�������l��9Ա��L���
�/1RW����Ɵ?O!-@�_p���r�$='	4�j�_'�x4�xM�ϧ�w��Y�'D�~v|qL�qcV�=����M���A�9��$�WC~&vn�G10*[�s<Ajc@Uنٝ՟m?�#���G^�$bia��쨙k��`�O�^��S(���H�
�F���W:>�.[��5Np{޵���}���C��Q=�q�g�l4V���]�ʅ��`N�{�;�<�e��+��<-���c�#�44/?	��� w����������M0� �5k}��x�n�G����_2����j��t1���'J���D�oCݐ������<n����̚6����+�d�?��Ȅ4345~:��c���I��������?i�cL;Ւ�N,���";E�� -O��h�1}����/h�����^�^]�"�1@%�5$� ı؛��^ '
����T��_���"k�0VMƌߦeLI0�9i~�V��|��Vb)X(Z7��n��f����{��p��,�"Ae� 	���d=�Mӧ�y4YT|/�u��d`^�w�C��'�.���M����l�-��$ÿ�v�S����3���A`��͗}BS�g�v�K�^��v8�U��<��T����;M�A�=�#K:1"�0*����$�H�F��3��Q��"�7��Lt;8�=�n:B���^ڽ��b��˭��M��^|Z7��]��v�'0u�%tc�q7 NRSqI�գ�)����z_�q���2Fҗ�J����ښ}�g��C����o�����5��"��uҦ���ѓ"�fP)�b�'� �[�ZoJ�7���72��,���[����2]`���dV)�!?�(���h{`L�l�ғ���?��M;�B�V5�`R���*Z����	
�*d�,5�sЇ��]�;�1z�:�gq��8�8�X)$�������hػ� �
�~�G�%��CS6D��q�i�m�p[��k~t�����vX@��7����;K��9���6���=� ����oB�<���592@�^���n���e�v�����vn{���}F��+���O> ��Ӛ�L	�e`�G�E�p�2[�+�g��578�C�\��{_�,V�¿�>��ݑZ�S@�#�Ai��Q|4��7]���_hQ�͠����v��-v9 .֩lq:�B�1�LU,�gI���
0|ы����@���0����0�n���W��)۹ۂe�/��,en���2B�׆F����ʱ`�v��ܼwQX�u��O}e��@e�]�������>%�h��v��EU��4򱒳��W賨�-��5��p!w6��^N�OU�1@����r6���V����G��� }��k�4	8V�Brm�b����tA92_��JWJ�і��U�����={�=M6@���=_f*�|>��=�U�:��F���[�(��~spw,�� Z^�l@�Ć���w|���a4we���
���1[x�<��pL�Ya�m�u�	�V�)�� {PZ�P޻n����W��2��{Qj��eHgJ�k1��@�c�*���rHf�|�E��	���zbZ�8#�S�Z�fD%���Bt�`��8�7��� q���8�v�4��!P��!�f��)��� ���595��̫2���B��2FC(F��%�.F�Dk���@���gT�L+k6���fL�Wܒ�Nt���T����y�@�/�����jJ��P�i/�^�L���R��VRc��%�m3����uRfs��m2�o������s�@(����Xb�N �\����(�:k���5[vfv1|��ה��Z��djn�٫C��X+e�$�����>����b��lY5o!YӃi�\ډ��D혺JRg����[�Sl@^Yưʿ,��_ ɯ����zk'�|�0��n/����T�ݼ��#1Y˘�j�L����)�a2���|�2�0m�0����
��)&�*l�ZF@����Fn������9��SV�����-d���/�u�&�E�c{ �]$*���Lw�iJc������6�o#J�L���(09�7�@ɎA����+�O�4{�ʚ�%�k?�sm���|�d�9 um�� �������:^�.��fT���[|�{���A��+�"��،mS����D#3�֨�#�;M@r'�$$#mwĸ=�Nb>:v�T�'��UB�[p���-c�΢�R6i����[�"��ֆ��N��k,�-�U"V�Y�s���Bѳ�F�R�!Y���,�L�T
0��Upk8�C�r0��˟f��a_^D�ɣ)BɁ��+s�c"WI�x��3AF�����%���=]'n��tQ��l����M�zvT�_N�O���НSw�ZB�J��|50=�1���ᎱW8���J#4�_���0�}gx�q1���N�{�~u�m�Mƫ�4�,u{�CJ8h�Dp�5^?m�+���!���@`~惖�Q?�wQ�M��w!�G��n���O�����k�����v+���<�֛v�7��6�`�dkA�`�n��/E�&��[��fx>���Vv�����c6�8'>�l�l�OpaL�1 �i׳�}y��Fq_ZǴnc��I�F��������]22u �Z��h+���Ĳ�,Ե��_ufB��;�K#����"�,�D{� ���TsY4�lG���^G���w_N ��߻3.{i�$�����2Ձ;���r+N���qX,<OLǃ�g*��Ʌ;�U�e�2��RJ �����_w���l�9#�Ԩ䯌�d�'����k�,�#J+�}֤���(y��NN_�T��+l�{a
h�.����fv����|�u{i<��d!ې�2��|Z���d�r"�$+5M��������Rz:
���`����S��%�-Ֆ �M*m���ha���V�8+O_�G��!�,�A�N�Tб{F�p<�l)��6�:ޚ�%ך��-
������G�J8�ڐw4�f��U]�5�����EU�r��aL�-���2��I�@�Hb�VN}.Uu�>?��q��w���!2?=@�v���;S��'��v�Z�L�����ރ�@��K���-��
����y����d	Ëԋ��#ES�7�T<�Nl��7]�M>酽�'ϗe��|�F�_H�|�����>=��U���T�;��ڌI���
*�8�K'֔�Ĵ0��������
�9P�M�YN;�8���*u�/]D�E��Z�G+�䱝��JiZ�t)^]0�r�E$PS�5�hIs 7�� 5���.KJ�,b^�<}�C�����	T�B�Rt*
8ς���� �.��d�Y�&x�m�ac������ 5﷝�:r���(N������V�s�uzC���.þ�ȓQП3=E-�j���{5�E���c��3=Cͣ�lr���Jx�L��=ھ�l��KDc�,�+��$��{���꺚��c��G��Q�r���Z:�^o��u��!��[%�t�F2�ܱ/�g�a�"��oh��}���_�|ˈdX3��Z�Ё����Ї��_$2u,V���&y��K*ޣ �H�q*�n�w~��H(x�Or���c��bձ�4@ť�:�>�n e�Q��J*�q��0 ����o^�:��ͥڏ�\O!j�"J}��D�1�~r�I9�%����:+0���ﾼi�/���P��#u7�����J��g �Hʪ�(��������-Ӣ��u�H'�7�X2��o
�� ���SLُ*;՜�!%��ڄ H�e|H�,�K���"�c�c'�<:�@pS9���k��~���R]� �j P!D#-��%\���G��(G�Dܩ��i� �a�����Z�2G��t�?��P��w���=���Y%�ED"�3vQ�' �9QQbU�K��bP�
�M%�G��|DJ��q��?My�.�
��ÙW�<N��o�Z9�@w/%��y9c��Gw+B����,S���qH�{F�M�� Y��@�+���z�ǟ��KJٳ�� ��,�]&&8�=3=�� ��%�����5�ޒ}j��G*1}��~��^e�$,����W�'�*H��;�$�@����(y�G9�?�^�ΝF+���ap:i4���Ʊn:�.JG�.�ʑ�6²�����*h �%�.j�r��ဪ<b�\	0�bG3!�(*MZ��a�Ĺ9�vn�:�JI�X���;Ar��E*!��a�<�aY�f�l弾�A�a�Y�R,hj��V��X!�v�ȳf���u�i���K�j�(�����[]��=˳����1�u��`�b�@"jJ�T�Q�߾�=\c��{�l1����7������_���Ȝ� y�=�I���{���D���8����~�O^�?�`��^�\�q E�2���嗏d���!��j�9�����q���'�X���	i-I������h"�Mc��Uz��Tagb�c�P�2R�� HUT? ����rw^_.% �������F��0弑��>�_�v��8[_5]�Cx�cs5~y�&&$�����+�}� 6��Db�o�J�S~E�8��47�uL馄Cc�!�=㘣�F��e�hEl�?)��e�8 �l]������ɇT�XVQwJ��f<��R���ϙ������x�^�`��P�\8OK'�4�n�aB��L�h�2� ��e���h�T&��d�S�
�&��XO@�KZ����t5��z��Gz�m��cv����˙�7"�=�HM�j�_�~�,�Ls��u],3>r��Z2r���0������HuB�}�Pw�;VlM���&&Ka�4�͠�F���EQ���P�c6w�����s]��.�}-�N
:�Xqn�3�ȏ�c︨s6<�4��\�y���U�Nt������9��9�*Ð�v����\������:�+��JNNF���r�w9i���u=�67��07b�Q��rB�ա��C�}�es&�va:'�I�г��k�����;�0��4��W��e��Č��-��={���b*T�Q��+E�� ���#|�oGp�G�j�?��b>F���C��u��ˇ<f�]��gU�W�H�u�4�̀/�Ѩ�Y<OƮ�Т<�������f���c�	��ot�?�r9��x�C������z��)����@Y�ׂNc�ĀY�Z`��}�&�G\�?A{L��;�%�l�3C��rr/�0����:B+���CJ�w�]f��tS�޵z<x�4�C���6/L��4�����}���@�p)��2hƉ�D�{d(b���暹^A%��N5Z4@�S�:~c�����K�9�ZD=�6���5N:���fο#1\wc��b�9�@?�
6`xW�����.��F�8���L���ŉ<�%M'��@��@�nDd2�4�/���;���v��&�!W����0(#�~^���T�\���:��>Sܾ���[�`����(ۜ!v}����c)l����Y��R@b�L�������&M���0��h2
8�_۾�KQ-�`�`_�t��3�,3��9�͗��AҜ	KW��>���ٍ|Q���DnEX�eT�*����g�7�ō�N)�/��cl�TL*�
?+��m�K� �g0��(-�D�z�y$D�@�����#��<6�����/��ϭz�o7_�4t'����@�~D�����8W#j���2��=i��}
U�b����]/���|��HՔ���9���L����EOT��Ձ3V���[a!��l'�Y�M9�,�a�5|��=.�9����ؘ�ۡ��@��/m�_�����]�2r�k�Ѧ�l�]�|u����iV�BL|�jbH�^t��u��,��EY"�<�:�D9�54M]|]�ѓ�e�e�n��%���ƵUM�i�XT�_�O�o��C� "a��+2����+)���v5f��&� �
�Db�*z[%��/����BQ�9~���͡����(��L9�K�4��[�%,a<Q8�:k���[_��6T����?O��ª�Y��Q�[kͿ�����+ǽ���dM��jC*�����/���xuL�-&��=�!��b�8b=�Ƣh*)��H��O�T��;|ՙylN�ϛ��vY��Ry�-L�KruC�[1[V��2��+i��5�©�+��X��V=�0���<�t�n����;Ұ�u�Ϥƿ]P�[���4,)X�������.~� �i��$t�]��˄����G�$����a�CM��ϷHx/�:����L�y����!̆�qx�Ђ F^GO2� T�&t�?��Q�
����"��^�q9�M��EWz�[2�T?FDU$��k̟��/[��S�И�����]������N�nM���"��g����?[��ڂ�i`�̌��R���ٓ$�^�2�-L�������
^g�j{�ٰ[ƙX����;L\P�<� �z *���VX�P#�x,;XYGn?n��$�֋C��8ia������l��Χ�1����3����j|�h��p]F#�$u��>SV'5�,�r��3�29�g6��ⳅ[�K�@֔�9%ڠ�!t~a���QڻWdc��=8��{ꖗ��j�s�en��qS���u�}�!�B�D��'e�{%L�#�B�w�����@T)���#���S;	�ԭ_p�qt�-����e�����x�5�rƉe�:��B��eB��KZ����#�5k�Ĉ5�cDC*��ed8`cy��Q���ee8���a�E��3j2�!$y-/��:��2v�h��F���b�몠@ץ����a�AμD@�[���O�o9W Ȍt�mX�P��&B��Ѿ��Ǩ��b�;-Ųo�$�'�|�!%�0�%۴�R?o�a�_Y,)��� g�������q�Z�{�z����2�[���^l����@�������wf�YD��M��Q�L�m��x&���V�����+�ꉜ}�pC�����SA��	�,_��9[�$�ٴ#���N��yM���}�/k�����s՗��OQ�/P���2��Mk�dtz쿴���2��E���0���e�`z"�%=��M�ڈ���u\""���`P�tŎkSF:�X�:��`h�	�1o�z���;��!�LݵF�V�lI�k��Q�{��rE�����]@��NyU��`�m������=���l���]��Ԣ�9\OB2�O�ש^�5���L�V���lX5�94w�b�t+�p��e����!�`}�������X�dJG��s�Y#��4{�4�r&�L�� � �^:K`ZGp�k��V�'wgA��~���"uK�N�A�Z*}�5ۭ�[Q�_��%{4`_�휥 ��������1�h$���n�rv�dǾ1�uܾ,�~��%ZdU�x5�rU9Y�>KN���x��ez#=;��M0\��������L�˵������B����x���6+����#2�l.�VY�V����3P����� ���(�i��&'���ԇ;��)v�_��B�1O��ȼ(
��9j��TpS�"�KE�8�l��z1@&\�g�]c�� E�jE(��N��A� �~�YFrц�V��![{��d� 5~l����}��JmVв�oz�S�0�&`�Q��K��xtZMԥp4Qt�s����nM���EX%+��߇����=�I��y��\н����k2�Ӻ�\�{�"^�r�pW"U|H�~v��h}w<mE{�[?B
^91Y���O9�}qm�uN���P��;���z^QI[+�����j�=��x��d�ĕ`�x����;٬�����2��9=�2PNM&~�z9�"-C�Bk����X��K��PU�S���� QNC��#��oL��Gx,dD��oրy;*�+p�?^1�T�^M;ʓ�o���ݯ_���o����P��
�J�&��-���Ͼ����N�͎��h�Ez�������n�YX��*w|�Y����f�43��%l���|�V��/z") ����|e��N|))���! �C���͟�%��1��6���DW��Ci�Px5��c������N`��V�����qZ�A�S��hJ+bQw/����@e(�e3/�>��=�k�������d�,��������?9,��j��|�S���)�Vx���f�g,/���@�f��l��_FE]�H�'�b� ���.%1?|��x��xA?�� ��?��+Ŷ�.�su����yr9�������6 ��<g�I0����U�&xP����_%H�H�d�B�|V��2�%�#�~_	1�C3	#��aB+=}4q�����Ԡq�U̫B��i�%��xAy��_P��	��[����*��J&�M,R��X���1p](f(��<c/g�ؽ��Ѿ����[���inXU�jU����Ԩ40F��9�I��%*�ʦ�ϩ
ۧl�ۖ�A�v��z&쓣9��80)#+��:F٩-u^�MQqu;������!v�Gߵ�B�[v]�S�ɿ��3<��s�1�����j;�!`�N&LNj}���d�����1'y���Yӱ�0@׈~�f�w�Đ���mP�^�4�Ϯ<�c�eq����Qñ�p��?b��U9.� PiN����&05���3tt?����XI���#E��JC�E�c���������gS���"x��.mm�ڕ"1�e$d$<�Zr�8��?(�w[�;�ӿ0����M�H쬺���ԐB��x�-XtT�����S�.b�k��qpU�*[��I��g�c�p��$��������.�v�nUND]�;��؟]�*ց/lּ6r�NP7_�B�܀ѐC��F��r�^@�S��Bll���H㬆���l�/��{(F��R��22��@�l��w���3�\�t[k��$���R���~ 5�9(��VG��d����L��[���+Ѓ�Y�q�3������4T�p;�P_�fZ��c��d�0P��� J-�u��6E$����t�E_]����=r+���H��K�h�$E)y���"�OX^u-���6$-�s� ��W�Kd���.��y�N� ۣL��Y^�?�V&|��Ψ�0.�m7�*/p"z�?@��]k�C��#����<CA����%������S���S{������Um��!VY�x�	=A!R��v��;v?D@�/��b�n�P��5��,�5�YP
\2Z��O~��P�L۞��#l�(ؐ�u%
W):�ߵ��iF{X5���ܙ(������ve<"�g��HM�Dӝb&�Z��6��|���b��W8��;�+�H��g#�ߓ�����G{�1�룘��G�M�9F�o0#�W	�x�\������4��^ت-�`aI���;gr��Gd���O�.,���p�O���Q�O�2�ʼkS��
�����Rv�M�@���n�*�0�P��6/o�_1��Շ� �柺s�g��8'��1؁�`�E�>�6����<����@m�Hw�n��RKef�8�-�������v#�2ͼҦa�W��?%�E̾6�1�;�ZJ�Eu{�G�i���C������K�Q�AC���	pwy��qQ?$u%��$$LяԦ�Wm:}��l��ͤ�dF�|������Q�
D-�?�f�o��Nʬ��I����y|�C�_CQ�&�~݀X薶Az�����Rܷ^���������Lx�MY; ��o
a3���W!�J�
T
<dղ/���P�SA��n1⠈�'ӷ�EV�I��Ig|�*Ĵ4��K�f�����*����B^Z-1���ݻ�W�9�(ֺY��:�wp�Z���s��Cz��z2���=�8[̱����� _�Ĝ�n)yu�TDk;��"�]��l��8oIt��ܟA����C5 Mc<q1
�����?+=�q�o�m_�dVA(3�H�&\�j�{�J�%z����h�a�Кm�4$(5UH�ۚ�玵sL�D�Gg�r���HG$qP�r;�:	L�}�ԛ ��|
��q ax-j�J��}�'��WnY����d~C�<����f��c�\v�RQ����(he�㞆�ܮ�C�t����{0��%8��hі����!;rϠC{	j��*�"	)���u���W�u3����Af�Jɗ�����7�=󠧅f�ͼ�s�KM�Ae\���ܤ�T�)��JF����N I(�S �h�8@��ͭ�MAWej�-��j)��� �y����m˚��d� q����-iN��jo��%c"�UoqQl�?
��C�x�.�<�[�k��*QG�}�����5�)�(v I�Z�t��-��мF��wؾ8�eO�T*s[�<(o���z^��VZH����-�P����C��k�V���6_�5[��޻�ɦC@i��D�.^U9�^�?�Y܌�=lI�@���w�y�4-����LE�<��������w.�kP��J��]���\cXʖ+8Q�t2B�"M��T~�޻B%ɺTtH�A���M'�ȷ�w/�!��0���t��lx������_I	�������
|�@��d�#�a��D�CS�ʠ��o_\��-@[I~g��0�`��?�חQ�����	%��AIX*N�tǭ+�~ʾՑY!a�װy�50D�w�u�Eg�ֳ�u�����D�y�Y��QA��d��8������//�I����}%���*���?��Q9�������#��~d����^�(L��}s%���J�^�i��2	  �@�6Y�)D0�Z|6d�*Z���U��T�?Q��M�`r��_�yx{R���)�H#�ެ��]�>d��+k���F�����'��+�S"������C\�ړoR5��H$��Y�b����O�%.N�� H�ZR��n��Q�HX�R��Uh�����������]����{�9�W-�f���"�SI���G��S	DesA5C�w��U ���5���]B|/ahks� s�j��}f�,LĆ$�n��YV$TT91�w`{9�!ɵY�|��#��H����>�i��T�g�Ƨ���.ĩՂ�H$��N1���xr������c�k������Za��Y���:�g6R���6ɕ$�uzg������8][Z��z��ۻAZ)#f`�}��[Ɨ�ཅJ\5{2��9����v��p�|���RS	�!<-���1D	�q*����]�
����Vf������ c�i+ |�Ls�A���������n�[ъtT����ݥ���<����L��-��n���?�R����S+�hpIy�6���	dΖ�^��|��}o�)`�s-٤�u�t%E�ul� �U�t�R��������Xmj���M.=��b]�USZ��Z�o?�[}�X�cBê�.�<T'j����_B����Ӂ������ҕlᒓ��b���Cx�AA'$�m���m��ښ��4���Y�gS��%����t��� ��GK�o�=9����� �������d,��Gǩ_CKU8�>��4k�t��_O�4�4�Ԃ��Vks��]��g�c��`S���������� {z�OL��#����ܶ��J�%�Ðg�<��R��Xx�Z�%T��I�T�J��+;��i9e�@���|_֌u�����x�x�u�l�9�yn��6���T�U��*��p�ypٜ��$�<��.��A6E�C��n�]�4L���zۭ �01\��L�0KF��D;��½�Wz�QfH���l��J��Zd�݋���Y,<�p��������7y�	�`��P�t���y�`Z�*$����cx��`�Vn���a#�A�T%Qy��؀��m��,��'�*��J)%������Qg�vD�A���u��d-��\́�'Lq��j�nf�����/\K,ݠX��z�b������e�%x��&���w2$b[A��$��Fp*�Ȕg��j�Z^J�֤�/0����H}�����x8�P�QI�Y�:��W�3�%Fc'+jNd����z=JH"��H�$������o
i�-1� ~q��qxȾM���<��|ĩ����_��à[�%q ���k@s�ʞ���Ƙ��M
^�(r8u�91uh6)���Z�D�}$C074�S�C�VPOBXŜj s&Ƃ3`���7��"Ey�m��_�氽�UX�d�^wN_t(p! �Ϣh�lR<zkכT܏}���1�"�vA�(��p@`v���Z���0��⇮�T�94�p�!��!�kfu�=�k�tghn��#��_���S�e�2����n�B(F���E�L�@�*��i(�
�!sL���/�;�¹��GS����S��5���N�]p���A�E�"����Nͫl��I{�j�B�e޾ W%)�pz7�ȕX������
�E�݀$�n`!�oD��8���m��6� )W����{f.>�������Du j�6Ÿ�ǒg� ��ʥP�T�����#��[��΋�U�� Q��y_.{:�ˣ�ܽ�v�n
#�M��# �zo��89�x�nrDI�	ȽG����j�����|�H珀3�[�i{+����on��O\���ZbT��3p9;�I���tP���h�Ik�����hq��J9��?ZFx%�+��χ�+1_eB�D�;х���اv�����/��j��'�O��z.t��IիD��Z�}43D���U�j����h_(��`�uT�T)�"&0mTNi�����=f�q@e����u�l�p���H�'4���Gxe����0ꜗ��:	�/Mf�t��Q���T,���/�Ɠ�s��8?伨�E��GB+pyӇ��Z<bC��R�eж��<�S`\�6��
�_�۞��#ÒO���J�(���I5�H|31S��@X�Q����3��<̋��ᨃw��ip��D��\}X��k�[��͔S�D���Z�0��5$k�)�o��f�Ѻ�j,J���,S��܄�mXHat�!�lM��U�\�y�_1���0�N|�ф�ԫ|��t�f��̝�������矿 b���Y�Qj�	vW����]�g�ЀxbΏ1y�mGH�w9X�"ݠ��yj��z.��v��Ɂ�%<IA�b����{��N
D��.yV�l��(�}�{u��R��hHa�H$�/���ĄZ7F�O^�3f8w�*UjNx�����5���2aOV������Wi�ٱ�X#�δ�ۄ�(��tg���H�ͬT��c7����(�&\sn�����]�'S���/�������EW�9�:N�x��ӄ9r=P�#@����ٶ��F#������Ɉ��=#������F�Uj�ɯUݝY�O7�ڮNX�[���4wp@2��KҟD���ұ�ÊF�.��W�����zQ�>k��a麘���9��~��������O;�p��0�0���E���=C�yVCT�ssR#	�4u@��u{7�!��D���<��t
�F�E.x׸�NI?�B����YEv=N��hý�ҾcP��kB�(к+Ј�k*��d��1��w��%�z�<��Ғ}oK,��lYL�i�>���!}{��5.�=�S����/`�$]7t��X{yq�羛�|T7��8��anoD\1yb��y�O���Sp"޹ލYH���d#q��Av�O��"K�&0Ź��|Y�}�H�׫3+� �}�lN]�����y�M��@����D�L�î��aSԽ���1�����5����)��>���ɰ��no��
�Ӭ,�$�Yz\W�Z�0ao���Jd����v�ǘB"4E�D(���=�hlR\˩�7�ߊ�'{�>�t8�5bNݴ��=�0q>�Ƨ���e;���h�Z>���{]7uM?.L��G���b�=���f�̰d��UZ��Att�=zk`�eћ'H���0U�]��bEk���?����q����P<WW�(M��vK�ӑ��b;3��V©C��hG�=�o�� %|�Y/,v�8Rg�z������Ra��Fu���!�?��A���H/),��΍9w9��e.��	J�yzO���]��s��;Km�~�:4����K.7Ͱ��iJ������7�7mU��Yߣ�.l��Q��16�9$n�c� wB�r8�p��Jbb�M�a�~���������s%���@N2�k8#V��| 5��x)˖�n�{ċ����t�I�R�%)ڔ�X����<�FC_�Y([�کy:��L�ϷP�ku��^g�TiP��:�/'�+�r��?����en`T������c&��@Q�LR�F�p��� ��;oTJ��8��䫝g�k���p���5�x[�C� �8IWp_�HW��x�ލB�mUE$�슀��J�S>Pҩx��.��#r"��y�:�T:`VQ��)���u�3bY�l[BQ]�s�1Ga|<VCMvy��Cw�}+^��`�(�G�ɂ38����s��wY�J��R���l�E��Mn����s>en�o\Wc&ø��b�q�@ĩ�+
e�j_�OL�\y�hĄ��d\2C$�}*�sO����vc��{�A��x0.6��b���2RP���:.E�V��ֱ�0��n��%�)�-�`�sk�4�ڒ�{���T
h���P�� ͒��W,�@���:���0P����p�ʮ�� E��_��䕇#�-��u�g)�s�?\%G������~#���Z���#�٘u�Qw�GE5�ĸy�J6f}�M��+�ǅ���R�T4y[09����u/儍Q�!z��\�t���h�l��$�x���}�50�5Ng.�N>�[���1sp�_�^�[�(��| n��0ޣ��%�2�L�=���\i���g�"?�>�c�{ �}�z�:�Q�#�ӉF|�hDJ�|G�p�3DJNL��{�s5�[cI4�s�I�������d���k.�+W:^�!B�H|��z���HB�����;X��]���&�8���2�{pF�@�p��U��T6Vt~��y����)c ��W��W���a�?]u}��l7V�R�!�Bʇ�"����T����I.-�6��0P��>T��QxE����lbѱ�����|�s�I�+U3�3uڏ�omG��eAp����o�yH�DbU�+}u\<ǐiû����^�b�(�O�5=[GP٘L��
�g�y���8�:j/���:	O1�Xm�8�=܀ըM�O׳���2LA�rn���V*��o����#�f&c�H��D�xЬR���3){RH��Dx���:Z�%���-���r���Hf��A�bA���*��x�h؛)O������a�q3l!�q�^��[��~T7}�}X�V:���������	&�w�،�?Mr�ȿ[�a��1F����7��\���Z�|��?���ΐ�N}��{��>��Toh���5{�D�'T|�8T�]�G��@��([�C�J J5s��i�:��	�8>��f������W�j�: þ��[K$�����HY�ō5�"h����,{Q�`��Q�u(�4ŢZfj��5�����7--e�\�p����y�K���f
��7Ѓ>��,"L��>AE/��$��hז����|cG3h��1Y�����8����)J�����u���vM)ݦ͛)�\�Mŗg���2qE�v u�v�;�a`������ ����c ��a(~��J>��� 8C�9w,X.Ke�Nǃ����s��\�!���+��'��Ņdǘ�CF��z2	�����ϒ�~��6�!$��GݞA�e�8Zj�$J�i5�'==�\�q	�^Fu��]����:-����h�ʻP@f�+l$��?7yi<�w2���(�,���Q[����j2\?�M;;���������[Am&�����	���U����T���.\r@/
V�g�])�}��(���%����u&�m�P��m]�~$�]�]�2^�Td(*�e�~�z�p�;��t����PR1�'� ��Ta�豿�	+���ǩ2��@�d�����t!WU����\"���?����`�4w5(ɨ̵(�\I��c}���(r���'oQZ
�h)�_�m�26�Q�=J��X��3r\�ji����3c>qB>f��<U���2l��������tF`M�rB����ZHJ\���*�Q��g��������s��L���Oض����ј?�����ҘɧC���� �2�8{��*Q�|(��)�5+8��y��1om~u����=J�Jf��/��x��."��K�2�厥���'��l�2�k�.۝���+�p�r���	��ꅦ�H��o�E���p6��n�Ĩek�x�ȓ{�j%�Ejt^�`R�av�3���	)��8Q��!�7�yrJr�b��IF�ơ^I4�p����$�Q�[� ?E)���)n��9| ����$@�g�qb�+KӘ+�me��2�6��K~��R��2��h�B�����Q��
��ŔK��c
��������Q�L���G�үz�"`o���s�@�Y�u�����f��~JchW���4`	���s�Ё֍^]�K�m.���e�����$��	������ ,�F�ŶB:�s����| ��7���X�S�A� ��6Vv�%���z�q�f�������N=P�p-C�_<�� ��/[?��Q�z��Gr�ɿ��vʧ�Ƌ�7+i'���6D�?��sK�N�܃��=�z��߂��y��26�����ޅ��UL/v�z۵E��q�9���Rs9g�N�v��ID�ʭe�{��̪�V1�<�ZS(9���8~�o܃q�T��N�>9Q�R#�xǔ�o\�k;B�fpT7����h�S<�����h2�͂��%]���/	uw�Ȕг����2�%�5vϮ��T!bp-�b$�ɓ�g�Fp7�:��[MܺE�����|O���o��l��*�\����
���:YtUJF�.h��q�ؤ�fBqG����e�%�>-����`��H	�2��7X{�D�`��WG�Q��\�ܒ�	��.�t�X�.��gF�=���r�Qzr��?�ub����NbFT�,�ɣ���Z�je.��vL4��۽2nPB0�P �����'롴��
��4u�t3�*��E�F�
�@z�C�b/̻��������"�\4��Ǭ����?ufGD���N��ٴފr?OD�L��4�����`��9�$HS��~�Jd�N��h��@��/��L�Z��Q��*�kDZ�A�����9�4t��Z��f^-�I8ykl��$�L-S�2��는{�нl�d9����"�����������y�H�f\�5�� ;��b�� �o����>AV�)�P�I��/y_�����d��qM ��^m�^�H���|�gS^������<v�e�̐{�h�7����$�XY��X�4�aEw�`�u�C��^���@9mT�$������>�cZHu��/-VK�z��iZٖ���m���7�`,��]�޺��w�[��z��`�+���Ϛ
��(�t�����.�
�ñ8�F$y���B'lĻ����ա�;Q; �#oyǠ�G��w+a�. �a��w5	bv�w�T����I����GW���M��_��q�v�?��?��[	�"�j��Vd��u����Fm�o���?��e��p?�< ŭ�"4�7��_�8�[�Xv���j�ww��<�M�W�����\�����&����3z#�Qъ�uZ ]���*N�'R��=�FULK� ��8�6���XP��=a�08E��S
�o4������v���I���pf	��M �{�`�E��Z*�4�<g�k+9�?^�bz0��6��GWޛ��W����XkjLLj(Оo�Pj$�G�O/xxx�KBɹ-�0�4l\��|�xf9�xr�4�7���/F�[�����v�N�5�*�Z/�/V�S�{5&4s�OW�`o�_��5G�0}���'`��:�_���Ù���8�K�����'����׿�e!�@���f�n�l�>^�ea��̪��5���b��ڒA,(�/kti��\S^v�)ÿ�Z+������;\j}�5䓼Ƴ�Q0
z�3�#���H��!��T�Rá�̣�q��)�sԩ_��?�i����|��i��nq��d낍�q�?��R��=zg��I6�r_��o�0}7��Z�qqx�2�<˶�N%��RK��G�Nu����q��;��S�6E�|4��`/ʖB�x�h+�['��W*̀��7�\��C�'�,䓰{dp���/�C^�O�!����3�ƱXq'h�+z����(�͹Sz�@�|o�*�e�?�>^�\fN��m���.�&'�l}eY������^��hi !�U�>��-?'�����X?�}��Dj�zVV�1(���-MQJx�x��mc��yAͬ�u�������sNllęH�R��x���7d���)�pUC��ۘ��%��Z1��hFx`] ,��J��|3���i�؝������]|�,��җC�0����<��S ���O�ҦSӽ#��7dؖ��L>`.��~'��A��Tk0��h�ê����r
�����s��h�����1��a*��7逄\����;�4���@��?AY��4�`c�}�(te��b�d�I�����ӎY?�qVB���j���2�@Q"�Ǧ�$�k����+��G�i@2�z_`)
Q5$$�7(Bau�w��O��R�&I$_,>K�H��4������iۿ�a�E�X2�~�{$���K�B� �(y1!���S����יϽx'��g�T�Ɯ`:T����������!u���Q!����7A\�a]*؟�/�4T9_�|&P~^�m#�fΝ�����km?��5"���(�Q�u3H[��"��$�p_,��_�#���h	�e��@ghV�atOQ|���ߠe&�9��)!%I�uozB�E�!Q}�j�W:���r"�9�4��45�֋'��S�H
 ��ȁ��~h�E0�/���+�1��˲w��D��h���8��7��z���
�F�n�g��g��ɩ��3�a��+-�{,(£���fX��$��"��'f�� |D�k^ �ȀT�I�(6շ�B��TO���u�;l�.�=�T��k�~jee�/��d>xS�ErD���I������:5�.6�����h�g?�H�[w� ����%G2t��(�x<�B"�Ws�Ҕq��L����i�j�	P*���B�_����
i��)��Ҋj9�r�,�ZX�_�����I�Xu�2�B��m sWW�8{i�}���k��@�p�o�@�KC��FBfuM�D�q�wN�� '�Y�E͗?��螵���{�)T6��z+��]�0N��wrCHQ�D��nk���G�D��N�>)�~��m�JtP��q`���`o���1� �pj�Lq�s�������,�5�Y#�X�2�����[x�M_R&:~��\�B��1�^$ �pLB���k�v3�Zn�SXD��ܖ�U�����-�Sy��� �=����Xs�����)i5�<�C8/�zQR0+��K=&Q�LG�ӴYC����|�&���D��ESގ!�~ �Dü^�Z�P��\�$�vݡ��>�u�6{&��ԛ������7�$��/��lx������J��1uh�$IOr�`&�N���`R���� 4�H�����n�Oq<"�4ŧ����˰c]־;{�4���k���&�ҹ�O���w����bJi�t2}���&s�,<�UG��n���!��S|CP;�����YL��v�A�H���)�FZ(��"D���$�:sEc#���<��Qi���;���gG�i��U�M91,bŮ�(1s��[[����A	S9̳+��j'�{8b\��x�}���.��rp�>�7nst*�:��;R)Iˠ�<Y+����5n�v	����8KW=,���#_u����/3�v�C�t�f�M������rU,F$�3`�,�cs"��{o`�۩V���&?�����f!e�� �rl@���^�mڳ�d��$��l�*�4����B%�"��͗�>G���1#�J(�E$�����w������x{*!H�4^��{��
�H�(1�A�Z�Q��lS�	�d��&v�50��`&&��%�1�i�l�'�@x�KoNν�G�8U�F�!4���0!.����z{Q��QŴ�ΥĽ-e�~��yX������c�eN��Igb/F�q�y��k�7��@�2�{��*��eod�s�-Xw�h�2F;���,�+Wq�dS���^��Q*p�r^ު��S\(� ��0���=�x���!��D{0��D�.�9kU��
��b�������1X,�F�/����ln�'��2���EhxJ��-85j�!^�5ޣ��<w���o�O��b7�����t� ����C4��BO��2ߨo6���9���U5I�'�x�o����	Ry�A�5��]w؂��~��� �0��)l|��k�M5?��O��g�	S\��h%P3�ǋp&{?�k��죁4�~�������7���#���8��I�"4���>qN1���P%^��M�h�M7˩�����[������>%�V�Y�|�(W� 3����D�ՙH�$�
~��Fl��0���/b���WZ��2ˠZ>c�?H���~����z�4�����F؋�����"�8��m+$1�*6D���pL�p�<S�v�ޒb�һ�Cr$c{��}�مg��u�u���m?|������%�iE�Ѱ?R�1��MFLk�tlm�:U3oj���HKL`���:26eH���A0"�O
���wnhkN�m��@�тpdv�K�
?gSo�/RJ��<#4UA�䅽P���/��>&�L��g�P
H�0��~��و~ų���4q3��ix��fndd�CS�[�J��|nE3�אg��oaEE ႃ�K+Whe��繮J5�y":_P��A�p�ZS^9�"H��+���v��7���$(���$?���Ƕr}���
_��D�f�W�%R��q������Ϛ*E\ZDO��`܉:%����|X����ŦfŻOf�ji�-8EG��L��&u�.����gt�a|	l�K�=�O��9��;N~�LK��w��M3,���7�=x˷İ��[;k�.K}���F�9Ӈ��F��7��]�-���h���f���RP��;����D���E���%@[��Ȼ ����ڧK;6����|�['\�����!JQb#�C\�sR
��inz7��ۈ�n[92d$��s�!���sK~مU!_x ���J~�:^��O7���qNC?����d�L���]� �!��l6q5=����/2�?�M�+����ï��3���3��9j-�T㜉 ��F2ђ.�^�z�,�nx�I��`p�XG˨��\Z-9J���|69�C'���/�u����/S��eXV��r앏�jN�A�4�I�L �_��jk����͵5pw�3�.��*��۾���dX�O��OPٸ���]CUW�G�r�:9+Ii��5�C�)-؍�e�J�J����w�q;1�í=J�t�I�NL2 �]�_ȼ���T�4����-z���y���ʎ���A�E����ż����A�@��6hoy��	u��S,�ރSS"��єV����H��הd�Za}B�J)`���,����[1uw���Az$��.`���l�/����bN:�����W_?�4u��'"�ځ����="~~j���+"�9�Mw�[�	K��rY����	g_T�e=7���yF!��
3ʯ�"�*�t��1N���~[�S��ËOg򬖏� ���':S���bZ������{���$�au+�$_�l,f@=QYC����w��OU[1i�P~X�g�"�6={I!�ρ���_9S���D�iߦek�x��ŲL�b��޼f)���r�b%R/�M����`����S4<ҳ݁"�Vի蒤4r��x``���G5V�ǲ�m�{s\T��<t�#d��w	*Nyk)�Յ�����#�&�r6%=�uC�ݶ����a ^�K��s,��:�Q��y6��j�*_cq�/C��@;�y~5Zv!�s�Z�\96���M%�+��HJ���<����O�jF%���[����Z�=U������Rۍ~�ľG���l�i�n@ԗQ8�F�w>���<K^<5��� 2�_��D�j��:�8���x{$����NbX>��s��j�ɢ�3�&�z�7�уp����b p�T�4����=D�ɢ����4ȍ�ʟ'��?~�P���ߐJm�BE��p!��aC9B7F_g�p|�X��S�mU{�y�"ԣh��wp������ndBj�SH���t~ %�|/���+���(�@?�lo�鴝tƇ/�K,Mu����EB�
�Я��/�;�┟c�HX���g�x�i����p*Z�j���r |��wBn�p�	x<�Nc��+���p���j�d�r>���􍉑�j�)	��D�ap�d�����o����J�=���^/d=)X3���@8W) r�� �㎼lcra�p�g⃯�D�t~�`�4�=FT)T��4�FE(���4Y�IVw���v$JǂzI���7��H�0���)dD�]�d�P�8J�����k���5���}@8۲���u��arwA00�����������{q2֑�Uq��B�q	���%�Zv�}i�������eB-���*�Ѝ^6���g����,|�\k��ft�ß��~�3��%��5VS@�kʤƦ��P�95}�;ػ{�'�����SJ��*dr�D^���>�mw,�d���9��Jt	�Վ��R�P�?1i�MN�E'�5ެ}y�~���]�)�&�l�+��dnS�FzS@Gi�YW���N��{���\���y�UdE��v`vVe�:!vJQ���Df��ǣ;{�Kga��x��/Ĳ��;���&�ƁW#�_S5u�z2�E#���u���-U��	V���_~~-��+�?������%I�����l9��䣵����-XS�QfA���b�*��#��-h���'�����#�64�1���Ia��6��qlSοY+}s�L	U�N�f�}e(�?G��Z�v����@}�H���dfvo�I�����>h����G��b͚U^�%	οi\�Z�ǇG���)m�cBbv�K�X5Ὲ"i��Ǫsh�Wd�_ �uh����('�-�h�u�?�뭐��\R��,Sˉ�l��JR*�+#ׁQ`��?ŉq��0�&}�_gRP	���bJ����os��3�<�c��(���&qQ��$j8O5����(���D�av��~"�DYȯov6�+��q�e[�HR[���B3'������a�5�x2<���eh�Sw�l�c:��	��OJ�j�l�O�N�W\w��4%�%�͵��������N���Sm/���n��6���nI Rz��B-5�w����)�q�+�lj�� س�PT�q!S�&̎�>Ӗ�Ӕ���/E�^�S�S�|w����6��Q@b팾�Y���H��)俣�9�i.dK���dۛ��d��1N��&R��[䖗�m<u�7�,J0�s�}:���⢢Ⱦu�P��ьj:�8����`$0Tz}���2�확��|$#F�<�_���Z�r[��Uq�&b`B�5Ԍ:q;Q�y�ک��;Ԏ	*�l#�3�A�y"(\�hJɵ��Y���H������-,�=��R�i;��S>��ę�<�(��8�����|�Ң���smS�>�f���	��I�L���M�hܧ>ﮔy�AI�V/��<;�;2�#�&�j 3�f�"��`�����2E����f��spX��]�}�N4|�O��%;&f�˒Чf�FvY�x]����[�x`jP�	��M����{K{;��#���zQԚ���T��&�r]�1�E�(��1��c{W%�g�����B�h�/H���\�L�	<�x�|E���/	��⤞�Պp)a�\*�P��G�'���k0)��b�/�)3������H�o=�z`YO9rXZ��<c���\�I�c~|�����g/;���� ����_J}'����'e��}K�]����}D�js݀!,�����@YB���ꔀ��.�ڃ��(�E��yfsq�,J�r�z��F,��K���ϛ�3(�׎Q� ��\;H��j��Ϡ��0��uuMM������(��p]���d��_�y�A*����0HO�K��w򺹜�)Ŕ�O�&�)��QZBȵg��y��ʕG�0�)*}��e#m���Vg��E�
�����7�O�3�^��(���_��bq���D^�e�Iz�6�}~4M�͟����hO����c7���_9���,2�R'�~� �t	P��<zy~}�Pr�"Svitm�us������m�7>`>�F��J��]������!NG��m@l�̓������K5�#|�y�ʙ	�_c囦��Ea��!�\���'�����; #>,jH�f�fХ��yF���{{������}s���h�Y ��ٖq*m�gء�=P���n(q� �� }���}���h[�d*|&b����xo�J>T��:��7M.�-��>Q���ye�).�������a�_��ަ�>����v6���1� J|V~��U��W3N<E��M�y�W*�DI�W�F�XʺW� ���7q̺��)+ֻx޶W�p9u7�y��B�YPȾ��(J��*6��ПX�s,��� �o]��=$��`A�]�G�;5�M�-vuC��*�fk#U|X�9]<s*v؟ao��,&�m�2�fnF��9b�~�>djc��,��LN�a��E��"�����<�7B��;&B�>�攔[U!�o�3,�]�j�m�����G�X��� ���r�T[����T����P��$��0o�Ӗ�t�����1e�.G��n�1��`��DSJ���Iau�s�)���)KE��� ��C�6���Ӕk8�s��*��k8Z���U��"�M�	�� -���M=Ub��%u(��[C�ɳ���so�e�l\�t.Ek�1�$��#��+�:���ϨD��u�y|ӄ�AT c����]V�η9,��hx24���=��kI�ц2�ņLb^�F�O+�=q}G����^4!�,�K�,�?�6�J_�x��d�3wq$����!aGp�N����X����'��6#���]�nS�R`I��)a~��>	;�V��f�D�<�W����T Mbt^l��M����W�~���'�,�'7�Mn��4�iW^���d�otw��2ۚ�'��r1@��Gb>_7zo=�d I|�N�����s���7� ���]o�YO�-�-����C�®���N05�rx0b���K#؋]�Q$����O��Ĥ>��~�t�Ѳ��J���
,��U�It��0i������$J��G�W�>�ϥ�	�U��2�Y�P��r҅�v��ο0���8�BH�S�<\���F�2@U@��놆��Nه)^cD��o+�P	"8�Q7���F�������w��M�WE������K!�x�b���_5��Fw��Cr���c`�K���,�϶�&5���.�8�	¬}켉����.�j���ָ�];����ٹ�՟pm�����+������.�W��Ѹ!�T��DéՋ��v��>�1�vG�o]d�Q��e�ᖼ�����y�����|u��;�!�����"�S��lS:�= 1��! ���V;��6g����t�
9�ՕT[��~�և-��;2x��q�L�FW��DB60o��	�ʸ�g�;��g
����3��Փ�QD��i�I�@��DhUn�ܮ�Td����F��nQ����kdy`�.��b5vYb�B9�$�_)`~fw���|iAD-³�e�o�_�n%��0Q�ϕ����(	�z��^�I��~���!O�=eEUC�5��9��[j��{�7�V#��L������bǡL�`l0h7�I�S�a�2�͟~�-{W"���-�O 	&�%p�Ñ�^ �C�s���'M»��:��5���I6`�)�mK�ž�ƹ�ll���⤕R���)�H�m)�Y�N:�mT�� ݱ�K�U��Y�=�Z�,S�M8Odʦ��ł�����赂,!���ey
hMħ�e�5�	�:����7dȎ���ٮA���� 'CT�W�{g��-�^so��HU�=��_��i�<#�����i~yˋ|(�Ja��r~���s��K<d&�6�Fd��x_Q��3ח��ɱ��n�� `���a��+��|<�WZ��h�Z¦h$_���@>B gd�ҏq�W���E>�FW�d`����K���\�n���o��������fg�>1H?<[jM�Ce�@n�Md�#�i���kX߮���@Idřo�vj���IO'n0%�ځڰ���|�6x����p�"z��}�n,x�DK!woG�����G(�&=�;ԧ���BV6��+�U��B�.W ���t��zZ�����GG��'�^i�?����s�Y_\�,����'!�0��R��������fV9�I��)s~e:��jN/����"��O��y��q�Dz���%���^��X�:�X6Ѝ��l*�
�������a�4`�B�E�c�UY3I.��r_3�`�bĥ٣x�S\+g5��X6yY��Z /�b����V�T� �Q/��"b�]zѯ	u�L����[�� =W���FL�5K;�`Ç�dZ'%�둵@]%#�	6fq0\%k=�E�k_, �hߝν\�^S��|Y�-<S�'I�<�	.y�l5�-6_Ǿu���
���L�� ��
�Hsi��/��-��bx����O)��C���<{�V��&4�H���h�@�u!n��l'jШJ��"/�V9[��{|U���1��	��$J<��K��4�Q9
j`u|����nb����M����`Ca���Yve� z����Ng,2>��-��e��ǯ�W��O}6Co�ل���,��yz��a?e�������0�m��K��VT>�.;n���g�j�zp.z�g%�2�P�U�F���*��G�&���|��d�ݘ����J�aN�	W3��� V���J�ku�_�XĒ6��0ݡ�Up ��Ԍb���>��ȟɄ,g�}���mr������z3P�rx��3�3��ԥ%1淔��y%
NPC
���0��M���f`0X�>+�><!˟zMʼ�P�#�`c��w�<0�o���ͷ1�g�N6Q8owF{�y�S�#�h�<���T����n5Ǎ�o�3��Ŭ���,���]�8�����h`2z�r� N6��7Dl����CL� NF*�P�;�A��n�~�+i��7����/�_?W�*Z�� A�C5Ql�f����,�<�8B3L�g(��D�X+�_[��,㓪Y+Ѻ�Y����C���:��A�hsd�z���-<\����v��T�Q����mJ�)��޵�XЬb�EnD�|?�翵��a[&�5�d6�/n��6�f#_��y�|_ ]�p�q�Z�H�^�^�R�}��~Qv�e��tћ#��K��ud�Y����O�wI��{��AC�LE,y=�~�>6.?�)�{�^�Y�Fġ��u�]�4Ļ����U����v����ʾ�k��a2vu���:��L$^��Z�]
t��Y���(_�R������:����9& �%�'oP���6,Q�Ơ���ɲ?����E���yV'�1���?	еs6^��7�z����`S�ܵ� �qF� FW�"T��XN�o����J<Y�ٛ�Qf�ס��$#��@opt�q�����n��`��4��kⴭ����-��mŴ��8ͩ�� 6��t�z(:z��<t�rx��
��4��N^�'t�i�_���`��^���
� N�܎��t7���}\���a�_2E`=�0��,mz3i��
��ZCd�[i92^�Hq_��. )��E׀x��.����������/��u��`H�F7,_�
�P�${�8�ɋ��6w��F#�
��i��#���o�b�D���!0����eC;Bb��$���`_�����UM_�H�%�z�����-��)�����q��'��;�mI��ud@�ϛ|߶�fL�q�>��'�F�	k����x���|2�����Q]#7fׂvq|��=�k�F��fP"�V�.��@�2����mX)&J)�J6
:�������
�d�"���*����w�bm�K�:�	0Q����Zd��tC�r��}0�W~�����Diw;�x��#7�*:u��5@�ː�T�x�֜�7,�E���D���vt�u
�,�iq�+�����fD;�fc
�� (�T���7U��]�����h��J�x>��9�2���ua�.>1?*�A~ա���dd�9).����6B!(E0�b�5�Ǣ��d�Ҝ bMQt��4�%�Pa����i��	���-:wq�����?��(�j=�B+s��6zf�Y�#�u�X�.T��|�m��t �����{b1��m�з�C��O#Yj��d����e�H�P�b�O�mB��%�L���U��8Gu0�zQ����z1Ҁ�v��}d�{���ec`�<V'j��|t�A �nV}���}!PL�,a�L���q����K�G�>~��<8�|��)����t���;�n���.�����0Cs�ո�)�4�_��|*f�71�w�3ca^~�L���^"8@�綗��Sz�EI\�Rq����Tw����I���Kَ�g�(���3|�3��V#|��Mo��g��|έh�p��(�{ɂ�_&��~N<~�����g�.9(FJ���aX��z"�����KY�L����`�9.D�JS���_WސC����P����#`�s}l��)7C̫��D0��v��l�O�G�(�4yB&/�l���C��t�h��B2��yv$bk�-��Y����8�G�p����N"�N��x�*���p���%2%E.�Z�1q͜e����8�)0��쮐P=�7��/01͓�0�A h�?���؉.[p�n�A�4O�-��7���?0�<�5I�x:d��\@e̥О��O��cI���*ɯ8#�5�h�A�4JOt�60U��{�`)B��H�ץT�e��
Y"췍$x��l�߅���K�"�$x�mLw�Hk��d@�����G�&x"�m���#X��&�� �)��1��Ⱥ���M��ˊ!d��J���:�g}D�
�=������?��AX���"��"{%@�)����TGa��_q$��Xx�zހRګ���m���W�efJ�7�U�Ö�����1N�*}�3t��Nͮ	M�����+�;F+�bn�W!<�m��E �)=~EҌ�33�>����'M��A�J��_"�����:�2r �B[4��ie��a��2�}i"�Nɬ��E����9��7S6�XW���%�g��.�]C�7������.��IW5@|�b��r�tU��L)R\�U�����_[%/ª��6À���U��쉦���f��+����'�e}�:�����J�B{���g��O�-�R'�cݻ{�	Ћ�c⢹��-˫��\g�	��LRR{ח����r�	&�v�0,����0Y埕�k̯.T$��h��^G(H��m{�\�S�a�qm�ckW�l��T�3p9���js�<2^x���t��ޡ�4�U�R�,7���P'	��+�[i��ܸ9b���{�jE1��&�F(�e|�q���}Y]�+�}�H���y�gXg��7��GrD=)o�_����ǉp����XN�Vu��ϙ�qމG�A+a�ऺA?��*=�5h&�v�H�G��D��,�f�_t�P�fH�[����D �Q��^�S�L����d�v��;�&�;�~�`)W�L�3�=oX�D��	_���E��+"�o�}�8��&����Q��~��#�Z�z��=�M���y�j)�_�YL9�kC@���T���7�឴e��{0�2�r��:{�>�d��|6V�EX�4�Aɛ.H��ة���֌Ѝ.�i��	�㺅0������0�}O���ΚF�&����]�Iu�_��7Q.�_Z�K}�G8 xֲ�ֈt('��a�P5�%��#k��*Zqv���z�>���K�� �/4��I�8kE�o��o+��9f��l8��j^F��GBE�b�D�*��>�42����DDE�/�~l��H~�l���f`;	"[k����,CS͘�C��������a1�����0.���UnYtn���(�o�aŠg�����	C��X�=}�Z�M�(�G��I�V
l�`���nL�qP���Li��6���&O	Wb_ղ�xdQ�0BU���P��lC���I"��n�ҩ�~���6^�`�z&��2"eU��8�vQ����E�#�H*���4�	��vb���x�������γ���YM��YR�@E���Z$��_�PD��N��^�:1�� �L˥���ظ�A���]�hU�B4K·m������m� _�5��7���>W�h�-wc~���c���`l=��pa�H�<�����*-���x��H�i���	�b�'!o��*z���&j:�@4պ�����F�pD��x������S$܃�>�b@ ]"v��eS�P]�5q���.r^5-��'�2�y(�����-7=p=[�(4�4�}j����Hɜ8Į�V�Z��	0iV��%Ie��C�؉h��(�?�?�����C]	s��:��ђKqb��B��VI�7�奈���ٽ���!{�-��盛I!���-��l�^�6�x��PM}��Aq���Vy�k�b���\�^n���=`s6tLf��I��K�KM_�̻/��=��nf��T��ˋ`�@�$�566�Е�R"�~��h�l��K��(�Pv�K9&��NO3)�3�ۀ�j��V#P`���þT�!��+�c:�	Y{$�<t�~�#�2�����u���	+�"�@���uaa[��O�Sǫ9�4J�Hٽ���i^\�K�xoROx�/nOg1?�',�g���'s�^N�@�6�K]��cS�d�s���P��lG�׸^v����6D�0��f�yt���=Fk���P�|��Vc��3|,�*M�16��Yr���(S����񯢍'����ф74�1!q���M�~�9MgZ��C2��NL:��[)���n��Bn�f����|����oBM���B�����f���8��;��Ѣt��N�+�*T�eMO��(�0mg7>����=��~��v%ʏ)E�)2J��˹��#9A�lO���m#��4�>
-���_��s�e1RK�^� ���Rɦ�#���heś8�F�e9O1HrӑN���q�`�	��*"���f�*�e�jd�O6���&�I�༉�!�i���V�Y�B���-`���L�B��0�����U���Swg"�*��W��n�˳Հ/"�-���G��J�����vc�\���3��`m��@���A��h�^Nl�1�u��bt	]_�Uc�k{�>4�B�&O2y��^� ��b]�E�2L�Ƕ��y>W��������N��-H�P>�����S�9�W�Xh�Y1);�K�������E��02Bo��ln��+��#��>}
����M��V!��v���v� ���IZ�*f���D�"YV"������4D�ՎY&q�B�Tt�zZ��9�����Q�e�&�\Yڪ���]�$�&��b5å����.*bp�Y�)���M���}	�BC��-���i�Uu���&���=�d��$ۺ �|l$�wޢV�"ɬe�ݿ� V\��UD����� �����T���_��4n���Tꜛ�O���*��|DDn�'_��Cl7S���5-r	�:�"c�%�˿)@Dߥ2��E��\K�a쮿N��pJȖ�����r+t��f`؍��bO�+k�(zYO��</��Z�5����S�L_��T�X�#�bb�1l���*o�(a�V,�[jc�{�\����9��]&�"۶1�F�c���{+<��y5���Dԏ�	�;��/�ڽ�Wk�'��2�k�7A�iG�z���=��k��0I��#��]�ѿ����ӓ��y���8�M�*�mR�� s\���]<H�L.D���9Յ!��?��+�r=E�7�%��<dFQ�}~u���>�z��P	! V/��c��S�i��S�>'V�V1���<���f��LH�M	BF:BN8i�����RW�U�I0{�$��� /�K�ˇ��&�?=��uD��ܩ��!Z_�F���h���<������}���ͲnQ���v�V+�ⶫ�il+�����^�$����Di>�<n��j>��oT9P_tn�wx�0��z7B��x��yQ\�,����(��LD�:U��˖6�+h���:�����[�D�?V�"2KAq���/ސ�O�ۈ ���Mk2������A��ޥ�]�,��z����ζt���A=�Jr�a�"�ˇ�����H�O���§��=o_��<9��t�P�/-V('{�!��.h��Q7��]�rO���U�q���;rt��������xa����_�R1Y^R�>I(���Ȱ(�A��
���C�$����_��=Lq��p/v$��v����_���+�i��RRZ�UK��4���+@.���<�&%d�qf.W_	�nT�_ǣ&�ͭØ͜ۊ>u�MA���e
]u����?��O�w�o��VA�+�E� Ww�-4��u�9�wз'\&�E��	1F+�����N�7֒�a�����!;��Z����K���*���l��У���_��T�;�:�?�m���0vZ�r����W'̊����!�#1�jՐ��w�4����Ow�ZÇd��ơ����e�S㚪�,� �����h�����t�IG<,
m�(�m�ew#Ud�����#�b��ZN李*_��i�>~���"�]����c���\=xY�S���}"l��E%$��tr*�YجR�:L 7ϖ~eR�s�v�����H�*�"�H(�)����ԑ����X�Wb׵w�B�ٖ��l�ֹ��L����a��l� �I�/�z5(Yu���e���	e�
�?�Y�L��4r����h���U�%��m���Tʧ�f�FaǇ�<�j.gF�ͭʍw�*G��Dc�ipog�졪�<	���/1z�hb��sj|��W�Őd�>���M9*�tz� )4��/DE���	j�|(@��;����� B�re�K4�l#�ݬo\^&C�:��ELP��=�rHo��G{�4�����c<ѷB6N?��!V�}�7��+Aᬫ�O�#&W,�U�^(`�#@sb�7�!@^��]��}���� \�"�%�G?L�&e�R�]
m��]�ޏ�lҸ��X'��:��|��_>Z��.��z����(ʝE�C���~sD�����$���kĥ�_:l�  F{2�ב�����c�QS�i���p������b���.>�C.@@�Ώm��Q��K�4�JOq�6���X\�s��F<�m=��\��\a���7��Ԥ��=i�bM�E+P��y��
�)������DB�9����J ���h���������I�7��a�^�Vr���$rZ&��Q��='}�#v��=�����g��e�\�6��ܯ(��|4H�H��s;R�PO�� ��B�}���a�u�µz9c+]�������ˤ8�2-49e!�<ge�4�u����eJX�gw��GZ	���]�zƖZ�g֝��_,���v��&U�#7�?̮:/�i./�F��,M�@붼7
��++��{B��?y�Hm71����W�~kN@��TZK�+�Q-%%�A\� 0���\`N�hu�@�t8M�H�w�0H��6�`�����(ݤ��eC������ߕC/['Uv5�>�)�Ѝ�]�����$?yk������0����0�� `w>��o�F(f��b����[>/lE�+���U�W��㖡1�8���|��-�Ms~�N�-�J?�M�=8
�#��M`�S0vr��a?��`D[M��2ʣ:�����a7�\&���i� c�&���W��A���>$kIrdD,�Q�����j�Z!�Of������Ήje%��S3�E�4#Im3¨}��tj �(�_ANAw�P8�ּ2L�(�mN��ܞ�F�ϸ+V� ���'�>���{8��.����<�aYh�@��F����j'z�I1�>�z"��2CTju����嫃�K�	�m��>��ﯡ#�N��"�����Ǉ�H?g&�B�glfn%�*$��/f��b!�`տC�LjX����z��c���\c]�} ��`�Ҁ�
��%� coB�S����`�X�P�X�A�5���'�����w߀�1̟���&B2��%Q��9?�O�R���j�Z����>����u'7�i��\p<��Wh�{c�v`�m��͑c ����06��Pa��*699�])P�^\�@��Ґ����m@$�h���:���(M�-m�20a��f�I2��>X�GYd pöc�^���������Te�_�%��o�.u�}���r�P�Q��%ާ���L��Cr� � f�x:K����!�>ٞZL5�D�� \���MEu��H�j"Pq��N"�ͬw�]j�y��)�N:psj�9���O�Q4ޜʝ�p����TW��"H�u���4�4��U$��.QД:4��݋.��72��zN�q+�O5ܾ��*ٹF����Bm�38�bգA� �#�T2���~ dd2S�:���s�5r���A�_3&O0����t���V��	jɃ�
�Z^-Uwg���l�]�7��mBDy&~(ͶW"�~����ʌf�}��nE���&��(�k�H3b�&�&�h�A��lZ�w�Ji����� �z�qL�}�<���;�Q~MLµ]q��$���6�磲]\8�ձ�2f.��vT}�&�]w7k�z$�M]B ����:���4�K(����W���_S���G!&��<̫�g�����g���=o}��
�ߧ�i���RH�~?tj	��'�
�9����?1���h�ްj1���t{�D�)��~��^5+����Z�A�ƥ�0�� ��dumO�X���#N���;U��bs�m,T�ɧ7�i���ac�\��J5I�ھ��wK깊4�]϶�uS��ޖ�����n��W	����zʱF�V�3(��� ˈc����&k ф�������,L�x�g07gk�p���+��Q����Ey]Bg��L�_z��Bz�(mަD��� �h�o���Զ�t�x�2�͌��Y�7u��O#�Pf�z���@�%�b݁��ɑ�T�JA�_ɨQÂd�*�+�
��甡E�C�;��,�O�V߷c����I�Y8f���v�8�����A�U:Ͼ#5��xƨs�	Xc���u�(�}��<|@�R҂��y�B擙V�(;Kf�z'���v}ﵖ8Dq��Nj�-1~#=7�4�Zvd�㪄���@��9	���]meVL��|=�F6������0)MQ8�R��*!0)-N�%G���o�JVM;��+tR�i��^ˤ����m`�$�w�uW�eV,� �Y(-(�:�K�8����X	���^�PU�R��Z�1'M,<0X���i+9-�o-��^��s��K&w�u���;���Ƣ��k�l$^�1�Û�Do9e�6 A t��X�	Ť��m��dRپ��Tow����p��y�@�՝�(}Y	L5:��#��JȚȟ���b����-�8-��blg���W_�'��mԱѸ�(Jcn�{tʮ�ZB����C�r���`K )��2��c��T���O�EP�P����F��/��´Ļ*D���}9}�vGx\U�&��~�Fא��K�:��&o|o������@t�'p�|8�z��-�uO�m�*��8g9�_h��E��˚��yG_$�)]�lPx��4�G���(�3� �L4�ula����:ub~g*��8���F[�驷����C��P�S��:����c�qt��J>m>���0q0/���A28P2ۊ 3�-��01'XwB =�k�V�xsn��ǎ�~#'4�5H/ܚ�O�J��$��#n�v�R� VX�r�J�[(C�Ҧb��a�s;�����
weե|r�ހ`�|P�p��i%���D��f�\q*&���!pK�w>��ō»f���ň�oB� C:
e�}w�h1�d`Ǖ�MV���|\n@J�j�:��Z���O��o�1e��������6��/�9��(w�\;��boi::����d�p=Q�s�q���[�M�����*�vNy�]�'͆q�#Vl�\�+��K��H*�?��ݚ�u�lň�8��v�:I��>r�[�����4}��Z�������E<���֤�!.<�n�&�[��qh�O8�����MR"��BA\��<D�F�wkB��I^">o��;𑶇V��ʛ�p�s����YgAob��Tq���&���L���ɕc��lbR���d.�ǥ	��-B@�[������W��?;�sB,m�~�"q>V����p��@��4�`;I�IĆ˓�� W���u��p�ư�ƿ�ѥdRQ8�x`���;?��eztE��JX3��"�|v�3O���Ⱦ��p
�����s@�
���{cl�L<>��&�>�}��	oI+�?��F���T���3���I���̡�D��}��/]m��ū��,E�y�h�v���S�8b�-;zm���V�R�W���5�l�VMƩak�j�78d���M�Czu���^���A+���KQ��gc{b,%{���=O��@���.Gm���7�8ԳQ���W���r�p����|V�U�P�q�-W��݀�(Cw��i�7#�����3�5�%sm�I0�8K+s�ס`��&������[�JI�ə6�xU�1zi���o��p;O/@_���dJ�G�u)�>ۢO�@��o�P^,�iϣmLR: �S^.��툒�&����(0"�.:ϔ���6�>�w���&��Pv�r��CI-H��l&a�L�����J�S	��I:v�*7���w#$K>�r�k��sa�SW	�"ڣw�s�KPg����A�u���������Mj%n�ni裒�������u;Ƴ��óC;���\wkը ���y�	\��&Mxb3�Kq.O��gܴ�^3��5�η�eEu�?�g�)`�3��&rJc�؅����]h�B����̵OHo-�O~J�a��o������rI�׵��˶�}��yc0|1T��K���b+H�*�mo�'Z����$E����5�g[g���$F����߅�U� /�e�����d��?��-��%�)/�f%GVSpQ��}��T7�o�e��p��N�[S�+s	��$�yP�N�	-��w����˱i�٩����CV=)�`Ŕ����j��	6��Q�����ɵ��m�d�)1�\2���헔�3,��X���*��=`~���$�^��9������,.<�9���e�ߪ��6܀gi9�)�<_��d��5����G+��))5��M�,�]z�'��<���>�SrF%p�,����Jr���5Osr��R�䓯�Ku��94��F��m՚l�?�:�@T?_�v$�:O������7� ��&B�RR/�W����B�7ž�+��^��ؓ�b�A�&��U�rݷ�|��b���:,nB4�]�9��9���'+�4"	�֊-�/��Y��b6ଙ�	��A,(��^zz�m%����|F����5m�ʦ���}UC7��Y!�����?y޶�_�p��J!�O�u?z^6�'��_���3����?f��e�Z�	�(�5�*e�s��9��/!a#��W@n��ૢA����|@]�C��!>�jf�J����=�Dy$�t�gm%�ĝ�&o*�a�ҝ>>P�0�;e1-�Y�^�6�~@ڎvO=�7`�[x)a���;�,e�����t�CI�\�&ﶴ�D�:;^�fO1\] *u�E\ŧ��!B��QY:���M|���R+����#J�%�>EP\��}%]]�G�lp��'�7`J�g�ʞm�Vc�,�,b����wC��f:��a
O�!I����sH�Lw��VQ�{k�g���+�$��f|j�r���k�p&C���guJ�u��EB��7��]�Y/]�۪���Q|����|��@�.U=b�}'����ь&8@}xid?s�0�ނ��z�.M��3ڕ���1T�в��V3�-���#��W+|1��y�ORsu+���o]Flv_Cn8�3}�`֓`R÷~�I�9i����Z��I�q�J.���.e������3C���;K.[�U�P��8�H�b(�1.JG,�%���8Ra;	#��qu�UJ��`��JT��������yr�:IPr�;5c�D23��B6�M[ߍh��k0�5�u��w�8�|���%��<����u�RbcZ�N+yΐ6&���m�O���VXĹ�fB�ɸ���k'��H��1�	F��M�Љ}�3�<�_�~�ë�<���r�/ �M���e����^�$���}���^G?���
��?d�_�n��BC��a�0_��£$&/>��~��ۨ�{`d�҄f���{��1�(�>�3���3�����zm�"��J"rG�$4:��X�T�:_�Tǵ$����օA%W �پ��'A#.�+]w3��H(�d8��>�k2��>]�^��Ƅ}����v�E4�
֨�l������ecN�CGá�auo�����/f���	��c��F<V�v�`�[;e)��h��*�{R鈎	-�Pə-*K&��x��m�z���#��N��X����Mg�d������b�q�4P��Y˼=>���]ׇa۰��\�8=~SaB�xWdKz�V�K��>��M,�hȊH���j�#���,�����)��ƅ�'#$�0�	�,�V>pоxQЍ�[���4ڲ�޶}К3�7��l/6���E��6'�YG�TQ�ǽ���MU���UH�;�n���Z�
����1�d�uAƀ�	]z�o��CH�%� x:Z�(�_�h�$R�V�����)�?�
I,j���]?Am����k�ՖKw.�3�
�8��b�F}Jq��V��`W�н@��2R�|GRFor3	c�{��᫓�D��X�?	vp;?q��ݯ�EH��Lre/fIB�3�Q���ds�6��NY�ّ��L��l,$A˨��ǻ@'�n���ǧ�<��'���wj�\?�{��1��K,�:�ؓ��Gx	�\~��5�(.��O8	�(�&���*砗kx��y��aD_��g'��@"�Q̟UU-���/@�&%�dN*/,[���F~\��m���ǜ�	�oN��O6�7��IfI6gN/�7��A�����(;�{L��VN�/��va�qނ���{i�]}e?j �4V�hM'r�h���jZ��w�И;&�C��c�t�?��QĿ3=8�I
�S�ҵ����+lT�d��"��|Bߓ�l`��g������	Z�+@��vj��]�q\�u��l��	�] �0��7��k�tB�_H��Of�g��~5���K�j����zƳ�=U��������Cx����=YN�I�=�v�j|��W�N��Ȉ�Q��)�/����޵	�����t�v�r4�&���ｱo�l���9�iڸ/�Jg��-�\#5���F�c窩�r��j#����5�٭\���9ߋ%���p��'�U���q�5�kѬR��:����G�1�\	M�Rb.H�n��_�~#�����;3�z²z��\�L }E$�/z)���Y��/�����J9Ì.
ޢ��KK!(��O��䕡��I۞`Y���<p��t�B�\�+�^�Z}W����}�P�H����&�6&�u�_-N0��Y.��Ԕ� %�xʲja��i�^�D��&Mb�*\bAd!�\�
��Dx�2+���[����%(J�4H�9��[n�qv>}}�Fr�bSBW(A��J"^��
֔?�"�)�iLh��5��]%�,���h6q�
�&���cK������&�)~f��7S֢S��x���U3�����k?Bs�:cΌ��ƌ�$�r�2�h(<3�1��%���e aS���G,�?�:��TIr���٥,�-%�-6���1.oI�6)as���ֿ*��;�ib�wS^�H����Y������%�u�_ko��J9q���,��A�U��u��l]�A��bm5fc2r����=�t�0�c(��eX��?K� M�+Ѱs ��2���ȡ�E��0��?mӚy��	dS�᳭#U��G�b��kT�����$�ScW]�z�֦͘}�AK����6�aN���l6��d�������A�Ja�.���B� c��ϔG��f�7R*!�+�Te/ !�N��=a�%��ܢ���A:ť�>Z����;��[����]ș?\+�a��}�b\Z�PHaI��雊�'493Mqb_�P�%B�Q��e+���r�oWFG�$��nA�Tn��Aᵯz-ڋ}���Gu|N	�]l�B������9�i��9F������׺ON�>(��\HN��R���4��f�o�cd���TODSS}�l1�o2� ���X�U�7!�WzO�;�<�/2��Ba�P���ȶQ���bq򿇂���\���{ɒk���>Ђ)�p�٩7��ϻ�v?�E����˰��qJ�WZ:�H>��Q�;�%	:�ɿ��
$����~�F#�M�cK|��d� V���.�K�W���(1L�,��+ݘ[���)n������%4&+:J�P��u�Az%�cK/N.���Z��H ��ku�v���zAG"/�𓬾M�=�A�@�M'��"�`JZgU[i9X&@lYA|�A�|�7Gt���iL�^9�SZ��E푤^#�r(Mt䕊/���� ��虒]����E�w�_vn16:L�3��4X@{ ��Z���6��(I:���挐�=-SpqBӆ ���\��sÆ����@`M�G���vu�o��+��hN,��j��u��X�P����p��\߁έmb��j,4��|��=��^T��ot.w�gXf��&��;�u�\����%���~.򦘔�12&ZX�O�2n���6}l�����Ux��u�!D�	�y^ZD�f=
d���[vK���n��z���+��r�L�ɺ
e^7˒�QC����p�b�Vk�	�ϻ�^y������x�ο*y�����蹥*���b��������49;R�$G���-f�ϻ�;�sE1{+n%j�8�,�_e��~�-n�#������TU�r��c�N�k����L�h��]���
||\10�U�QC��z��ٝ(�d
J�E4lg���I�Q��zu�fw5���[�͝ڥz�D#�-i"� �#RY�	�,FhK3����{�\ O�s�t��T�IM�%�ړ4�фJ��~�����:[z����t������䌕�i8�i~)ҡ~
K�&1cg���IZO�V��Q�6���x|��2��U�Vc�Y����@o�m9�B�{�KMU�sG��Ià՜��{7s��S2e�����>�OIN��e+�y@{�G@���If�{�����RzG�R��L/y�]񜍇I��l:��2��w�[���R�j1U'��^���x�~9@�.U��Ý��v�ѝ_*�˿�/p6W�m�TQOZ#L�'N+Ҝ�x��W:ig�|��	S�̋��f�~u��.��l%�Y�l�H/Л&<4���{�<sf����0v��N/M���q!�L�O;Ӧ� �ئE�J�?ΰ��+ɡ�T	��-���&��,Ln��aa"��F�� UIB5�i_ɘ��L=�_)
��|��Aٴ��#�/�� ,ڶ���������!۠�ُ?��>��V�L>Z`-�	�@�m��!�FK̡CH0P�6�Qb��T[�x���2:�8�.K�qTm�|:�̌�����m!�>v���A&yĄݷ�����͈_d��^b8�`@�o�L�*�r�9�F�:f��Ӛ;I� �	rn�n��/X�^(�=�Q����([�-��W~�C��@��JkƔ|$/O|�YYV��TG3��nz�G�T%c��F{��1%�����Q]U��"5��Ү)���e�Q�3n=Q �G�1�}b�%2�a��L]q��$g��?�n7g,�����$P<�Q��	lI�V#���0�����b�������"a��l��в\rBT7�O[�.'"������;�TF*���<������}��=�5�ym�m��K|�uTI��\�Y���f7�7`T��YՈ�`xjCr�kt��бV���%�� =�y�L�{!1���P�t P��뛾uBo�ə��Y��~b�o�V�D������	l2:� �2��2�d�+��0O$�X8�>ǧ���[b��'�����V%����z�YN@��Z�ʁ;�Aʍuj�o��'T���so�R��tM������� fD`ľ~�V{��GO2���&#��3�s�M������Fo� =,ϝ�w2�-%iQt�� iW�ـ|�����b�31���/��Jyk�<T)H^�����%1����3��_Lj*��~4���q31N�P���g�a]?��3{(��ow ��:(�S�M;�?�n���Eu�xl�Jn�v�_tx� �T^z��G��)��=��0b��� i`7�Qv�Ĥ�}��,f�ʑ�V��)�~�J {"���<nT!�\��T���ѴcXK��ޜ���N��VHl-�<a�Ͷ���/�Z=�[)ޭ�7�>�\���$~�� �p�b��:%4>���ox`��ܯx���M�J3\Y��e�4o�PE|)2:'W6�O�n���c�#�g�m��V��rNV��N�;���~��Qaʦa}���z�u����K�翥cI���#S5��A�?��D\����/[�Xۙ��~[�� zOހ�I�T���r����T��v�Ͳ�CAw$������&��l��,�1	p�1>6��i���vV߬�t��#�P<��N`��M�ړ��áu��mBo���ZC@��fY��7��S%���)2�2"X[h$R�T��7�<�(QMԱP�_>�KaQnL@��P-��DϠ�H�U~����$�6��ҰAy`�$�����P�9�d5�����Őׇ��Oc���
�0/����t�ݫ�𩎫7�y�)�����5'����c�`����C:.��\�ߝ��T~��=��}�{#��y9ݣB���]�p�_j�n���f��D�zS�K^�c�)HR�O�S�v�I��%=Ȯ�{}C^��.�(v����)�:�W;���g"i�bu���*�� ��@ ���#i�M��h6���������U>�1;?>UȰ��r0F7=�����}<Y�$A�]�ZD�Я��ݕ��a
�УJ�(O��(�����5B��[̳ʽ����	Qw�e�4u���Zh!���`� �����E1ʋ�o�� ��c��_�+��wf�$��b�T,��	����Y�t�����G�F���8UX����a�,�(P�/���(�ui1H������"��
ph��r_��׎��jEl�<Z���"9�:ڋ����O�.�!>���<�U��3(�<H~�Y.H4U��t��Lӳ �����(��Y��@�����ͨE�%]t����ܭh����)%��P��E*v0ĝ���pBŏ9�?<|Xy����ՍF��3�s�jv�?�]�{�3�D���+�Nq~g��U�����L�u��&���
�����/`��G��+L9����7�rMn���&��]�� 3%%H���U�	������|��>�R7�&pPM�c��o��v��7N!��xE�;�mC�F�pt <^��t�1��r��ౠ��ܩ?�>���7��S�7U��$�xJ�K�$��XZ%�)%m�P*�ݭ��6Q���"�<a>[� �{t��RȲ�$+z���5�]��ۣs}=��\�+S���)]�]�z�ڊ�#��:�͕���[ڷD����`w�0t�4���"�p��8q �yG�O���)v3*�6}����@-�Fp��#����Fv;T&s�����2���F�#�vC�-23��ǽ�Y~Z�%���5���U�����4?u$�B��e]�!�v�r�8H�S�Nq�P����I<�S��_1�cAU ���7�}�t$���n�U�M4Z�������̯�����w ��~�8�G�q�N������	Ժd오�m��+I�wu�v\�@ -.d�:�gU��!d���"���3��@��*����Z����%Y�@��Ah�蠮��8�'I�[�֬Ia���a�fi'JD��͈$�Ojr�������5B|��+Z�C@�yO���k9�F���?Q�W4d=)�����WbGJ�d�/��(:#@���KǍz�Sl��Qg�%�(?�����}}Z:5HyJ�d��Wxs�{���~�Ԍ�CZÖ�caE�w��2��,����ڵzǽ���2{� *�����sQ��R�I�4��-k�^~����+Ncp��ԓ�������^��q��Y_%�hs�<i��J���eѾ�|>�t�?)Z�1f�A�$~s<��)�*i�ųO ��xk��o Lk��5孓��˛�ɽ4Wh�i�i�*/U�;x�'4x��v!ѾD�p��o2���4q�5��"��'� ����%jy����� iD��p�&��/����>�۔~������,� ��t����b�~bWe^��܃(�2j�٣��~r�Pd^��W+h�|��¤e'/���n>�ݢ��(�D(t�A�)�V�7��I��n_3	9��PU*��>��T�L����&���DC9d_����)ꉴ4�#���29v%[l�VxU�r�7���c�ɐA7����Z�R�Ï�AJzM���-�F%�@SE'�-i~�g\�^-�2󞂦�Y��>����,
�S�v&��BrN���:�-E�]�Ði��O�G���M2��d�y{y9���_fq��X���v\�wR�@��"/�2���%	P"�� �,C���M����?Q�{���G}������Ǯ�!i��!u����'�=c�"���@~6��-54��-ɾ�O�����u�˖�5��,^�=�\�Q�o3��L���C�o�
�P>St���q��>�e�Mu,���'�����~�Nk�L	n־���L�@�B�U0�9"G(s�U�
��>1>uD�=>��֪�3���pH���-.
���? ~�9dI�X%����*ȟ�:�8Mn<�rĖ�8Ib�ZN��J����������v<�(�L�8�p�+���k� ga�T�ϋuc���q�̊�uL%O�>a�}y��PNd��s��?ף2��:����� �X� b�`5>��o����T�.��I�^7P�����Z����V�m~!�X;���jH�%of��	�$�ti����*����iM�o$/b�q����T�&��ex�-�80�v�`�>�
�zs���3F}��I�Qi*�����㾣�8��>�Ж`G���W�m�E������4l�B� �˔ ����6ߘ�#|�l่��NsKo�e� H(�A�RN5b��߯AӟR7��*B#+�}�.3��`ؒ�6_�?�A4Xȗ��[Y���G�@�1?�3-׈Ĩ`�F�[���m�M��q	��	�nT|��
L�]�
�+�9%�R02���xK�'M���\�1���ũ��ݯD]�w$E^����LH����ˉ��>����~�F��(��޼�B�R惼�P��@��t�#���9��\RW��-�l�X���lf�!24���ߖ?���3ɒ�j���K���	�n�2��@�u��T��daLڝ
�����>�\��g��aY�k� ��t�*(`�~�m�O4��k,"�n���c(�К��F�fX>Lo`���Q���L���k���?����x3�#k%FM�ZpI�ġ�ĭS1�m�:��Ö%�ݤk�����M"�XcC񐱹�j�

�s���B���w�T����$�� �ʭX.'0򜊍ֲ�hA�H)�5��3���5Mb�I����X��U$�io*���Q���;Q���d�X�12$
^�d��ع��ՇT�e���>K3�*��`�#/�O�Q �` ��L�FRK]37Z�U�����T��s�͋"M�I> N�I"�]��1*��c!�.�<�����`�l��a��,��OJ&ޙ�2�rmGQ��;������7���%z��]0���iB;Syi6����<�����ЭY��)w��Z�}��0@Y4A���25�0+"�M�Q�H�ڗK,tfJ�;��И���g������x9N��A��Zn���G�xYL����d;?��)�E�33�E��4^�F�����6�u�'�����BdN���g�H�(�F�a£���n�h�R�"���y��-�����T䥛�o�^$�N2����R������WX}��T=j���w��On0��g���[<���^��6��d/�3r�%���*����_;"v���}J��^��m��ǠP�zbL�p���*e@ا�X���uG����i첒�af;+H�Oq4Y'>z䡐�?���gl�{۞^A��j'\���%�-�7�L`�vl���O�6�1i��G����h��^�<���Ք�{j�
� �wr6��XbN	k@	���y�b����0�c|_���8�a����/`�M�.q�=%2C������q%��Q|�97�9(R�C��?�Mƞ�[ֆ׹K��-�+�x�J$kY�u)7���ul]�A6�����^�غ
���d
�p���n�,�M���
}��WR����t1`]�����ɟ^���*_V�>)F�vV�֘O�皧h0��_E�^���&z<9�͔��^U�6�G����n��D#|U�q��k�?��� �,<ܨ��yΨ>�㧾,*�S�.{�B��%�w�E�4G����.�;��;�h3��;�4j�	�@L���>.	'Q���ݛ���Zo�$:�mk�yA�h xl�z�\�?C�pސq]����%8_
�)�):5�<"�iV������O� �5��ߏ�� X#45]�Bw�y�^�2I���@SP����J��g�������jý�PNKI��I�Ts�\��6����I)�;�aO��]��[9L;"��N�y�+��%�;�J����s���L�
oG� ��E<���{���#:7�ݪE�h�	��ȰȺ�0��Z�`�pZ�Z��#�Dˋkl�9��ݓ���`��Q���4w/��FL�WQp'c��+dP�P��CG:�"9ky{�$���r��0�z�]�.��!�2�Z)	�Fì_A��1�R~ �Z{��ۃv���6�O��0����4�ĐŽ�m����ث��{v=u���˙��(��q�G���C�No/$ʡ�*�� ��L>���A�+=<��1{��HP[�_ۈm�9�"������b��nK�xu0����^��<������y"�$�:R�ջ�gDcգ3#�#�͐��'C"�7%6�q'w��g��a�А�������2��,���G&�H�}!|T�qgI<��{�b�^P�M-���w]J~��y6b�GBXz�е7����	l�ei���ի6�"˸J�}�0Z+����E�\�����5�o��jk����Fw|7�Eg��Z����g���H��ZV���X7�G�-�Zo{�^%�>�t����ܵ��>*��o�����mQN��)����wp�r{�7j��5� _�����:�(�)�'��d����HTJ�6���%��~7(k���g+laG�zݍ \�6���RE�aLZ��^45��)ʸ��͇�mOr��s���\P�k
�^\�;���S��>� ^P�>��ċ����n�U����n|�$��<�Z�E"*�F�cZ�M�� iu	O�Ä�,��5C���ｎ��s^��v�?牅�6s�*:�փ��?��a�o���}NEj.6��w!4�n��P+�.>o�e�50�����z���U�Y	��뽯�,���&S��� Y,l��z�_�x/9E�(�|a�?	d���n$[v&��}5ZJSTf�n���-�U���'pVD��+��f
�a>c�ڒlLiyP32� T�H:�Y��(�<݀����U>�xŇ���S�!09�^`�o�?������+��x��-ъ�c<ѻY������s�~���IXPB��|�-8���.j�+1�>s0�"��s�:=b��,��M��'P#�V�q$�q�9{vDޤjZ�5t���嫋jД����u��j�桛m��a��Y������P�,Z��V�<����:G�St+Ne �n��M�A��i�rN��0?W�1p��a��[w.:��������8��{�Ϸ(E�f��
\=�&���tr�6N�~S�X8Dٍ�/���^X���R�~ྉoA,gg��&�=[�a�#wr����B��V���ב������!��X6h�1I4����%�8�E
3�8���e�J��i?�����퇆���[��c3��\����"���=�A�L[v�@p��i�I|r��F�+���tVX���Ȍ�i��k!��� ��i0eg��o\� �g�L�?-i��tn�] *�%!l���1��FbG�"��zZ��0�e�� W�*	���Cm�"�*�Қ��0�t��!
߼bc�El��CA����8Ւb�������R��`P�+:���	���ۯ@f�z�`��M#I��6��C_��4��HM>�ݶ��@tj7l�,4�AF��6m�
J}��Z�XR��X�cY�6Z��t0q��3kAUS�K�&bӓwq�WP�.�w=�6ܻ�`��ىv[ka�҃i���v�
�1S 
gD9��{,YB�kD�m�9�n��ra8�!��gB'hMIfUg1;��M�g�`��������.��}U�ͧ�#6��dzS��+�&U��!�;ۣL�c0������ :`/��d�����/��@�kɝ_K@�O�$1X�=ߎ3KR�� ���P�2ƒ޷�%���f=��{��לx��4����^y�z�Ӝ��,�n���!w
]�kz�Ľr�j���sl�R�����s�nR^��2��hq��ځ�HJ��� ���-����x���`����sw��{��FL8��riqo�p0%��Gș�����T��G��e����x���,����-�!�/JG͌�p�:��T\ч��<�#�	���$~X��ݚ��O+/U�:�8��u�G�]n�'V�LWۉ�X~���?�NӮp�����u���,��o��ݦ-�|���l�������g��N�vi��_�aPG�6k%��b��s�*|9P���vl�!���	�[-E��.!�Fp�'��"0��FT��
����W~L�*h(��;��U���s?�	ƻ�E�,mӞw���2�XXk-u�aCؚ���El���Rs	;o��� ��0]��:� �A�&7<Z��"z��W��ٓd�Oe������AO�"Z`���j �ݗ�͒�KX���4 �p�Ԍ,�pI�m�J^���n�z�L�� 	�1)����t�к���e�	��kB�c�;*�� eS{y���j�������
h@f�{6ɐ&��}�;����'��顃��W|�BOm������҇O��Ev�QԴi���n'��%���x��>� O�vp��^�r���4v��A�7�WA{#=�З����7;Mg��i�f<�������n"ԍ�̿f�$���(��)v��{y{Mغ"����e�`ξ	��f~U�� <�C�~�4��â�e{q|24��Z֟c!�f$\�af+��
�(ܬ|� B#)Eף& qۋ�E�"U�>��R�}��xWm�-���lK��]��KT3]�qb��'Ҍ��H�����%G�ȃ��!q{�+�L��I���Z��:�����2�%��lú����d���|Q��c����+�31n/E���/\ �
l*t�	��OH��8�ݒXv�������C��ce���D*}�\��|����Cfޘ#��Ru��]�~�˖�?|J���o��c7߆��9M�.Y5�����s��MQUk F��~���e؜����-���G���߶�zAK�����8����;��U�U(~m��&�,� `���<�9�\g3z,7���K"����U"��f�'�Co��u���}�{�rNX�$.�/�}�$6SB�̺��G�^�
,�y�ӄd�����'�V�:�����H���������6	�
��Ss�4�ߞ�P�0��ۖ�
=F�*�(t#�2O���g�Z�rM�,�� >&�ڔ?���(�����rJ�6x��~���?)�q
�~]:W���l�ݐ �C���1�hb��j�4���/	�R��uP�9Μ�|M�N�m*���Gl�.�3b��6��=fC�%b����	)��ɪ�g�a*~�Y¡�.[c��Huv��b �C�2����֡�O�j�-�h,�O�tm/r��;|�0;�ðS�D��we}������z"xHq�1Vӗ�?D ��ƞ����O�l�)���d�pd��:����*�Ȉl�:����ؤ�!eV�V��`��AP{���)���jY�3/��ٌ3�i��T��\:a!����������쾶����&?����\� �;�\�Ѝބ(�c���x�zqW�Pj��%g��� oɇ��DW�#�P$�����^�ƀ�f��&![�����a�e�Y�I���
����9�h\q��L��B�v���nC  ���$��`����Z#���/X���)�Mo��g|�&"BF;������Ư �	�����ƙj\��k�{uF�9B�ϒ�6��vߡ��y�b�����&�FX%m�e����ó�j�f�Bҏ��}�[�j�QU��l����B��Q��ߌu�ś�aS/�f����6P7Q��~�f��!��N��興��ٹ1��ϰ2]�"a�80֜�o���Ћ������R<y'��3:t<P[�ɇ?>�ZG���=V�wh5+dW´*��Du}-�be*HgoNO	�?&u[�0���*'ܬ{�$��ma"X[����X=g���)�����F��d��D(Y��+I��ƹˢ�����=~.6�J]��:;㟋:���?�҂�f�JI�%�'����.P6r89���<`ɽ�S���?<���t�Tv�?��x��t���A�$�#�.bP�q�l�7��`�~k�����㰤8�q��_PI�w`��>F�R�JS�����vč�L&�.�I�M��A�2�Gb��L�A��y�]�+\�%Q�xN���o���,�✳C���ʛ��������R[��5��ӓ��=�dK���b��	�[5뙕���_",nˬ/?u(gLb����8*�<�C&�0;\ȥ��d�g^�kx.����_�Y�	b���cn�4>��(���  L1N����@�F �`k��cd�l���Y�����b/Q|e�
��i��^�0���^#�]v����W�q�:�.3Ҡ#Mu���.�R�|�p_E��Rn�E{? �,�/�Z"��5�a�G�X��fԻ�k��|Wu�	��`|,m��60SP걿����<׬)��L��XF�y���|_��Y[S������HK�����56#� �5Flq
���M�b��7$�`�d�!��s�us�Ғ��׆~���ޔ��X��iSϥWGmY�^���-�|ec�gVdͪ���Nzt
r~�9���f�Kζ�m�w8�M�e�P�V���7�"��zP{��9sA%�u�A
͒h^e9b���R����2߸,!��{��k�90$Hכx
�i-�
�&`U&f2xҶ���{֏��J���9���s�GHj�u555�E���[����0ڋe����憊�1QN6/�I�V��x�w �wof��Z���:�'����D&Q��w��0"�N���L���es�垸�b��8��CNJ��2%'x4���.�w�g����[��5�F�9��Х
s�șe�/
�o�AXN ,R��Q�D�\�%�6t�p g�M�zˍ>���v�494쮔��$a���'�xg]����L�A�7)�T�O�+#�۲�4�2wo�A��s���
 }�浗�4=�$;�v���;%��R��/���Q�*��s��"ߛ6��EZ�dQ9m�[����QC��(=e�K�EU~1�N'�!�2�K�bݙ���x���א���{'(,�ǳ��X��)��ܕf~}�ǐ�^C��tR@�����/��*D2%�~��B˫�F���4��i�nBj�m�����B��Z����(�?K��Z"�?>�nA�!����KO�R�ױ�Q*�)�pp٭�D��bCw�^�\Мv1�T�TK^�9+ !V����j�_�.�z~�Ɏ�5�~��h��_-F�l�(�@�p:OӨ��3�
�搢c��m�5[�Y+�]��gdS�wZ�X=ƨ%Ғ����O##�m���{�#O�L�%x��R��Q��=����~�*K�x�qF����ǉ<�#ZJ��_Gʠ��p�u�����.뫵�%��0�\!�;�����_�N\%�?�x���賦ڽ�7M�H��o}��.��[�42�5�|�����Val�T�yqLl /+�1��@�ѩy�������&���� �1�^�^�'X¢ A��/ѝ�|�
'E5[���N<��n�$���׍�-���(e�S³���T���Rt]7A�����L�Zh{�9m��F��΃����g=��4i9Gڒ�:t�l�>� (,|�\�~ܻ��Q(j�9��R/���WRF����B�N�ֹ1V�%�?�]��!N��dw�<!��*��1�2S�|�l�)~*�#�br�(����f���|l��b�����'ׁ%����V2��ڈ"�,ˊ�P	E�:�u��m����߯�v.",j�??�\���C �{��<�ws�U=7�3�7ȥ��(��DKR�UIZLn�i�O�ޢ�9�|�"g<ɱ��YyB�����^`T���, �������_s�a�����'�>X���Pt���N���Κ�� �Uo�h����.�EI��LiD�pMI���Rv��CVR �S�� ף��A���
�*_'v�����u\���v"�,��FB�����J<�)Ywϋ1J���i�:��Etg����d^��T�v�<Q�&�ˢu*��Ù�|��?{�������eH��P��w��b�@���:ﾅg},A:�C (����D�Iy���y��gZ��:w�ͰK��q�`E����q5
��X�$�a�/�/c�~�m�ܨ>��"tZ.3Ϩ~�j��U9����f��凯�y�q"n')�����e_�f�m�����ĸ������Z�ܿN3��Hּq�υ�-�����fÙ%5�"����A]Cg��[�ؤ�Q�M�P��l[G��P&	X�A��C`J£CѤ<�	�h�C� ̨0=NQy�����0��X�G��Mݎ���	�0��������f{i �G@
k��ny�C��?�ͪӊ�aڏ���g�W\&Pr�qc<y/�%s�����e�����n!e�kY)yG_��9�B8<��\G_�i��E��Q����I��	�L���t[i��"������M��؝2?�ChL�Ǎ)F�D�S�!.�t�*n�ȻE�-��^P�6�[�s�����"�og�!3R+׊-��Y���%�7`�MM�y'�gN
���#�Z�d/��L�E��݋�a)<�t!�O;eʑ�X|�d�vd x�i���1A�2MOBB�P�7�i��l��֡V���.��8��`�i���i-.O�^ն���7�S����8����� �?(�5�Jo�&ȿԿ�Ӂǎ� u���d}�f}3�p�+��7���^|E��5J;F:b6:�E"�|����Orӯ.{O{�������|��`:A*S�\��`	� �n���$���"0?�:�<�W	�n�Bh��x��x]� P�B�\�5~��u�:�"@�p����|������.�2�R��朔�Ey{`��M-���>��bJ����N=���eݘ��&��M��qZ��u�����1v�<�1�#�Z�.�o���ndA���:�"�>�%D���s2�J��8N���T�X�Q�/Fm#q$��<0��c��۞��,7KtA���ݭ�@��S�y�	x�&�,�3��5S�?G����:P��A&KYs~3 O�} �@K��+J��$�/��#���!a6�]%cAU����L�(�-9�Ѷ�TQ\��n�����?�QXS��W���I�Z�I�*��B��ɡP���p�ɻ��l 2R	 �BgAH�\f?w�����S�[�t��x��@Ӿ�h�{�������_�̂`U�T�H��/C��ƌ',հ�<tPZ�5>��O	Ճ�����_O[(s�q�\��*��y�7���v���|7� Ȟ��v5wf��mu���
)��_���Bѡ>��?�+���^3�g�
;�M��?6Ty��8��A�`~F����y,]X�h	HY����Q��d�k�\��m^�خן�������2ix{O�k�}�XB��f\*�8U.Fe��'�@�ETog���n�M���&G����8��ذ���ףz^��aC��ʛ
�p��Fk�j�Jp'�-הx���P�&8�����y����w�7��F}�8��8~I�v��/*X�U\���U��k˝x���ܦX̉����4 ����S��k��b�2�|���.m��ؔ�6�L�>��9Q@(A��ѶL��SJ��jQ�	�᱉R�,�n�)��1(�������Tr��M\}�qdc�t��|��(�x<����<[�C���hlo9[[f;}@:+�燒�X'K-a��d\��l9��4�I�	�凨���i�VR7���Sf4/�7�15Y��1%�G�_=3�a��xN2>q�<�ê�w�տ,*�1so�u�0�w�y9Q�q�����z��k��3ׂcE�E�Єl
�"*�̍�V?��Yn_7�y�C���A��B*H���v�CMD�	��&�W5݀����~��x�it��B�?��/������]>�����6��i۸Q%$���H��u�����;�����Nn���F��p���DEʦ�h�u�X�O��Gŷ���H�w�T����sSh��*%��f^�g+�2&� ]�AS�)�� �j��0���P@���w��-Աs��b��+q�O�c�o�h�U�,��.Jv����ܜ_��s�0�d�ZM-��LbτZà��BiX���j�+�D�1��`:��}��m*D�5H"�M�N���z%��,�����I�� �I`G(ASi��f���^���\��Ql�>崷;L_��7b|�3��b�"Z92:v���;�����i��Y��a0x���Kj�cS	%��?t{0͐�I~��'Y����D�����:D��Ţ� ќ�Зб�N<�?_�b
 !?I��_��2֗1��6}�v�W�1��Y(��a�I��/���\�@�LpPu^��#U��}8���L.�˻�Ö�>�?YQ�ks����:2��=�S����HN���t���0GK�	����E�NZ��݂���N��~؅�%c[���W<y#�t4�D�h9a��*��$���k�q��[���K��������������j!�+,y��3��箾s������c����|}����q����90@�!�Nut��3Λ���\�V�m1qH.�B��c9�C�%��̀�!RiQPWw [�%j|>����'/�����36�����]K�(��,VXg@���E��&��!�޿$E�X:�Q�噝����F�Pj,�P8���d1!���N��6�R$�h�@� ��t�L��P��y�9���2V���s�X{j��;��z)bImDQS�1=̋��h�ZO�n�qPT}�P�fkW$���g�8��Q�(Z
���J�>A�9)�g%d�&A!��HA��n�O�0�Y�l�����`z���֐��v(*s�.�������Lfan<ߺ4h�h8��5�]RXx�h��a8bFٷ�'8��z�h��>*�2U0@�"1�����o�@��������I �R4��t�ugmo�DO1���TA^Pk��K��K#�d���r?���Pg�/�wUT�%YsR��n���_gQ�H�����K����W4P��|H��M�EqO��փp��,��'����a�)��L�LCm0K��Ű���e�&fq��ż����21�>�S^-م��c�p[q��)��J�������L�^bf��@
2.�b�$`�.:������<�T"[�]��qQ(�:
k7��͛�.?���������#_��GXY*y�S��&��?W�5uE�d:p3�)`�5��i��o�7�^���������s��s��[��Pj�w*� _���qz�,ߙ60W�C%�g�Ҭ�e�I�m�MQm���I�C��Wr�}ne�>a�o��*j�cW��`�f4�9�����U��^\�a}}]�����K�ܝ� �@�Q"�Z�����{���y.�����?��Dp��D3{��j�/��ȁ,
jR��ԧC*O�V��E����ư>�(���*��)�UG���`w7����v��}�}���

R@�|�:�c�p��~ӈ�J?�n?����3�6��'_3�ǯ���eG�J�K�?�?�Ⱦ�G&�dT�v)�Ǫ��f�X�Z﬽J��۱a=�\}⩚�W�������)�?{�n�H��oA�JOcr�tv�b�����q�vgO3���#S�}s��i�n;ѵ�<8e������"�Zt�}�������5$-�8�k])s��Vl�����+�"\��f7ez4�H��YC�[�ԏ)�e���2d��sdh�#�`���Z��%����(v����T5*��s�v��j�7����J2��������_DF� ���9Gt�n��N"��P��D���;?�s#m�7lI� ��$y�<SVF�Q;���f�r[�1�е?kv#N�RcB�~Zrʛ�������R�@:�W3"1!&�_��3�Z
p�&p5��_��빥|��x�ǎ��#)�� �ߢ�*+����*u�j�q�� qP+r���JA��?Z���I�<�������x��}�Ţ����Pv��?�?BR��<F�$g�K�@�Æ�΍J�b�]���^��A�L�Q���vl��*q��Ɔ��d*�������g���x ���4\
s8��eJؤb�D@$��_��'� �H����o9/D��� ��-�4�X���A����k-i)�$����� �2t�3Ux���,'r�[+���n��[���j�8�A-��|Gi �\k��i�bp3@V�t�8v�s��g5��H> ��Yd���8�H��gG�A:���(�5_*4���qk�e�|GGq����.���c�ڗ̗�U&�i*`�����Wf�4ߏr�b�β#���	O,R��T�0nōï7>���%�}�C:x�d�|9�2��q__�O�
,��j�����U1Ȭcdp�m>f����bR/W��#��Ɣ�g��F�= ���e�4�׋��f��g('`"l����F|�\T���C���`K��҆Ԇ�ׯν
�t ���| >����
�^��2���mT��D� ���D ��j��Ь�u��#~�u�}U�y�GΡ[�(jE}��䘇����K�*�}T�i̓zT �3DT*Ǝ�c��p�-@�'�?��S�Ŀ��B�`	���/aV���㵯��l=%�a{�.��`گܟQ-�_o�L�8%m#p�E�X��4�;����\
s!�Qz��&%���ڠ���_�6�&�������ffKW��|�W�>G���oRh_�b���SeF�3o������!T$̚yxsꅰ/��X��<�I�d�ؖ��8>>�ڑA*���<�x���Ё���
�up�g �����7C���vf��a�)R��zy����6G�/��H��e���s_T'�O�si"ʚR�_�O�#PT1�r��CP�C�'���D��\�{��w�s`�=&�S�<��	m����p�na�<:^�a��{�Y.((׮���
m8��R"�R�B5_ɬw��}(H(Oh�쓟a�׸o�X�5�(� ���A��\����/( �(]v�r���?:Y(�=�0ӗ8�}9dͦ8U�HeM{���U=�����AFFAm�,�l4�Gk����1���Rz�Y�J�#�����d�`j�/����G��#���Y���z!�Ւesk'�����H�7��`:0�1v�{�Qm�q�4�`6X݅���37s�),0a[mK�bC�O���|��w��}0��<i4ř:�+�K�i�>
����I�w8T�;f�N E�A��87�M�2N҄���[��*k��<�V���ٟf���DkJ�}oT���F�����!Ƽҩo� ބ�.�[�D�J؍�ޥ���" fe��*hť	鷦>4���H}�����_�qCy�щQ}�;֐���b9�I%��٥?%��"~/'�%�����:��h9q�R�]h�`�K����L�	��$O���}
K��b�����[ͩ�Ա��^����O�8-N����w�QZ�b�/�DNϵa�g�zv����6�JH�?zK�-7��O��;���=E~��@^��K�%�6�<��Y��)���v?E�##u��;�xXA�l�_����n;�)*ІI�j��n\�㉙����₉J:8��������p;�j5�ǩѰFpG�q9��?"	���)�+%a�<��vG#���&h��������|�vH@�-�/ܤ�؇�bBȇ[�e��Ϟ���c��8�:��-�'��a�o� |��.z�w��t�}�N��K(�zIkAi;_�N��� ����5�y�ѧ�ՁsV�`����.��	��X�~Ұ��������iW��SD��)��N��Z���>���u���@X��>f<@f{�a��dQT�냬�1�:#iR��-աw(� �4��9z�� ������[�s�F:�0_R�l%N%���X�&T��!�a-�:o _����$f���ה���4�Bݖu��ʩ#��EoÕ]{�����3w�`0�H�!7jSdx5uo�36I����"��o��Y���s*;��|^~�(U�]jg��]q��jJ�5 \G�߉_��='d�ǐ����������Iьp �+%̿x3�h_���P����y�b_�ls,��C�{�T�
�t�kg���B!�ߝ/$��d�.?��!�ڐt��E澑�V�$����þ��m W�;r�+0.�z�ŵ�ife1�P��K���D����xP�yQ�E���+Eܴ���]�ZuxQe���da�z�;�n��L$��t��c��$[H�)v�z7µ�:@Y!�~��|<�t�?
�_>�uH�,I3Ãe��:;�^T��jl@�Bn�@��"�^��:^��[�,W��Z�$\+�|N��L1t#m�|p���d����T((�e~ˌ�ss��Fg�腶Z͛y^}��YL�!��E��k%��˅����g�(�Z�W�j-�|���)	_�B�i������ �,�8�F���<���G?��2��e��Z>2���x�]cf~b9�7�
)S���7�D�Nk��o��0�����isH�ߪ��n|��q�m�S��i��wߩ����x�����{�1[���;c��0�c8��5x=�2f#�fQ۰����l+��> ��1�,`6�U���r��:Mkp�����K�����c%g�9��je�Yv�_Q�"�f�<�Ji\5*�&�Kc��+	&4�ں�)�qd�f�!tSK�6��$�?q�^��aֳe��d� �}���#�>���
R��4%N����W�I�l]j+��Z���K��._O�KV}	{�'����VBk#.��rϙ+2�{�P�GПq��g,�V<��?dSRT��ڣ&|S�{�9 H���u��ml��Q��DL M[A�PE��m��=k=�߈��96��RX���W��(f���u��
\��*�%q�|�;7٨��c;/f۩�; XP1�g�7]���p9%43�7�S(���K��
��D2!knC�bH�C^�V�3���#[I�[bW9Chj�H�f��
�>E�*�#B�K����T��m�U�N'O4��Ɣy��֨��M8�c��De�2͌h8Tt�1���Oᄘ���ҙ�� �)���N�`�.��8;�h`h˩ș��V8�$*��ނH�h�{�_��#&IZ��Z�I���$��"R~�]�H��S�0FƼ�X;�	�&a��hn�G*d��Mr+&�C'Ɯ��oB�ت!)!(���H�~��K)C���砐ś�V�[��ه%U�y���������uv'��x��4����l�o��ٲ�.���c�)0��	>9K �D�{����u_��U4��Ts�uG� �S����:sb�� ��DLq�>uȺ�Oٌ���Ixv��^��{Bu��#d~"�1F6�@ >�Gj�'=	�Bl�4��I���ڵy;��e(v�� sWQ� M}��i���S�?9�;����ų�bA����q��;�%+��r{ǔL�5���H�Ǔ�'��Hzݐ��A��m@��5~S[��ڤ�j=\�:�:�n�mV�(�������c��]���Ȱ�]�|/v�� ����/&w�y#l��W(គ(C����W?_��c��ka5��L��T�#7�9^K����.�X�)k�ik��e���L�B�Лo��p�N$�N#�1$�Z���b��F�H���Q�,�١ ��f�x���r%H*YI��B ,[��0Q+�7H�����Z�w�D2�?����hg��_�DO�<a�>ɭ5�!ݶ�sv]ܷ����>my"�V���8��D�_@��x-:�+	��b�5���,�2Qo��Odʹ�S��;�������߉�16�G ��^�}o�Ꜫ���ȧbp����x��^����x� �r���A�����4V6�}�9	���K���^֮<��Ǡ�-�o�����(EF~#V2ȪC C#^���͵��Ϛ��}������{�`�H��jW�
+���c�N�ީ�,_*�ˌ�ja�Ȉ`EOzR!�ʄ�r�*�/��M�k�|.�M=�o8)��2��^��s ��+��8���,+����j�ی�+p�?�/Ǽ�;o-`Z������._��S֮$���j�d&�8��\6�2@���rZ����ͭZq��@�S����[d�腮ʞ6E�.(��M�:9G�H������K���z?���7��!ݸ�Q�DG��L�+4�']�)�+��`Y��ベ����b��^��/�e���cR)|7���``[�34+ϧc��5��E>4���;)e@�f
u��^�V��T�ؠ���%z:���p+�Wgkv��׸��6y�g��D�t�w�s7*D;�GK�s�=o�>�:P>-�5J��H����qM��>D!�%Em�G�@�Zѻ�/T�6�$zM�<N9U��ا���qY�����ں�$�6�N��"��x@��� �>���zzH�銤A�`��Gc�T���]���:qwԋ�����]$���y'�~^�͢�Q�k>F��Э�LH����M&OJʱ�<��vU�FiFo=�o�(O^ւl�^gԕ�G��a�l���%aK�te&H�}w��%��~}�N/;'�l蒨-ʥ�FMA���GeLOϱ���@��|���+�s��=���x�Xѻ\���c�Z^I@�=�F�Fd�v`������K�ߖ��ݏ͈���F��9�X&��Ā�$�(��t&JJ��p�@
��ڔ�Nrt�^�Tq���"h7�ƪG������;\78U7,�Q�%`���1��J-�k�?{{�>Ͳ���������1L�T���|]2����W!$ˎ�9t�-�Q���e�/�Z�UnA"W�չ��$�(�~Fr�T*I�W�g��Z��c��T'@O�����u���֤�-"��zK�Mq��ۄ�N�3Q�Q��3c�$�kLfn�Z�]tŏ�u{�5�9.�/�b)��*�æz���J�iSZa^�]n��pv{��)��������������e{+6��6^z=��/��$��QH���/u�{�|�\T� ȝ��~+�6p[F���5��pԶ���[euf��U�b-a-��Wbw��mE�*����I:�5�I�
D�mK�0���R�_�ϯ�2�M��ɒ�u/jf�}�H�Fc�s����+jg����j0hŴ*��v�n���\;���Vy($]M���~�x�c���F�τ���]��h {��\y�m^�W>PKTBn����a&�i�B��lT�[���|rջ455oT��ݧ׻�rփ��7�-K�
�~�Y�6SK��_/���,+�<d'��HI�K�`�Mo�5��Z8^�&6~������("�"��0lbMLί�i/Fr'���#"R$w%�7�m�4��nl��]��Uk����1��4ҶS��0t�ͷ���Ǫܺ2,�O�k���\d���TT�r��!�c}�&�Ƿ[y�bF}=E(h���&9Y�d��S��~z�ѾqE���k"���Ѯ��I\�G�л��ԖIЈ�0(@a���GT��()��$צzܟw����J�U�Q���7tef�b���R��<����~���F��s��^�������M^J��au�r��mj�'X�@��ҙ	6�����滆y��6b6�W�����?�����B��r~�qP�H�x�ţ��^b1q�U����Ҡ�^F��n�n��7�5���(�Hɵ���Ml����^��;Bf�%�ɘ��4)��T�'�Ŝ�`��F�Z��A�{R�9|P���
���?���K�q�3%e�!P�������U�h'A�YU�Mf�F�D�� ����,���	^f��P��-��5����t��Mb�P�Y(쭾�3�,���`�,q����n��&�a�E����F�6	���ǯC�u�E��� �R������2��Q�o��9*��Gg��Zf��M����f�3��T�)x).Yȅ_?uN�>>?j��vOb�GAk��n��W��%!���?�K$] �j�eۘ�Z6"���ĺ����#ʤg����Ⱦ����qh�i�C��%����뜊�P0�iG��B�{�Y�dщ���-B�lN>�Py�������{�����Q=�ů:!*h�1��A�K�ճ�P�zǃ~h����#@���`b�X����D�^]�hE�8����G�P�P�i�%����5N,����m;������l�����d���HX`�<����n	[�όE%��R;`-��{�xFX��M_"X_�����Q��}�@n-4��Bo��H����^�e7?�]Q10��|�$�	 "�Զ=L��T<$+�4z�O�=?���V�/����*�H�]�m@��Љ�I��D��c��e���&Xeg��Фa]6֤��rU;�@��^'FPj���dl�[��;e�n�=a�GP��W�{f�$��~��t-�v�.DH��o�DNj�૛��2yɘ�X��主��V,�2DG�,�>���m;���#���h'H����丆���� e)lM�R�Ai��"�N��~�g�:0\<����F�;��P��4X��:�JFʕ�k����X�˅įܐ�)�<!�����%|�JT#l(�4V�}Pf�Y0�؏c�2-̿�ج�r9�+h�â5s�hm�����U�)"0�2lnESܙ[ݕ3�JP�G%��B �z�֫;�Ƥ#Ƞѿ����MT6�:;�	�]��:i��@qH&y%D�ɢ��TPg�*Q6�eZIm��(}�pI�D� j^�d@�S���>T!O�Xb'锌�� `R�@_A���L��8`
a=b!�i��c���n���q��5'OF��z�|�3�~�ͯ4�˜*�ix`�6�n���l���0cK�;��蹿��o�������r��q����(���@��-��zS W�_��3֋غ�Zi���)k;��
��b�T�.|��rz¦���L�zs�a\���|��?:¥9�C��t:Z~���qY)g�?n۹B�3�)_��DU��������"ҕ�l� �@E�U>��+O�S[���ޞW7k����KĔ �/Y�=c;���f��Rō��g�	�� ��-� ��O��ѯ��r���4b���?��|�Q$�R�Y�Sy���
��vk�%���+��p��k�K_jH;R�A#�x�E�0@�CX/j:���P?7�믬�创�z����Cxh�N�­�J�Wd7=G�)|~ĚL���b�"))�8?�����x+t�S��:��Y78m�r?=jKsme�q�39��Xa���-��-��1��%����:PW���Z}A��[���:;�~�bx� X�R�G�{ɂ�Hls�{��܊\�A�*���W��R�eAR�2"��Sq���:��UT�*��9��O}N����}(�R)�Q�n
�p���3���uǦ��6.�RŉBjFe��U>]�EK��4���*QN5�ko?��7�&��=Re�X5zD�A����N�^�˕B#Q���тFm��`^�G8xE�{Y�n̬�z��O��
9d���^b��Q5$)9&���c�'�!��=�[�K����v=��}J�#~*f �#�B�b
���v�v�OW�9x����j�6	��
#j�DU��f�$��T�X�KR2�*�����yCO:3[� �u���`qT�pe@�Ɓ	�O�(M�H�k+/�3�V$�uD7TU�����}�`5�⒒XU"%�Qp{L���Ia��s�L�X�$63��0���Ի���Us{h�?b!+�)�2k��ʋP���2B�+�ո\<�C���9�l�����@}�h[���S�Y'}P�n���8�W]��v
��Ǆc�A�d�ȩO��f�;RS��?�Qc�� ,ի��'�	��r���@\��e�H�.��Ѕ��>>�2�Z�H��mtG�e���e�p�C,݁3�Z��)�(��Jm6���ǩ�7`ju�������Ok@C�ث�Ξ?���P�y ����X3JwѲ�u�ʹ��̖�ؼ��[�4
�5������'�;$�WC��eH�]�Q$	�%��&ym�'�����8�v���Mw�>����=��@��h'�Ȍ'��)�����͍]3�� �-���1�<���B���?G�7cHl�K�G�M�����df��%�s#*:����D��0Ev���W ���7��%4V���/�26��=H�� >2�7��0��B_+t��=����N4�'Ђ�&�aó���MQD�l�����p�hOm�%�&�Þ�3�HЦ�R����ei�ImI�qJ���9;3һ���E����0)N�bw4/83f,�e�j%k���Dg����{f��q���g<puiX�a��x�3S������3n��.u&�>�Zz�W'5.��m[5`ؑŻ���"ë8@���ʲ���856��&��.�ݾiӪ��Q�/~�`:�7U&��c��ֵ�Y|K��Sd��
��f��j��e�:���}���x@K�PC�����c(�^�E>�3�.�n��#h��#��s$|�!��ҳu�B�S��B�S��!�h�j�w�Bo���g�C��{	�(ZB�'LƜ� ���K��ޜ:�Ўu 3SX-E��t�a��{Ϣz*"�ޗ2mSAk��=�/��P��.(�| 3�ET'����(�ؾ+�����6���-��{��I����5�ܘE����yy>_o���Fp��������WS(�F$��ځ��?�d�n�@jݪ���B=�~BY`���zs.�׻zP�uV�:����،�%��q�W�ؠ{U��FC������O%0�M=ʥ|ObM#<$g*j[�B�:���ݴ��!zHڛ�U��/>
/׶�x�9������\=M���c�:��S��w�-tw|���C��\e���| X�	x�b�p��>��&Z�luZ����w[���:aC�f���	�U����B�AO��՟$imZ�u�ƣ���Y���.4�= �*�E��q2�j��&y��S֩��,�E�����n�cw,�qe�������>�I�R�[�V�bB2�� ��E�x�#��������ÆB�����B�
'Q�J���UU��ڹV�C'�:~�H#�Su�״�&BŞ�MU|�����`�
��A���f�¡��+Jd:���J��ؔ��"��1��c
�20}�+�����%�;�97S��<��������3�L�_�h��ٔ�uM��UÜ����5�d�d�a$�s{d)�l5�j�c�[�x�����g�N��!,-PD�f撟`\��%Bm#�c�Ҧ�R��_e�R&�G.y��L4�8N�pj�hJ6/�:��lCf�����I*���<y"�d�&���ħU�q�嫉`��ۅ֢%qi��{�G��K
����ۀ`��f�1�ZT���n�ǅ��,\M���i��;�[9�[��a�D}�� T���B�`>s5�o[�|)^�Y�Ǉ��g�o�+�
t�[��&ݽ^�j5�b��-��̴Iq�1�����Ʈ~��^����{����[k�[!� zo����<�D��}<���Ֆ�Mt0�J�)N<Mi�e����a��i�@T��h< I��2�h��;���E4@���΢�v��x��`�O��;V1��7��*n��2�^�꥽�v��HS�V�Ð���[��EG��.x��1��:PI�d�T]�w6����uj��\�<}��i&dY��M�x��(����Q%y^����K�P��u�c�K�YU/�A�ᧈ��2d����KS?��Q�Zi�/�R8,F_�i�g�=�JQ8|Ζ6����sL����E�[pk�=�������M.2����2	��m�0��`/C�uʯ�����4�?&���!���(1��,��E�%kS���'5��g�j��B%�&O,��90���rG��}2hg�R���ؿ��9V� ���Ξk�O��;?�g�j��x��hKf�n���D�q���ܳ�SԺ�������~�s'6��5����?�{�=�'	��i��b1؋<*�ۊm�:�`67_0�;;ǯ��rzv��w~7�ł�lT~ d�B�.��-���K�b���L
z�Q���8_<�l�Ǡ�iN���]��ɼ�#G��>-H�0�"L�M0`�q���d{��Z4SW��Z@=�M�}y�J�r<"�C� 0b�7iܖ@XI�*0��� 8��Ӗl��g��y6˭<%�SB���q�2Db���$B�%��4,.�����h`�/�K�#�0�n��3�;�ZQ�pB���ϵ%Jy�<㈨o��&O���������,7�s�ͅ+�a����Z4E{7�i���a�y�'���M���ٵ�)u��|6�?��J�\��ls�>f���e�4|3{M`-�0���\�;H��f#�O�	�1Nz����*xTI4lGV�_{���]�A�* �������l;���i��Xp=�#�y�Ȇ��6�	��s1z�n|�m��@W�����n.��[�Xㅤ��Bʳ��G�3c8B�EI(�P?ud��t ���'�ծ��v���Ʒ�p��E���4�=t��N�Z��n/�Ѩ� �r˾(���4��W_p�
�{%�@�T\R���6i��'P��樌��`�+��;�� �g�$rW�۵��(*�/��h0s(b�����Z��HR�BP~�5#��!�=��VE���ʿ��	 �rW1eR��?G�]�!W$d�01�[��'�nE�i��z��!�Z��qZfY+s��M
p+On��Ss�WMq��*��҅H���'��1�����y���𢽧�sԤ�
p2��A���M�Xk�B�n�R�
<�����y[�i5a���1U���Y񐷇AEI{I3��� �Xo��wB��ashrOol"��[�ηǟ���-]�K��Bb���&Ю��k�Ŀ���?�}��1-�%�3�����m��_��;�#&=�ۋ�w�#Z�)2NWf3��]pڵ8�Vh	gd�¦M�s�GE����?��F�nu�Y�+�Y-ʢ{��;���u��4�(\������4C��������-��،��W^̇��ز5���&��R#޸����h�J�|������e�FJh�0�z�( �5v��#Q:�z=mB��[\,�IH�If�3e���:'�{oa�O�<�u�δ���A(��"d���fn�qV�2O#
yp}�j����_1����a̗�K]�![�o\����@DЬc��S��`�E=3����Լ��WO��j�����QM,0������B�����Mw����8e��(�%���Qɜ�� � �n�L*����k����]f{�HJ;;*��%I� �Q���)��עhz�ʾ�b��]���%�k}K/^E�	`9�]~e?�٩%����Z�`$5�Y[-vu�.�z�F��"�mIY��n�t��6�!�<��vP�48Y1u���q^����+�u�5��:f4�qC}��TS��w[�9��<��U���͌�lr�y����5��V�N�Nf�eXn��QM�i�e�"
����UQ3	S�Qx��K#���T��0�b�3��9;?,�-o(�s���iA�F.�9�����#~�l;f
�	�;�K��-s�|�G��t5H����a,oO6�M�FO��q�;�Rm�TP�r9�b��Lҫ��A9%ݪ������bW�X�}�����º�+!j�k���D�C��:=kwuA�����$+-���pG�Ŕ�ݧ�NfV]���=j�֓*��T�4R��Z��H��L���2�S��˚����|��>/F��U-]�(��(�+�&�dJ\�^�תw啵T��e:z	*D���6HFO��l�����)nd��U���TwgI{�^�i��f�����"cY��h<�[7�D���.��<?U����֞�ʸ-Z�|-�qe ��]��sS�<�s.u���v��Oi�;�-�H�jiAo��p'��Π�QP.���"�A�>��-KW���R�[�� ʄ�um���Sg+��0���z�����;��Y�	U��s����a�����+���Wn0O�i`�.�<�W��ZI��d�I�ls�1������?a�<���
_me� U��o�9z�naK�f�p���8���sa�L�cC"��*���l����JV
�}T[xp�F��˓{�tՂꄵ�/�K����<R���+�	)GWҭ�IX�m��m!����o�0�W��ܿ����gQ�S-��W�H��T�^A�y�-CF+5�Op�����k`r�4�T��,B�zm�P=�TW@ ]�V�ty?���w?�.�_�,gvbA_�p�A42����	P����eih�ژ��u@�.�K�wޭb󅹔U�4��@*�%�}YA�Cr�����,��%�Y)\-��KĢԘ��'�4熥Ĥ#a��4�m�2�JLX� 3��}��oH<���6H��vM�.�"�R����T�(�(T��Fg��y%��A7����x��D
v�pYu���D���Q*�e���`�D�{_�f�^p�OK�:m�t�[�Fj��	��D�S�����٪�S����B�¥�)(��9�Wr�^w��P���B�[X�9Ӭ�z��_�:���B���J׌rTb���2�
$�����s� \�p�Y_���.�%ͦ= $[� 5OA�=o�+_rn�����@L��i �|'u�zH���D���J<
��� �֣J	&IT_C�5�|E%��3t���BȶZD�VO�ɴ�gq?At�=�����3�8���bA���y��Y������r{"���|&n�c0�A�-�u$��Ŕ#��_���u�2��J�s��^u��}�;�7�����OqyԒ/}����45�(�*�Q �`�%���}��J��o�^��\�0~���j*@�>d��:%p�l*�bTR��cL:�WZ��Hk�a���vt}��B$��{�r�7��t
�x�4���cbG�U%�,t׉E)��uD�v�ܗ;be�N�$�S]/��_pag� �	Z�Ǖ�*�ٱ��a.�g=N�F��bw}}�G ~6I�>3Z���";�9�Q0{)h��C�U��waGL�%'�"R�V��.<�2OM�2��ʔ1�ڪ������'�P�oHb�Yh����O!�W�\�\�>�OnI(<f�F8��՘S�ߦ�E{�S��J5��4���W�Q��<����tܒPJ9�2v�C�ABM2������մ˫1���%\�;�
�&�V�':�?e��V;\�m%����4���W�10U�>\��LLwYyi��yQ������Gn�㵤�P׉�y�������Sy�J6��"7T�9���J��<��w���u+oF�W���T ބse�S�}s�o�dW�F��`�NH�u�_�7OEi��q&���;�/I1nX`'ѫ��Fxv0aҽ��e&)-�˦圙�{Ds
�\ϋ�bF���b��Z䁄!@�~ؖx��Y��b@�ZP5�[e�`똥8����5��+�I^MW�<qa�\������*~�{��L�ۣJd@�z/G���1w��}�k�]����d��eɜ�m������7DJ�<3����ǟ���sN�VvJ������1�"��������0�6K��P��_q&��U�=g픪<�1����b�b�	�1vn6�E��ȑw�H����<�m-s � r�F^{[�AB�0�d�Bw��(}����x���^(o)�����C�k7Kƅk�R�
�+;(vHҁd��_4E�]��;��ثB��PQ^
ۯ�z��,�-3�o4E���,u߹���ހ�y�ܜ<4@U,����<$<����%����*�����^�7�����oƷQxb0��b�ĳ�|(^;�+�]1���!)��l^�����^�K'�ҟ�gLyE{�7y�?C��=əCL���ݡx�Va��ku�kצ�����s���O����y�i~��@8�d~gFQ����E&�ދk�W ��%�As��Z�8J׎�t��UI�>O�T�k��!���J��/���ӵi��o�4�^��P�J�pȽ��J�֦7��%��l�
w �q2��](�P��5;�m=��F�rY�g�P���d}��Ê��OI�E��M�x�I.!i�	$>L<	U�Ukͪ���1�
��!p��x[��d?l{�5+nwRɵ�j($�4�:^�Q-�[�����蹖e�x7�%ZqL)]���ԛ6�=x�+��_jj�QF��c��O&�W�K�	�a��Tt�	�5�=K�Ho��I�U���u�L���렔���r���ֺ�>p��C���K"\c�"�'V>F@�3˨��["ɂ��s�9���� dE�4mZ�(���(_xw^}RMB�v�^��_[���c�(b���r �rg�+�a�2���P�X��u?������k����.�wA&��Q�|Cڮ9��X;���ی:Ŧ�E"$������w F��wu��czE !�-��7y^�Y���
�V��1��|�O�}�ĒO��Y!��t�L��ܯܓ��S��M���������6fB0n)�F~g��ϐW�Y�����[nO¯�@� 
َ2�,��@��ai�,�nN���*F�$�s�Dzk1��z�������h#�f�Njc���y��[��ƽ{���KnH�����3Q�5Z�n���F�*��L�rkk8�ދ1�߁�����b�6�Ґ�2*P�����ށ=�u��
��q|b�{�ӫP?ַA������HJ��峈C��e`W��0e��<�J��)k=�e7�G)�W�)�p$�u^2Dý�EO�N$�n�,R��{�}�C����mv.�8�jj�t>*a����04J��c�5$Urs�8qMϤ���ԵA+o�5�݅'������z�r��m}��OY4��/b�,ā�;uCU�Tp
O�@��
�-Ir�<RBZ[��DVu6Xe��#��$l�i;�Ha��D�I�p�����2��FJ�"c3#����kO����[O�̓C��uI�'0<:�J��G�9*�8G��f�ia`�r���x�f�����w#pԱ��X��d�mxB�ٳ>DL�i��v��#�
��7%�-��&�x��j@԰	��՗ܷ%�N5�  ��Cz��d��<�	.�W¬����~�eT��iv�C4��^ˬ�B�E�3�ݙC��/Մ��j���1�ڰ~'uh�k_b�{�"��������O�rJp�rT��	Q�0J�g�%D�>��=�6��Q�����5�:I�dYQ���=?QX]e:jh[lE��O/�[�ʽ���'(��4�N�k��.?��%�.H�uPI�>�9�\�j��\9��w���KYTl)�[yg1QT�X���jϻ���:�K//C]y������JG�̃p�h�6��S�����Ѩ/ҕ��P��oa ��.�D�|r�2"BsTX6"j�5�����pW]K`�Gp)��\T���m�Y�C����4Մ���Პ�,�V$`��cŤ��m��%� �6����-�`[b ��9�p�x�5�<��,z�w6��y]��sl�9uO�r�� ��l�dq�	7r�Y&���5W{��I�=~�\}�J��$��8�m�0�+4���fOd�+ד���1�w�;�A�h7�ކq�3wqF����ůP����&��==���!��Y�U'7Sީ�y}ZF�%E^}��(�h�Oa�9p�?�p���{���Sü�8���.ӭ���<y�?�xq1��&v��Z5,�	Z)��y�W�
��`;Y��j&���!s�����#ģ�t2	BjQ�8ڑ�aO�F�	���W%�acC��R5����mUC���x�ߞ�&ׄmG���tp���e�����T'?/�Q�С���ӕ��C�2.��,��)�xL�T#qA��Fpp�(�I5�"k��"ׯ{�F�� {
X-A��I�y��Waj���o�ϊ[w��dl��O�"v���b̟,K"�4���(-��?�id�^B}'�H��YF(ʛ�j�/U�to/e�m�m��W�B�__��)gE�*���0I�)��&<�ƌ�`P�Űh�9�w�N�����x|2ŖFSx+�D	ܧ�)�xk�Bo�O��]A�"�9q��G^i�8��z�]��@*][*�����d$O��4�-�n*؃o�=rQ,��t$^>�$/_c�K-�@�٥o��{>�_�����ړ���[��fQ�,�)����z^�2�w��y��g��]>�:��N1yyڝ���Й�"qȏ���|���?�#��:szO��V�*?e�y���Q�~���p���En��%�X���{-rɷ�p��Om.W���� ݄�(#���.�.n,{M;����3�"T����k��U��Ø������XR�Z�?�W�E����7�� �M?���ªc�*�἗~���h�y���q4V#���,}��{�ǹ=�R���O;�.]���̟�mȳa�Iv�"*���9M�Bp��Y��M<q�+�*�N"w?�*��,����$���u-��r�9r��P	�TY1�u?,������E��?�u���Ƞq�`u���f2W���P��]&e�x5�$\D����M��\X@r�naٜ(��I�� �\�Op��D�W�I�m{h�ɄNܺݍ�}���Z�
%�"i����%�(T���,Зƿ�K�Ҳ�M�UE��澟��J[�b��o	��Qp�f�1���s^�0�����"�Io!{1��pS��)kU���=�+���U��i!�������m���6�#��#���,[="�}/���7�b��p�Q��N�����s�VC�kcL-�A7�7�a�2���Z�;���S��!��0F����8fo��Dq��,B>�I%���k��ؖL#T,^4:1}:)W�`�o׃�:�Lx���p O�>�]1yxk�XY#�'�
�f5$X��� 
A�H���v�p��<����<�;2��T�['�*@������f�(��eֆDy�\�֌������%hԺ�@�u��O�QD�xԶ�"�Lܫm�;�0����Y�`͉��ox]r	��`G&�V�o6��?B�����&t`˯;��U�A�����g$�' ���������I�\�E�2u��]k�>���5	�SWo�m��rR}���{�}&������i8��/�{���QI5>�K�ȕ�}��nSB�8K��z`	��ڷ+�d[�d�4�yԄ���&�a@�.������`n&����Z�[����/Hsc]��x(���C�%�1gF�q���8[`*#�).�8º��	��(Rԣ�L>V�6�����'�le@Z��"	9X�O3��q[��;���=c	tj��s�1mfב��:�M�E�.�Z#���c�����IȎS򢬏 �����c�j�c}\�>V�Q��AF0�W�]�cSŃ�:\���v���x�:��^�Ow*HQ��e,��tp�3�������ٰ�6�(L�Oa���g��ݶj�7h���ƽ]j*"��#�PY$KC��g���]l�Z�퓺�nQW$�a��[��gLe�ic�T[�6�Ⱦ�������{������R����D�\Ɠ,�E�����=��nRr�� m+����ym�h��]*9�GPL�u���\T��y��36��&�¹?�ϑ��;��-�ͭ�Z�_�H�~�(����]�0�*��L֫��I��A&6�4s=��L[$y�����DJ���H�l�� IȁA�L���mVQ�D���/�a�
�J9����
ͅ��U���=*"�v���t�HI��	{K���L|P>>����9?��4\/��7�w z%1L����)���6������Y�ם�j�g1����� *�(�6/1�+�ԬJ\�D�R��)y�3wX;&��6�����-�5������0T�l���>��%�w�ȗfVvz�
�ԭ�����P��`4N-�@��w&��S��L��"��J63'�"(�B���%h-�p/(�K����}�*��۟�qw�,���*�j��_$�5Č��i�u��A�r{+d%�\4�b��F<d�6�$�ʵ͙�*	'��qM��q����9 �:n���� Zj0��D6�wTaxU���m��o&J��ꆶ/45��aWo��~�%�D8PYxa�cC�w�Ϻt�ǜ��I����;��U��y��Q��${H�z�k���G�C��h)k �(:Jb��1V�	p`P�e�4;ֶ-1'�8k�ڌ�|B�;zY��	������� ��P)�q*����pmk*���ɄKO��B�f�4C^bz����y&b�5��\^�$E#��d}?vx��}>��O�Kޜ�]K"#(�����a�d7��%�����zA&�y(s}&T����u�d�u8�U�ԧH&oizC�rƗm(��D|����d�q��OH�7�)�d���2�NIU�,`H��H57�z%-lcL�L�0_w$b펎��L�q@8�BHo
��VXO��ԕM��.�k����E��N<����?
(xc�D���w�V41�d��KѨ}4�#�6�'N���Y�t�a,d���uߧ�ɱ��y��ߥc~]�Z�� � �]sy&��k��R"��\�WI��6~�S�r��D��.w��RhV���]�ia� o�B �TD�&&9\F+������^}�,�C���:O�F-�v�dv׹�S,��>3%$���σ�O����v���3q�D"�F��5D�	N�|�j$H>�1�Cx�j��T�H�N+",�~cN�|�\y;� �.�����rѢ������[(��֩j�X���s�L�-��^�4}�}���ʅ<�:4��Y(ɤ�L.iN���3S�|��ëCl�h��l�2i�t9h΃@Y<St��i�ٖ�P�,�+�4�D�����Շ��Cz^%�/�P#|�i$���G����k��uK�R�ڮ�PQ�d�;1@���ˁ\�
y�� ��em g:'��f�ksBmF8�A��Ū��iS��&����P4�L^��������MH�>$�/|�|l�%hNF������*�T���o�Œ�T��醠Q�+��wGM�x#�Y� B�n�ne���j���"`���2Rur�&�8��=��2^7�Qg8��t )h��-ZMR}�r���5P2i@}��g����Q��YI��p�jWg;g�����%@�3�m[5v|"���p�T�ȾH�R/�C!0_KB�W���ٽ�K���!��:��;������p㺊���ۈ����ۛ�ނJ�=^#�*�S,6/��m�����wJu3���1���3�N5�+<���W��ߤ=67w	�[�*�A���ݮ��\#�s�_���J��f��("�RS0��{�-���w�O��}o�'��SW�C�B���6�F�*E_3 �a}R��kX�'�u8��0Ԥ�1��==<��3t�w5d�h3��ܙ]����wJo�v������F�=�gK�C̼�a�zG�A��M��!�!�&Y
,����:<V��O�Cp��g$n��TN��[��wϵP�Hv�F�_F\��Ӷ�z��+��T��1b��>v��O��fNQ�ԯ9"+K�����Rf6`վJ�V�������ԚF���Pp����B��@�fG��O����.I��mJz�FF�
�S�O�(>�2ȱ��Z�K��˹�Kt��|�2�؏�R�z��F��=����Xx��l" ?�F��橽)����g�/d�[����؁�tgrK3G�����0�$Ш��'x�2�'+�mNxƑfD�-��J�\�	vB[�G�|:���=MAQ���8B�.ԓQ$f�#��<�w�Y�4�|���8�ܩ�i
;]>�0`�W��~��'��`�����u3K����6j&�4�<}ߛ��g䙉�ON�"\͓A<4�dc.6:{<�s�B����H�����g+W��,���5S�^�����l�=X����7�M&��b;�ƭ���!��*��J�  6�1�u�%�5�X�^�b]D(8������5CY����L��␄��|O�i��L��UP�3���*�Z!l�}ť_\�� 4�W�!��-�*����Jm�l�U
�w�f�{ɼm`�S&g�#k`�<i����(����*\��I� ��F}�7RX����A�i�~%�(!ē���rf��Y&�����%�V� շ"Yb~ju�-s{aL��~�ץv�!,���D���2�Bwgi���r�w�am���Т�BЪ��r��}�sR)���3��Z��܃%�fj�եM?�0��ڷjY[��+H_K#Ki�hq�]��P�XS״�ۀD��8�`�#}����O+�+�`h'm��aQ��N��+bJXf7�&��kz�!#$D`^��,>s�.�y&�xl��sj�2a�WEV�(���uͺd�QiQ��- �ˆc.)��eC4�Q�\fy�쥫�р�9�7��^E�a��*S�.��B�3�t�����[Sd���u�'���L�{I�
3HD�,q������M�����;�J������ն)�>9p�����סI�	�P(~�bN��r�:te��!B�*��l����-�6�43����
\�G4���ƪq����l�:r=TԔ�C���q�Χ��L�ڪ�].�V�?�]���
����"��*����q�'Mc�ΉV+ԍ�Χ�I�x�K(��<0����h)[�=7���LIUE<�ޗJ
�bL�=�(^�m����0	��P{�x��n���П��ꇵ��CU+ܘ��š��������U�hu����oېs& �v�4X`��C-�æ1Y"�$
�7�q{:�v�얢P1��cF�ŀʐ@�txŠ�d��@�����3kp =\��e�J���7&�&���8-��C�$Y;�v���s渏��ݽyB�<=c�� FQ\I��{f��:��s��@E�s�C��F\Ȝl�+`
օ��H|@��0�/�7��(��̗��ɴ��d~�`H��lQ`�w-��`0����<�' ���;D��\K�'��~��r��cwn/8@���n��)����S�%?�Mo�f�R��r��e��^��2�*"�B��ov��-����D���2������ǈ&��j.��p/K�K(A�w��DO~��-�RU�]d�8o���{� ;d|��/�g�F' ��NL 3^���q�K{؟���l"];������� SvU$������wB�M��=���!,�7�h͏�U�LJ˴q\���pL�=t.��k�ö$�b�}�H�ᮛW��f��>� (f4�!�EމrΠ��Q��#�ZY���ݠ$�u�e���ໟ�u�P�g"��BW�jl��� ��z����(�A;2nIc��b�"C)�߂��Z��*�w�"9�����
=j0w�(�R�Ƒ�P�t���l�:y�6Ai�&�X�E��3����
nl������W�d�v��@Qqz�πX4|M��R��țS�e���`����Ⴁ ���<Z�B�{$����񾟀��������`��ص��b~v�iJ�7g%�ΞL蜕��XX4u3ikm�Q�X�﫱&lF2@W�	L�;2�q@\P���ۧq�j��#�GF�lD���p͆������E1��Qf�F	&e�ϴ^�i_�b{񃿒�d�]n:%��eq�ෝ՗����ز�V��H֔uj���k�>�R�]Z%T�/L��w���X����up�iGv���D$&��A����SO�˳$O��+�r!�gT�h����X��(�k���l7���'rGB%<z�J�
��'�no&���)>"%n�U�h{��j�=x ��fxls�(�ư4��:|�z0�ٮ!��z*��a��03���-��wsD
J�����Jh��2~������B��'kj�	��/��Y\�j�� �E(]�r��`S#�uN�5dz��V�\|�kNڍJ�FW(
��f���R=�*T['��۫�t��.�3�C������`^�����X���=)���8�\0+M���T5���c����B��~␃�P�p5�`b�(�\����N�%��V��| � �DkOHd}��(P{4�
��O�7������kR��]u��y��**�]���f�&�W�]��.{#]� �0�8�Y�묲��LGVY��|�([�����
���:�����R�8�d�״,�
����Ri�PӪkX�n�v��=�H�hޛ9{i��t�
F��ц��C���'(��]��6��tؑ��t��.ܖv���YE��x�`�|*HrA�i,�,�{�I,��NA
�/���X�y��'M�`�0#--��A�Y��@��4�_�����>y|���.������ҽ�fѩ�2����b.��&<@�*���ԃ�~#�sR��o���9/��;N7�W*��K"Y�l�(�!�>Kv?З�S�V�������7PsD�r�!��'�<(_w�����4$��\���6_X�'�?;���w��Zn�e��)����Px6*M���G�K9��k�O:��<W
}!���~�{��n�[�V�j�ݒ�o�S~��@��k�JĜ\��5 G�;�o"V�rl��c��U���u������hr0Tw��9�x�h&E�k0�����#����$[h�w$��ƶ��j��X?���԰�5g����\g���t�+��E�>Cu�Z� ֬� nM�z�Q��&��ǲsf���X<����DՏ��Y�]5��$�����_1�h�긁?Ɂ��c��D��m����H�N��� A@rYS)b�y�����k��5���@)�Ra��������i��E镖��QxӇ�jgt�tXEç�M�N?�k�+X	'J��nY��N�4���,��w�Po�����7�7�b�rJ��]s���
Z3-Ve-�B��o6c�Y�Wa��*qV?$��� 	���1dB;��C2���.%�8��# ��J�aq�f�[n���1�T%� �)��fą�`�˨���ǟt����?�=�(X��d���EiK��X�U�i��,UQ,�Юy̯�ޜˎ��'&SX|Ib!��9��u���ϳX �ߦm㼙��d�~�T�T�v	s��@b���8�=.0�W���:^a�[�!P!-�z��hc;�	���|ֺG=E�G�-7K&��aHp�(J'ĉD�r��
%&����	��EMJ��C����m��)b�RTx�V<�������V*f)��������
3�����F���P�>-�Gݗo���m��$�d�f���!c~z���#�)l����c1_��7)�����JlCK�Tȅ���W����^�\��������=�ϊ~���%��[j����oH�!��e%��Y�l���E�BNyYJ�NP�y�l}N�|w(ϔR����&Gk�Md�P/1��s�F���/��YvĊ���O����P6U%$���p��|=�$���2@�b�02��@����~k*��팊�T�]Ǡ�]&�!�Kg�Q���?��&w�W�zX��J��\���D\�����=�!�R�a+�P�����h2"K�Oa`Y�a�
G�*{��+��⠞s�����~q���$�>�]��:���ɯ�E�<�fϤ���!�@c�D+H�i�p�:}ï�)�Un�N	�=��	�lC��M�bEa����iA5�{Hc�K6��6��Kzyh3�)7����ޑ@�ӱ�fy*s�JO"�05��]}�Qsa)5Jpr}��pGV٢̢�1��*�l%�#�A8�v-0U����� \[�yҎ8��SD�SF�F�C��"ɭ�U�?�,1���:�6WG�^��SD�tR�&.ͬ�_���m�ކ� s���K�p��9�[�[��Ӻ�, ��u��c_�@$1P����>Z=�%��q�GP�gݾ\�d"��Ĥ ����nY��_��MA5���|�a�*I/��ܘ����������� �P�t�@
��Kīh�伻�tJK�Ry߇\~���O��c��V#�i����~� �n�iR�R[І�O��5a�{�!�a�_=��?ʑJ����h���*��`�eڐ�+K&�߱٬��p��$	7�������:�J��$=��a���W9p3z�0/��c:���Wh�� �k�o|�_���&rBj.��d���nU�/���J�?S��h�������r��QC�+Z����y���[=PX���R�lӅ��\(xa��i����T��z��(��Ѭ+G>�)-lf@���4f�mEC�t��bM)e�HSR1����&}s}���}|]'�>�y����%��-��{��Y0L
v�؀֤�J�цlk�>Mp�_�X��a�n�7խ�ݐ��+L	��b��Km��X$'�O{���Z��*?�oKt��*=��zH�8tw������z����j8�LFj �#��X����XّW���t>����ͥ%��>�׸5����6�Ɇ߶����0M{(��I�;��|釾\ث��Kc4���*"�gL�S-���+�g*����0*�ed3���ƭ>��$N�m���ˤ	5vDŭ�W2>:�b�2�Ҹ=R��"Y#��W�:�H�<`3k������D�"l�Zq�OK�ϥ	/��BE��U3�A�7���l0H�-�7���#�I�\�=˲����;�i���� ��Z��^���T��^��Y�X:�h�Xj$i��1��2�;�_���o�^�q�Efԡ�sȷ�j>5f	,3!:��W�����O�>B�¦�f���V�P�],��s{HwmC,��E��w����l�<G6�]�������w'E�Շ� Q~|Lz�h[�(�e�,ٶX,�ċ��=|�5��)��!"�z*K����3;�|)|9�-�4���¢��ʭBW%${7�B�9IR��j����1$���C{��o|�_���bɿ\��tK���G��7��A�^�����T��O�H���l�o���/>������i�QT�����Ξ0z2e�s%��z�������G��s[����7%���D��+I�����~O&��.Z�?	X���yY��uU�u'I��E}����ĸ甶I%��i��e&��v��Q���J3��X��
f)�����c���� �-9\{�X&���ӯ��E�Ԥ��SJ�`�<�>=�Ω_܈��-�j�z�����[�a��sIe��S��߾�����j��[/����?y������FV�pU퓹Pd�W5VO����Q�IH���`���3=����E�]��m���t�[��/g%�'�>E���h���򧣗҄W�ȈIa�Ah���.,J7m�,zR@�J*�248���*�����S�uB�>��r�Q�Z�b��D/��-���)�U�7[�HJ@v�n�,R#;A'�:��Y��:�W��m�tB����=L	���i���ܙ�8
z���m�,g�i�xv��|��|U��;M���?�>�Y��5��Y|�2Wc��8Ry9����� ~����������(��@I���zC�׈$>�f{?�Q�-������r��N-���O/����|�����R�yլ0;ͪ�,���@�8��z@�D�=~�)�,���U(���
�$���G�ä����Uaʱ\W�1-^c1�@�$'�"��^�OVI����R���zAKak�G�x����z��R9����+�2!\/��eӆ.�և�Â�bx�Xĺ�W�������gWoz�� *l�2��*��ܯ��5�bv�,\��ou(�
:6��])X�}7{40�p�[Y���rux��L�B�d���8��
��/�ʣ�2G��l�v|�`��rw�.���r���*���Q�v^��*�\��$"Y��wYW`��Ho&)�x�%'�"�	����l07iN�dM�[V�hc�a�f [N|�E�;[�:!���^�n�#A�^�F���������WΪ���0p?ő�@lI����]Y��K��1;�^ᆙ!�z�q��BZ����Aeuo��;�N�N9n�g	�x�F;9�.���bj�e�׏E��aş[��>d_\�.�̈́c����n��x��]륷�����(?���
�����ƓG�Մb����&�H��@��>��;�.~��{
�h���{Sm(�� �7�	f�]�x����t��9g5�j����
��"�'T��|}l�~
��#=���\�_t�e��I<lͨ�sU'' �C������%���׀��R��p�P{H՘��
����T�9Hd�keG.Vp�9��)_��z�}PX�j��f�a{��� �6�-���������l���������ײ��������E���ְj�����Ҕf�/Ó�G2^�ο6"*�	8R����ad݈���#������^p̾'H?}e,��]��3h�D��2�0D~�\�p�zHVKOM���cs��=�"j�^�"-c��(5��J$4�)ϔ�N�7�ʏ�v���Ol9]Ljѭy!����"zMt��W� �`?I���יЌ�m�(��k �eCg��g��u,����;�Ȕw㸊=6r8i���>*+l:F��t.�c*�%Kr�ł����]���i����2$�dv�?�{gX�܇$P��)sP���3��)��x���*;��K$!1�������L��G%��ǟ�����Z4#>z8�Z1t`���N�t�(��,V��̨�
��i��7��Uz��>�:�؛��~"���v���M�%w�[�G��GS5 �ϭ�T*�g�n60����φ�����6�({�zE�x�#o���7���1g�])w%����҇�H�v���"�O�F�p�LUB�e����+��hǫ:^���]G�/�Ǡ	��
3��������ځ�jD	o�Qa�G�;�����q�*��jB|H�&��!xt��>I��Z����p��⫗$1E����uD�U}�E�=�����=�2͢��
�=wG� ��bۙ�Ӡg�,�\26`�¼��D��!�r|*,�d���b��P+x�Aa�_����8-l�8!Y+�K��F�eT4��Ņ0H�e�T'Y�%�=�UJ�u��|D�&�n<m�����
��R21�N.)�?��/�ok��#�S�� �Q��H�[�Pҕj��fsf��e���mW�.��ɳZ2d�l0�{d'����t���)�<Rh���캢��w���Ц��ޔ��L^b��F��UН�d��f�����J�Z���&�2:+zk�K	�G!�qޑ��t ��~2��� & >~L�
�oZ�X��NV��uZ�I+�nz���X}t�f���b�D�J�>�>�U����=	_�Gq�l_"2 �e�>^*OT(6�(-Ae���Y�o�PH�4h1��bϔ*�i��nU���u/�s�)�u�0��*p8�2�᫐������5;��S5'A�:�*�`ҭ��R���VP����h�ڍ8������Yz�g&ĸFfs�(�xj
�pl}��v�a�u�F�ʙ��UD}�ߠ�3;
\�V�"Mn��s���Q1V�z��drR�;	)����1�)L.���a�[.�ȻD��K��2P"����_�6�woZ[��"'��K͞��0#��bz�C9��nU��P�j K:m6']Z�IPspP�;�����k]j�$T���Ou��s�������p�gM���3�Y�K�^=�G��6������ii��8�ʭ��|��p�:���lQ`3�-m��ܖ �f�!�$�]̐?�)��h��Ȼ�ǎ.��%	a=�?,�j�}�&^��������f���)�J�-a߹iuS~������_���O
����w�ُh��kU4��5� �w�_�i�x�YI�QSPM_s�r�IK�w�[4�w���Tj_��~�����7.x�D.���������� �N,�4�T[�g븡�ܦu�y�p����4�w9-���D&.	(`���J��-���>cE�K��5I�mz��$ԕ^Ϋ��ǡSw�ˡy��K?Ӕ���]h�~���<֜ �#��hLk�ݛe慦[���5����ѩ�� ��(x��h�[�-��p�:�7F��7_�:��A��zr,�`��]F9����w��l�E���<�=\��2��,/��Q3�WoE$��Q�����;���W�ԋ#� �B�0����oxn�ɰ��z4����-��1�xf��~��<೪��-Bc�5�q�vV"}w�⾧)���F��"R�,<Ox���yi����%��͗���2��"���n�k-r�����l�C����C��Vu)oF<�����(BM��*
���f^ۈQ��Z��Ç������1�(�l,��Gp�})�m�*�"��������$�ǽnmU�j��(v��M9���D���ve6�QT>qp�+,��A)�GZ7.i�Z��3����R	o�n��j|�	=�.�6Nw��5�q_R�� 9{�ǎE�����B##3I�Z�y��eꎂ���p�OBӐ�qD��{*R��vXĲ�2��k�뿗�#�u%���U�!t}'˂�j2c�f1l����{ޠ[�Lnt"�!��8���-���&�����aޔ��4)f>����|�fǙ*�=�݅�|��������~�衹����==�D�ɔ��_�jnn��
���|�\,z�;�]`g`i����9�WF����d�f%��[��� �_^׋�/0E�~�/p��ʾ�0���:�
��,*�G�Xu���4���?�gЬ+�j��[c���*�Bqd��*�f��tt�$}��β��X�`�Pn��\qQ�=U�h8f�E���D���˂W�14�jѕ������ �zE���$�W��ViYyy �r0��`��>�v��)��{J��2���
)�=����������R�v0�7&�f���~��͋�m��Y٠���O����P!l��ʝ��8}c�i/~Z����zZn[��8�����Y�`���+Tɝ�'5�:�B��B^$j��e��']KAܷ&���dsk��5�M�k��sx%[������57�n>E�O�A;�Ȭ�xK�g;�oN�{�ا3�����_)B���m����-o:	$%+k�1w�1𭁚tֻ�+l��N�ԙ��#YC��N�Iw�ΧE|�I�&�+���mL�(]���c��3�;5j*�1��C���u��hL�L4��q�"C�J��:�� r��D���
a���	�gYZ�w<#��y ���t��I�iD���v6HE��E��r�}�����K�<�����FUYr��~Ň��]�	�K�&_|��l�*u���h�QG����>�ͮ�,��6Ҥ�!�@�5g�/)�Fg٘y����S1���4(Gr�l�| �R�)ݹ�o��,���ٱa��V%5��}�	���'"&���\[n�Rjj�ͷ�t��\6��[k-��t��B�����mL�h�u��Z���C���ݜ_m�M �k\��7�tν$˗8\��{e��)c�A�Cp"�*��+V�@�+l��7��3�+g��A�f*�(!N6/AM�;�k�J�0${�5AAG����X�%��xBzo>����/E]Ի�q21Us�r����Ȗ!���K�̱G� �y�
17Dt2֐�7`Pn·�ɍ�z�5�G/.;i˽N�����7�����7�{#���IM޾�to��L��2؋o6���̇��ߦ.,T����5��Y��_(���D��ii�Z>^̡�%>6�,~�@Qtil_�����[�1:,2Bf�,�I��r�eb�D���"�}��{�^T	�;�(S�`ȭ�E��'��C����u�M�B���$��uB���ƺ*1an"B8�أ?a�^�{4���	؀���I�Ou���ax��u�_���^ؠ9(�L-3��(F�mT�-zhԌ8��Nf��"Vra�{j����nC����` ���LM4$���}0��.0����ԛ��B;ؠF���$u���E�c'�E��pY-/F����th��}������i����dE(���	�Tf�L��~�֪P+�������+��ZY�����2���`SKڭ}��Z�o�6-c��dg&3?�x:V��T a_X�+d��s7IV�9$o>�m�"�;!Ђ�_�|X�肐�7|���3M���| ���&f�4&R������@����i��;�"�kA���4%�#�rɽ�$�#ߋ�!l���'����x�U�����d�����x@=�\],R��6�>�<n���W� Q�K�c��t��Rb��a��Q
\tX*Z@�K��My��ƌ^�����������N��-�����R-�`��z�]l\�fŪ~�*��Ȏ�z,*L�-���D�!Ƭ<�W�ŏ_eh�����02��y�	�6U00�fZ a_�M��1Mc��f*bGu'�,jQ�$�̟)�%�����-j�g����L7G\�ۄ;;�"��;�V�|Н����S�$�v_���۳���
�B��լ���8�AHT'%!��p���i�jA��U��d���x���#w�ԘH21䉰!]�	�{��"vÎQx󗦯0���\�6c���	��$�w9G$�[��Yp���W�ʙ��ڃ������eX�l���K-?�8�
<'LB�S��V��G��_<���`�X6�Z��楯���(�iI��� 9�/�hp���^$������'��h�0�{�
��.�D^X�&�A�r�i�'>D�
�y�4�l��k��ɞ����>"�/��H�����{�Zv�yHB��㉭���@	^�2o:B�B����s�G��7ws���E�����V�~�L+B0�M����f_�_s�/,Ũ��,����BtyP3YVy��Ȥ��#o�0�ء0BMP7�Q�2�;ݏX�]�l����㙵y��K�V�T�/�f��C����F�&�(�6;�泴���q������Uۨ�O���]���0g3��b�W�CEh�p�ԥ>�b�JN��h�seсeV����M��.����f�`���E�}�h�Rx�R��V�jK|Q����2f6m�iQbF�Eح�h�S�r��}M���D��[����}�4՛�&yRv @2+��yxU��ò'R��"�����S���m�N� bL�����w�p�������Yр
s
m��V�x��N���-Q�5�
�T.s����<��	K.<,Ūe�qvA�w��a���دl�u����^=x��� ��9�n��)���y��7��X���ż�E'
{�3��� Nt�#*`�t��C��Ɉ��uo���Iށ� ��鈗	�k骣@ly�u-���笿�^��*`ֳ,Զ/6ʹ؇�,�?\��V�wWU(�Kp����.Jh�e��=�����.����/oG�dJ�Tj����w`��J`]X�$�Ɛ)�o��qt D�co�|컶E��<Uz@��I����0�B�Hr��ʪWwe \I�.�����_\�����J���~��B�u��*1�}�}�ءS&�F�A�j�uq�/��-��qӃ��I8_\��}^	����;{�z ��
v��+�K$��������Hvm�R�k�n��&-D:�Ƌ�ŋ�dV�(��y5�0�a�1>�,�o�S�����z��Ю��"0�Z��R6�Z�¾x�1��8DlcX��ң�����e'w~�M�r�� �ejO�m��

rP�E����琯�ʈN����*�� |���2&'L&��A����<Y�+ �����2�֗G�r������T��YT j~�0� ��ʬg n�I�@as����2ǡ�F��gg�R�E�ꮠB�
�P�}��
��'	����' �,s�Bna��4���5�F	�U ��ZI̬�"�1| ��Xy��A�wlm��5���9��� _$�3�cc����[�O���a!��|%�3�/ 0�g�Lڷ��w��r�%(:%�z8�ƣ0cE0����qyN���g�5�c⁘_��e[���ZGo��`x��^��^�YVf��B��]n�v��A�䶛լP��̸/=�J����@x�?߷��*�j�U�d�����q�K޴���d�����љrw����"B�T~��(^x�i�D���/B2T�B�p�����%��ʫ�����u����ྛFy�$N����2)�2��#�s����?�n�P��J랦�u�<h����h4����p^��Ƴ��k�S����<N�(ߞ�m ���jN�,�a�K �X������s��!�g�t���݇f���t�e�~�(�7e��̝�����m)I־\I�sUo ���4��)�L��r�Sŝ�p���Y`�C�n�������j�f��g�<���Q+����C,L�%o �C���dF�ٚo�k��x������C��$���Ǩ�|��gk�y���h�!����O�8��� 1w��a���Q���dE1�~��� !�_�����dү|O�U�rO��mY%lM�?d��ϛ�`'��ʙm��w�L��7����"^]�bOӳ)�r���F�x�:n�lf/�m]��.�F��f	(���X!�bu������߈�t)r�K�o����Y�AR3�M�T{}|p�{�Ctt��k��+W�����?0�S�e(?ԭ.�H�1����Cs�+���N�+�0� ����`����w��1]4X>U�;q��%zO���LƆ���B�vڶ�c�q�]m��bO���.���+�l��/�U��Hk�k'�q͂���q�C؀��?
����4�O,uh��'�p���|5��*N��V�o�Zq��턱����_�i&����A�q
�bB@�Ut�t'��L�^��J��2��Qs�����V ��af����ŕ0?�}��/���g8�)��KXm�:�ŵ����p�S�<�R�켏��K�;3fDZ�o˝�������(U{��=�^}Tb�����{)`�� ��䙟]G�'��:�؜�����5���G��P�s27�9 �?<�r�Ob�V�#hұ�_1̥9�]z-<k�d�^Oν���I{y�V��2��WS���&Qr�=Do߅ S� .�!�U}NN=����T����;/rd��<���Ǘ�I�T�g4�4�&�I��rx�уY	�I�a��~5����^��WrS:r�h�L�f�,z	/A�9�����s�U��͕���r���B�-���2���KWD���
$��G�Ɏ�	b���ߛ�iH0y�˭dM:�;���E�=@3P*@9b���Eh@�VB�.V��Y/�ƃH��'����"�d�L������X>��jQ
d�y��N��4D�� 7�|E�n��m�,7��� 9$�����?�Qz�W���c��wgĳ��o6�U�4&�0X{�0^��g�X�F�9����K/�A�f/�$Ck4^�$��<�3�h{Ɇ$n҄xZ"��hwޝ��yg�l��a����W����:��B."�ˍ)՗�o�^v��h'�&�Bl�n��"�p��H�����	9[��@�V	�Kn�,K�9?9�ā�R�Im`�֕����:튢	��mY��F�Y�L���A~���p�4�hoiq�����[����E-��a9�;��yc3y��X��=~�!���E4,!p1�7Ϗ��,W1�w�V�3H2x������:z�VTe2���G����%{t��$���o<�����=B(	ݡ�Zީ���	�.Ɲ���^	}��Z���~֘��௰�  �Aι���;�+X���5��}fŻ�@�3p��t�{	AO�J�G�� �z�4�e`��)����ѝ�
V�UH�U�~\5�h�3������7R䖮Dj��Z�4	��߳�f��Ʋ����4@͔��)I�z雱?�w˒�����UX)�P�a"�"��k�$�^�	A]�/i��y?�(��}DH� 1�W>(��x��-�]�^Y42�&�?f������_���1�dlR�8�E0uAO��#��W>j(<K��i�"���api���vhΉ"�\§Z��bG
�����z�K�
G�D��v����6BiȆ;4S ��ܢ�2&�`܋HC��Hn|�h�i�s�K&ة0I�}2X����e��)�-Lr��,r)ǆ��-0�|S�|�xb����/H�MN�m��r"U6	��lA�����LTie����/,�ߗ�;�11����Qx��0�3E9Q\wϽ7g��V�W$�*�.򙼩!�]�CeV����+����A��`)g��l-(��O�O�n���\��y��v�"(����00'@���e^��1��C�Σ~b�����,4��r�� $��v�DZ+�������3ϜpUW7Gd<��!:ը�g|��TD��ҝt�%�)ԤBv:�0ڮ��3�V�U�����Đ��>�dTy�Bջ5Э@3o���~pQ��$�e��"�(�_m���t��#Bs�+�������|���q���kw�x���P9�׵f�v�U��ԸA*g�`���5P��k�`_�孃�^Y2E��iɅ� 9`�;O"������|6!ޏ��w��BH��}צ��7�m�?Up�˚榭�`p`���,z�}�Y�!EǧG)KǂѤuZ���I��띒�-}�x9k�0��='猗Lͼ^�i�u��\aԧ|j#�4(��^�{�Ȩl3�����>?aP�O�)��N
��p&%�Ή��o(�Rt��D2ҩFoPl�����Kѐ��rS�(�:�Y@���>�X<�t��VZ�P.�8���% V�����ʬ���#~j�t�����O�rT�^3�����7�U��â�)
r���VʇF�<<���rD�htt�/
Kß89���!��IA���m�9����#i��жNBi��D�}M�G�A���e��g�9Ţ�u�Cv���&Ur�}1��T䑮9�g�Z��Ş[��@��m�=(9�=˨�&��T\��D��w�넽�hjyN� �߰����3��p��T�2��������Z0�[�2�$�9�M�)�E�%7X�;��|,�Hx:��o5ғŀ�ӊ-9����SOfJ*^�N�U
i��{��/�ʢm_�Ǜ�����r���'����;�e/V��:G ��n�M&.���1�2v���3++%�ie��0��Xj6�i����^Ƽ�6��v�Y��p̐�@�R�v�c�_ԱNv�@�)�mrk� T� L���C�P�of�J�s/S�f'�v�ʓ���z��Հ.�b��.�n e^	����X����ۣ�6Ya�ɽ.m�6��.�c_�t�y����5y����8���);�Wmn҃������4���l��im;n� B;�}Ne�����?���l��B7'%�ۃ�5gly�u�-��4�F?���e� �_YK�@H<2�@�B+X��R�,\�j��/���n�W�����4�ɭ,�#� !���guK/NP����;��U�:2h�v ���T[+�+caE�..��.R�He�j�٠���{fnT��	���BKt -���9���oh��A�Zj����ߗg�u��}B����&~dj��p�xM�����b�{
-+�2WUVIR�����Y}�Kp*���Y��'��ڠ,S�
�8���������d+�M��T�tw%�p���Y���a�?�f��A3{u�����v���S?[�u�,l�,k#C��ܗ
�/"؁`C {X���$�D��u���^�T�헆�o�+R-��>��6w��N�j�pk�j�f�-��_��	h[C|� V�y�7�3���I������K�Zu�B~�/�kZ2�>1��b}{kB��o��z�) �Ӈ�![�B�g�� N��׺����=�\5E��Aa����~+#Ǌ��|S��i��y��]b��K�z�u����.g����H�mEF�
��v�����/G++ �,gj�c��hB}lt�	�#nDj�6 *[��J�ϰ��p�!Nh��e��q܆��i���;���s1�A}j8���z����vk��񃞔cx��j�@�wJ�x��^���'�I8�<�=�&* �'	�` �w��p�g��*����nڡ֤/�	3���\��`!6��/��P0Ä��}}C�m=+d�(�oĽ�ښYV
�6W��'c�&�+�c!ln��u���o��Gy=S����;$�|��i�o���{��������ȁ���%L�X��t#, a�s)�_�Oq���Z���cܠ:p��
Aj�>D\_�,c�߆�	A���ɽ����|�F++7:{%uD�#ϋ��U��\�؅P���n�?hW-�{�W�F��c�R�w�V���2$��D=ū*o?]�]w5�,���#����0��T�!|�Ys�V�"��[�{�c���/�x8g��n�n��V�ә5��͐Ő�/吢��B��a'�[}�����-�Y"���4��[�����	?���.�9�nFz%<g>Q2��"B��������� �hV���F�bbi�g�����A�G'|j����H���4�u�v�,���tT�2zc$s1耭3�R���m׽1�#�.�?uQ�G^K���+�Je��Y�Ц�Q�6��>Y�7����a���L���D/k`�\r���W&Z��~�����z�S�o�'� ��ϧA��c�2���z����"�O]��Q�$�xm��e��ye�&SG֛WL<��^_]�t��_���<�K�]�$Z�V���h�]����1�`�NcN�|d{n@u}9�[��j�0�f|q�vo�`�Hqc��EY?�5����t����Z����1��%�(�"J�Ƥ�%3�>��y����S����r�E���v��=��ۅ4&���h՛�'�tԃ&�_��*-Z��?�f�P��iX3^[dNb�[͟��!�
��H�h���s��y�U�> �f`2���"��|�$�1�'��M�p,��Tƪ��g�aK2�ܔA�B�F͜YUMØ-	�HQ?Au��W����IՃ��+I��%����
�ocZ@�C�$�v۬n=o]�Ư����Ҙt<Tr!���S�Ø|��HY���~�ƫW�i A ƞ-��k�N�b	\�K?�b���|��*͜�:�3%*S�U�Ң\ S0����@�'hG�
���`Y�z&LS��S�����<�R��䅉���l�~i��"��eL3��ɪ�FvJ��ys��WX���{��N;�[nU���d��Y�_������]���Gy��o Q��>#�q#3t���Nh��t]����G�R���"�%;¶� J�H��I���Txݫ�g6'���)�jg6��7�|l����d\�|ރf2du�mm����Մ�x���:!������8-��q��~�Ơ��y�K���E�Hu�~��h�r����]"��.&�b��A�I���T`��F�bv$����:"O�9t��z
�ӡWKc߲a�g�%$���2��1�����HEU�HD�޼�w�~����F��C~�EV�?G+�`��(���u������eؔ*J:j1��t6�֊����4HA�����ۛ����Tbb���R���"�0B�*&>���H�6��=g���̅u1�p���j�dy��a$M�/�rW�3� l+ſC"#f��9��ہd`�.���Vq�`'��8��RMb6f"C��T�M"m��܁���yC/~}7#KSnqT�n�d.��)�m��`<�ģ�LE.H�a67@�n��~s���`\�K���;'������4%��9�$�*�梅�3�c���C5DO�p��"��ȯ}��3mI%fn7s
�|�N}�i��ߍw��\��$*�2*K�V��Cp�˃�j��,B	�r��g�M�Q�!�,|v�K�F��0C_aJ�)c���y�&ĒY�Z��㽻:x�?!z��"C�t�v��"��/v��9��@�k��z�8x)���K�h���nK�i�YRb��Cye�8XnH(������Zb��Y��N�9�C.F�L���U��RAZ�<^Z�T��ҫ}��Z�8C��oe	;�\L�Ì�l�j�i�%�Z���kI�����x����} ~'����օ�]#�W�9���9&�Y!���'� i��\�D�]�wZ�=d��;��ݴ90X�-���Al��)83�#Y$��������n�q��:�|&�(E����Wh��4�{��ݎ����8��د���p�K���>6� ��	�D�V����7#K�0���(A�(|O�����L�����^?����/A�����
v��Y��X����|����<�_$5��}���kf`L:1�Zr�'1����<xz�DU��*�R��g m�x#��s����N�]}���GL��2î�6��"�\ٚ��!��o�����T�d��~��M=�N:M��sԱfJ0�˂w�x��RO-S���7%h�If��=��<Ky��нJRЃߏ�����ʐ��D|�=_����4�����}�m���i<���]���m!w����R�=ȝ."cz@镇��d�H���D%Vqdl���?T��e��fӟ�=k��>3"�3�FlO���x/�w�*�-�8��۠t��EcP��������w�X��G�E;�:���0��� Le��b#���3�b�ڌx�)���v8�@��?9�,�#�����V�W�oA��Hf�-��3���Iu ��ʣ;��t[#�a��b��maSq9t��ϐ�Z��0�����ǖF�H0E Ɓ�0o�vCGQɿMP�?��g�3hV�ژ����~�DS�ʕw��]w�y#��ʡ��_�5���O��o(|rdL���QA�dF�����U�ƾ"*�i���0����ǹVl��I�X,M�ת9�d8�4�-�9T�A�5�����Tm ��͓;�	�+���U��]H̙[�]�[&�<㚶/�7�N�����QA��k������Eh��%�ee2�Q���Z[識�����9�*��,Y�*��W������&Y��%�x��o���c9�[�m��<r0���� ��
E��<_9z����m��z�9R��ȣc}J)��i���+u2�v��E��{���\<�x%D�]�9t�5��pp���A�����]D�> z�����o�r:[z�?�\#ﱖmZ���&�����cj���s���N �ge�pW9%�=E�9\�hqz�'u��/K?b�폜;�6�(��'q>���Xt�a���)Ů�n"��)A)X��-�`��������r��C��?G��^j.�)��Vo����1���W���y�Ђ��M��ڐ3���!Cf�\�) �Y�eoG?q�v��L��1p�u�Z��/щa��?���Ayϯy1�u���������s�	��6�����E&;�%`-B�ŧ>c�#[�;�duHG����biܮ��[�%�У[1ڤ��e'���2��J�����:����v�I�-���׮hk�jb��y��vh����CQ��u��<�*��Q�Ũ�^�f���/� �����E�=:�,�h
Dt�w��fv�L����"w�}w�,�����P��m���=^���\��K��o�gW��ڢ�ei��$�6otx꒚t�:��L!��G�D.��t^ts�a*���/��t�Q$M��[���(Ray����ѡM��g'X�O����_T3�⯻ <p�/�VSo�Ea|VS�z�]���/�9<�lc+A�� y:����\Q�⵰�
"/v�����J����F��#�1�����V.Ӳ(!#��_��`��:e{����%\� ����<I���w���)W�E@Ϲ<��å��M�l�{�+Դd�u�!�!ZTg*��#	�V��ڲ%a�t���N���B�x��0kfL���I�8��sv���R-n�p8�$2���p��J���|�uz����e�ɸ���g��⑳Dt��w��؉��x��^��4`]M�B�ev���oέ�9>O��F��$L�8�z}������D�~3Su�tG��?u��bx']d�|@�0*�
"�*^p"؀���=�$�wt�@c��
O��o8�amH���[�����W� ��O�/��1��7q��"B��4���5��b���&/�%7Gܚ;O5�%%��Q���np�E�`�-2 �#~�@q�e�$����2�'Ub09����p�#<��"C��^5:�!.f�Y�8��е
��#��y�p�"
N��ѐ$�vub����m�e�P�q��Y-mZF?��Mq�F��/e@�>���s��G���-�T�w��g�s�v�0��k:���ÃWCE4�S^~�ZD^�QWN�A��i���ȁ=��wy*᫜�tf6��������O���Պ$!|�5�Y�Q}�hQ}�Z��4M�p/g�o9d;h2̳���x�6�!��
20ÖY��bfџ�q�%�y��~�N0������m)��6*���(c��&Z�k��[M�o�xc���C�*F� ��)@��faA�����}���!���/oq�����aHq#d��Z߱�D�A��
{8��:4�q�튫�P&��I,;��X�N�H��8�:�v�$W���kmSx��C!�C����	��}Q}�p�iq����ψ�3���7`~��r�,c�߬YY|hصF��1�oι�QB.X)��\�Gt�n�O��S��L$y�H��}��>k:q����������@��ieK�ܫ?6C6ǙZ[7*=dJ��	Y��/shⓢD�3��(�Yn��(���~�6w̜������h:8jv���/���rJ+/ҁ��o�̼Ӽ�/4�{� s/]�k�{�Aw_���9w���k}>�k�!��H�Q�6V�M�Е�F��M�����k���-a�g��NNM�F���XԖ4��C�e���"� ���JQi�i���K�s��ۗ;�� �k�k�uv��$@���R�E�]��G�V�g>[]_:A,@h��uc�p���7xOܛ��ʾ]�: S����'ck�q��)WGt���+��ؒ�G	�y%�|�q�j���͝6�?.N@?�l�V4�Km���N��a�<��2\�� Ü݃<޽�*��{B�ɏ9�ц7���!�CV�<����gx���Y���f�r"/�@v�
~9�CF1߼�)�Z�' �A���`���v#Ѿ���_<�҄�j3�4r�{k�=����+h2"��n/��2�I��d��
ײfl{�ê�ʣ�%�QE�(�_�����
��k�[Zm��o��#�b�qR{'o����l"Vd�p9�0�NKM��uCj�(U��:��k�T�(�[HP-k��M�C~�����O�]:�s�w���F�U�P�hc�<�N�� N/�'C���BXnX�z���ʷ�v�?�B�/T�Vy�ܗ�����(o�,vR9�9�^����A8�t�r�M��nĎ1qc�t�%^i���Ǹ2 �S�cE �@�蓩b�A��BN�R�I����Q�}�Gn;���� ݌ ^9�BĿ���Jf\Q�?r)��1�p��?�t��{D^��u�楡����)\��%��^nd�������J�Y>U��_V5+�h���}+GhLR�С�����!Ж��ر��R������IR��[���TT�B�S�̹�_?�]��U�7�ꭏ��]�X`gL���9�Y�� ���8?�y[eg6p�7r�,Dh����3��UL�,d~�����(�I"�ם>��k45�`��������8�l	R.n5�k��1�.]�0g���vtX����	��Y��`9��<�(��!���p���k�c�̞�(a�܎g�y0��N��c!��HK�D�q�qHgot��k��II�y�@H&����+㵐(V��%�Iέ5��=;rH �4.�no��Z<�6�Io����OКT�n5D����G�fә8C���f�s������˴�Ȯ^�/�f���4ǜv�� r���僧W����0S�\��Ǳo�Q�D����v"<=�P���v����������t�9�'"�va֌(HŇ_(��������J	�sv�ލ�QrgFί=�xW�Bw׮ �g(��#1%3��4h��z��!e�}r����&���Q��:o0]�`EB�pSC�YS	�$|5b/�9�{��[����r�͔w�*.is!��o����-�6R��,NSK����,?�L�
hՀ-��.�r�ED���C�R�����Σ�ab��d��*�P�t��ys�YI��S7����{+�M�KkDL��pY���T��!$L���ZyI�k��� A�I��!���j�K�-��=��T�#h?�ZU�*(�Z��L��|Q�%�Z�-�v5fu@��B�TX:1j%���#����3ق�Qh˽F����P��"������ȶW��Ȓە�Wmѽ�n)�XS~����L��&..���׋ (��KV��g��֑H]�6m6'�ѫԔ<�|F%��	�%3���y�}pq��#عe�ˎ)�Ȓ���j��n�=9�r���Wkϡ�H����#~��₆���z���|\Ts2�5@�h@�\� a��|���p�[�Zx��@��H �H>���d|��P�!ʴj;B=�Oբ�~��P ׼m;���%�\ˈ#0*����֭,m�ub�������7ɛ���3�[Jg��%����o����~�C[ś]d��я������眥�!)�e-
�s�z��$'t4�H�!n�7b�7��b6U�Ӷ�:t
F�^
%�u�X9���I�4�̤T�y� {�ԉ�'�*��u+*�JaT�$"Wy,;]�T����oa�+*��B��Fks���3Pk̙P�:'�ٍ˛|��d��������S��[aV�*�v-�A�F5�=ċ�Ro����jᤐBtⰫ��/���;��	k�� {=`uR��#�n�����!,C�o!p��UpC�i�F�I����r�7�/"�#�Zw�L��g�iLH0ٿ�oiH ��'o�ZР�̴���t���wn<R�th��k��lT�R����οH��x��ZИ�� FSg�{�@�!>Up����[k#��B,1Nؐh�Ү���JQ#�����-B S��"a	b���o�6��z���tD^>H_{��m[|�u���Z�,�z��^6ޯ�gQ�����<se��񃅤�M�k٢m�s6"{��\��]iZ��_��#��E�-��[Sa���
�������0�hC����}:l��/e]%�\մߠ��.�U�+3�ć��U�Z�h{�D��YI0��f��sa�y���\�7����p�� �]G�4��� ��޽|��!��hV�㋥���>�O�Qr��ܼ\Ƌna�<!��>�72�?�ɑ�+��|���d��2A仓B��s9,����4��w�meN��7c��ւyVx��%�� �&������7�+V��ưn��r�g t�@>��dz��χ�@��-�<�Y�����ݣ���ʫi�[�n*�ޞ*u�:c�	)͟q��Osg�Ⱦ>��%��D���k њ����o#��1m� @؋_iR3Q魌�a���_W�yߜ
�,���E�N�x�H�d���#��?bV#"+Bp�����"���e���"�Z�!oҕ�� �7�K7A��͂��x�B��C5 fM�Ŵ2 h�S�#<yMCL8��	!>.I�*<��V�C���!`����1���f?�@�4�޺m�)󾜃��ΰ�l=�b��P���z��4�+#k�c�s\��rw��u ��|_+"�/n�r�W���@n���r�v�E&��y6���]-[L�5��q��U��|�^������b���J�63�m5����ޑ������˾�oh��OB��ZRd�)d,�=`z�w�t(Ϫi���h�,rX������q��e�Pµ��N�DvZ�ےЍ�w��צ|�j<G�	�HRc�k"8U����X�i�C����M����	&���Յd���k�D9ܷ���~�vmU�K ��u9R��Q|0r�4Nt��ʜn�[h|�����d*��TE�6�l�XC4a���Cu��8h���j-]	�y��q�}�H�[���2�g1�K?��	�ˡ2�R�ͮmdW��V�_I9�0|Y~���x��&���T�@}'�.u╡�?���kN��ZM�2���.:�:ҏ�c��ꛟ����o��4Zp��3ٗ�Gr�[���go}�kK(��;��>�L�s�^�R�>�CEl*�	�b�Y��z� ?~fD�����>�:�j5q���+k��^��4�+�i�hUf�¶q��I��屔���ēQz$�T���x2��$�V��ݴo�l_ڰ+>+1t*��,h�&�/!�^�`	U���dBf�U��i��!]A�&�����e�1�No���.`;���kC���˘���*�E��a|t��SZkC�
�y6���sy���[ E
���'@P[4P�9��A�0�=Ƴ������ 3�k[5Ƥ�z��������O��1rn�F�k&S+��I���b�Ӑr�_�l$e���!��d�q�:&��ܜi��"!��q�r��Gs�^�PCE<�<h �E^m�EC.�] wN��tq�x��S;y�����	��8hq�c@o����L�p`�&��e�3%m	]�����ix���@�R=��rߪ��q4;�ͤ�7��s�$�긓�~3��|�D }���bo���� '�X�o���LK�ڴ.�b�y�Rg��2��s��Č4��LK��+��?s+.�x�}���*`0�Y�TS�}�A#'�sB�l�Ds[�
�31����nE���)�,^V�c0�����	�H���NO{�0�q��-��r�"`g琺N����a��KI���f	'�t���١�e76�ؿV��à�7@��E'�ͺpqO��u��=��>�B"����A��KH_����w弨�f^�b�۵�/!�OW0�4ՙ�ND"�.�Ǜ#F��<��l�ӟ��Zh�g�A�G��]��}n�:V1�$C١�2���Ӓ��_���#ԯ��٤�����Y��Ag$t
�|/gG�P�wm�֛�W��"�0�
����%���-�rm�J��w�"8���n�l�y��lȷ9Y'?���U�����/v��4��ۏ	��M��Y������w{��p��^5�}�j� ���tA� �:�lbԯ$ӫ�Rހ��s��prR��^&@L�P�<M��M��j�.S�.~g�W��'����{8�nI �ʂ�H�-�a�Ui>��vr*{�@���;/qFL������쭲�6R��	�h�j���
��{��'���=���"�wĢ���:���(���:Vצ{�[+� 6�x	%B��ce4��jѻ1<������q�fq�Th�\��=����V>���x���,�ǳ
����� jC@T分;�/��7^Ҋ7�@#���Z�'/	]=���x5���-�zK"���i�+�#}��w��~ϭ	ꩦm<�kw�����<�Q�.���.N�G'g��H�RL#o`���"��p=@��Bg@�=�kS�o�+��e�O.��l���0k~W>�3����s�bL$d�� K�Ĺ�ixA�&�6чjYqx�T�@2��jy��/�t�R�_Yt7�e���f���*��fm�-��<����E�S��/L���?�>�k�]"񆈲����!ʫ&ބ���'�{?�	/�X�����v��T;L�
ϱs3��D�޼�T�#eӤΨ��P��䑙㽌�*�#�k�W�"t�5���!~G�,�,�OY9w���=|�C�o����e��7s��Tkw�]L�q� 	׆��)�K�cp|���G�Zt�`Zwvn������3#����z��[p2��<�~j���J�	��ņj�c�V��m�KRF[�i@肠aBL2ړ�x��֛���Z!��ڨ'��c
�G��X|������%\w-�� ���n�|���Bx�]����W!��"^�����5fuT�ӊ�_����fd�D�����	oC_ay(�ୂr,{�1����!sָguH��4+�Yěx�W Jwֻ����I��B��L`&ޙ�������2]C���2�E�=���UU��𷃚0Q�(L^M0�̈p����1C�F��n�.3`�d��Y������ix�czRD����Y@��́_A��ޚ:B��`�C&?+Pᘧ*ϓ��o� �M���dR��D́:�~�P`dH�ql�@�F�Jt�YMmO�_(�����Bc�Y�}K�RIq�G�����n�N��/R�	K��3�(���fj��K�$,7M��Mc�1)�ђP�b�^���5�����i�)od��h�0�r�/��Τ/C�gt?��g���c����O&�ۙ�֨���0O��@���8'����z�û�zט���,y~%���=���Z�D��裇z3c�ҵ� ^�^�c�1��v�%����q|�(b�D�%hO������E��ӷ�/�%*�l���`�˦�����T�U���Q'�.7;�V^R>�[�� ���_�6r���:z����g=?9�2���=��Ul�9��d{L���'���q�{,1~`�7����=P�e�ڭ����'A_�4,�Ԉ�A�{���X*��.M�KI�E��:=�$o�16h�Y��3�����=�G��5zG�U���F�������:���7\�sN(�H�9�r�� B_�R~5sH��D�F�٨:���L�=��~� ����t�	�Ak�_��	�6�Ag����R�y]d��ǣR�%֠8h7�� �p`�v[	lH��lؑ�:Z�$_㱙5���{x~38��+�苽��=�s ��~����D�朗fHb:��O�H����7��y��&�!�<Q���U�FFJ"����r��cr�^rJ��L���G��<��88)�������cL�u���7�&9;s���?��� 6�N�Л_�#,֮\6!ݛ(�x�˯rV]���3D��\��'\�2��T}l�ɗwڢG H�}ભ����s��j ��x���BҾ���6�(nX�+�:5�@Qr�<`�!�ZwIc!Ч�z�8���=�o�߀�~���Q{���3��ce��*{{���WGI$q��&z���e�ZX+H�|���ܳ-m���e�����F2�>\�'K�ҕ��H	p��ۂg> +����ו�M�;,�O
��Zx͈趲b!-���$����c>�T'�v=��;\��=��p��m˄�����Ku��4�3��{L둍[G������
-�&��e��؂�	vl���?[|Й�@`�{MP��!��p8����9���eW�d�����q����� ��K1��X�s�cI� Յ�
؜C5��&�?P�X�}�z@��)��5�I3��p��h��<U��D�۷F %��aآ�t�F�N��|�2D���皡<d�Ϣ?@quC�?�t�B5���q��5s8Aj=��f�4.��6zPG#�|�s�ĕ��f���������F=p:F�ۖ����A3J�KT�t'/,5���r��T�2P8c@ �c� b�q�s��-B���_ϐ��>cӭA� �R�u~�x��ک��^*ut��{]+�^�䦓���N�P�˚^�!�\�Gh}b�ua��I �`>s��a��.fQ:���e����B���+�v�s;�['9ƾ�w���*����(H.�[.�z�f�����N�C��'X��Ț��-�G�;�o�ai�!��R�euݶ�G^ıI�TaP�S� a�E�3o�-7�w��Œ �X�Ű�68��Ȝ�Ͳ���q��ρg��"��|i�4N��Y9Kq�`!<�I|r1����gV�y�?��b��v|M��M��\mҼ�S/�p�"��y�d���H���< 2CGH�#(�	�_#�,�%)���3�!��\�߿�(������M8@�����K�{ؾ�N�&c��2��ͺ��,:s�˂&
��p@���οi�>�jꗻ��u����zH;��R���`�B�4#`!_#
�}�������p�d��w�$�{(�s	18Ț��xMLl ��MK��Fu�;�ǠAQE�.]����V���k��%���vK+�g%� ������#�m�(z�%L�?d�ٵ���6ُ�϶u�q�@}]Nc��n��őKՐA�ͣ�rPR�:xL����{`jx��Թ>�N@u.4h��OXٜOz�%x��`qk^y�N-�ɡi�D��Y뭛�">�$}a���������=��W�$ :p[�v�0c5!��g�Qu��C�G�@l����뚖q�&.�	�2��C�y�-�W�V9����f�������p[{��������Mk�h����uT;�?0��K�n��ʶ�I����8�HF�����G�Ll6��ɶ6.(I���z*���Z��7I~�=Y��tA����k�W��lR����#8�g�y��E�b��}q�3K=`���s�F)�K��Y5��Oݬ'q��F�v��Fo=i�Wƙ���
���A�Vt�����d�h�"�ߍI����+d?�y���.�͸�We�)����͐�����@},M}�W,�$�ׁ�mmd
[Q ����9���|w}�r圴Ka��i�s^Vz4�K���cҟx_��2.� i�xMG���v������ۊ(����wQw��/��yu�P<���l@J��x�� u��@�x]�E���uLo&a���.�e��ݶ������y����^re<6[_�6
[���`�7~�e��6~�� c�ƺ� ��9����i`
��L��z�o��z��k��^�r�������Q��ˆʗre��؉)s>����Q;�H��?�ۮ�F�� :X���yl�?^~�ȝ>Lի���@��]��Ľ�M7�<.�s��e�T,�D̢����eY����L��F����7��͗�v$���݊-y��ňR���1�uF��d��4\�7��pW�O��>����� �7n����2#ĝ����o��N��� |�8�<�9)oj>(��/QG��Tb�����E΂�C2��b˷��]�5��=5�,�`	J��*�ArVpI,C{^~��.7S;�t�r?*��'xN��� y�YG�3u 7���+�o��<���E[|B{?.��w����3�&)���ӟʏ�bj`A�]�5u_�7������"�a�/g���w����#��.�5�e3_f4�^�?	F�W�	O�;.�7'�#aX9���	�qM���<��F��8����AN�06e���| �#pp�(��}���N�x/Ud1I�s�10T��n�������ȝZ����.��Dv~x#ӱ)�\��5��W?RqF}���D{T�.ZzQP_���cs��13�"�kI;V���v�>	�˥���QM��z�@�9��p;�]��yB�����#xlt4H�ѩ
�{mu��e]���|1��s_����uLQ�G
~�x��$���{�_��K���(ͱ�Z�|�L��uӥ�BM�w�����Nد��S��b$�	nj�pMߣ��C��o"'���=5�@�O��s�#�8z�1�%�]:��K���6��݌{<�D�?HJ��� ��^Ƣ$%�)� �� z��zh��_��H8�x� ��i�z�ե���HD�W�>{��':�1~��RG*w�{���$o� $��3��Nh��A�#rq��o�G�����{C�%�M�����ߤ6K�:�݆�
Fn�m�x8��?6o�C똌Pݖ�����}�4�A~E$�h�,�&�r�$� ���Y`'���Y�`��wuN��e�3 :nsB��y�ϧe��%�%���V*��R���b�gv�kt&a^:���dB=�
L��\��
ϰ������>q��{>0��6O��.���u���U������j���^P���%��G�>��&ǚ��S�znTH�]q���%�۝m&%&�
��:GG�jA4��e��3���`:G�Oh�ק߫��`�����2K6��h��2=���#	��g�N�{�k}�?�m���J�V�����Ю1�����tR(2SX�L��>Rpܩ���{�޿0�9Ł�N�>���x��V�Z�U�[N��/��*�k���P� �W�	��L�%�:����u�蓌]si�?͡ɒ[�]����X����Pq�FC�a<�f^隍v5/�Ż����܌�����kb�ؤ^��Qt!�iԣ�<Tb��r7�;ǅ��@9?2�n3fA\�!������̒J3�nO쥊pB��[kH���^1��$��v�p{k=i�i��}�̵�Y����5x��7�1��ݬ�|�~Ra�I�4�ߡ�8ڍ#l�GV�瑲���3K���F�vÿsxֶ�N5���'��?��QO��������7�R�����X��zs>Z"c,�<���&�}��w;{���a�%��/�0�k<oD�j�p�n$��q�R�i�@Wd�r�n�u�����{���⁸%H�I٭��ŔލD�a�3����q�TLp��ߒ�R0��v�0
�Y"bqZ�Ւ�u��k���3���'��#��ʢOE�\_ .�ߖ�w/�Fc�Q�+�4<5C�\��z�8���FH�mq߱[��0��է�*0). ���]�#S���㠜�����%�ذC5�ឬ���L<C;̈́��\isl���Z�2x����$�){(I�Έb~)���5�7v2��醲�_ʗ�7X��
/ͣ �mN��r3[�~x��1W��X}��ʱ���܀=Ԯ���?k��'������ڊ�����T[���o،3<����(�V��9�r���*���ڈ�R��f����pNj^+Ě��@�Յۚ��W�v�蒅ſ�4�9�Pɡ�Yd�-�D)|q����j~hvB)+����K����@~K�4,
��o�\,o[��p�dO��Ɉf�8Z�<��=�|�J�����xʾuF��F��&U����9"�bL:G��o�U���o�a<j��orf��
j���4 �T��~uEr����`x��4���d�b�����&s�8ex�0ZTj��o?͗9��EG�-����י�q>`���ܞ�{�Bs~ۇ��pۘ�*�*5��m���Y0;1�}�"��[�G���HËa6��	S�'�L�&smw�&c�gC{/5]�ێ���Z�j��9�`j���1g��N��7]�<�~�1��z�Į��n�峏���c�a�<_F`����+Y��u�B�S����H��Kn�;�@3�r�m�_@Fhr��
���;�E��i>�V*-��e�R�<�~�E=�yv��k��#��~��}�(��.L�^5��X��U��,�`���ˊI�ޫ����.h��"���nD��5k,[[��q�/�4�4'��)����N�E[ _p)(H䁷���u���0��C�� ���gL��Iu�°k&B�v�ۉ�����qf[��2�Eſ��$���J�';�.��^F��6s���?-���ҏ�k<̼��¦?���v?b*^w�4'.iz����L���D��a�K����hc�0j�م��w";.S��%�)�)3� �<	��9G�!܍`���'�S���Fy5|�mL����9�sd�
��lwh�)6#��e�pxV�9e��=�iX=��� 4�W��24f{�yQ��2��0=a��Y��8�M+Ǜ�����ĭ<�a��G��wccU���DzB	��X.U`���sE����@��O���y8=,挺���LT�9�z�3�~N��3��&�� ��eH�<��TJJl�ӝ�.d3������)���(, ��c���?E]�l���`��_.h��0�ࣜsiSl%�}�b�[�E-��	���{�ywp_o�#��j���~���׫dj����� ����@ 0����A��]=L��Q��·�^�PuLd��A�!�P�(��|X=G�}@݊����N��P%tݣ\�X$�-u�[�c�Q��B��Me�\?��:��"Eq�rl�� F}�"?t��k2 ��+������$�����]��b�A�S�a��~�b����?���z!kR�{S���X�"��F�vH� �wz2��z���X�E�_���U�؝��� �����Q	�5_G�h#䜓�ڙ/ �ɫ�|���L�>nrn�Ћf��t,~�?��� ��)v��@e�I˿��
@��P���R�2Gi{W��s�ϳ!��M4��h�����Mk���3���!�Ȇ�����.И:�'�æ�)�C^-o�����>��&	T�$�Ӭ����<����񍎹�y�5):$9��8z(@Vv��/B�ݵ��k!5���p�r��S��V>�u3�ɾV;�FG�6��Ã!�h�P��ئ��>ar��_�'���ȉ<>)b�3���s�c��P�Ц�����Q�:v�Z�rʿ�V��U��k�T�'�~���V5�SV�P�%�Ǻ����Rt~��,=�W���&-H�=%�OfFcJ6��tA��aD3�_V�B�G��"5��8`1�v2��Ⱥ��3.Ơ��2�ǽ��\����eT�V�f���=�TC����4=!�\)�g��d���w�"o�0���3+�z����2�'P�AK�!E�c���k	tN�'�H�p��h�9I��(e�Y�P����f�,Kf*�ob8UP�#�NkiK�T�����׍�Q��gX��a0��u���w�*R'<�'['K��w�7���P¾�t|�"�3���P�F�N:mխ5����������w$�����7�6�4� �$6}�zV�G7ĵՒ����ɋ�����J󍿓Z��ȷ��=�?G6�	��x��o��
��e�ܹ���p�e9vv0��E
_�
��W9���:e�*2�j�p�V�g[�e `�5aPDV$��79��=���t|��?��R����n�4[�;r�+� Q��>��{ �ǐ]��z/�������qB+���,����������XO�?Q�����*�`�%}	�bg��غ�O�4+h�х��b�p,�j�	�w����(̳��.��ǡ(���X�(�M¬���(���W��P�/Oݫ�V���V�Jo!����y4|�&"�ܗ����1�8��3y�?Ŝ�����&�x ���ݹ��O�=�\XL�3I3���O�,0�}��FuA�{��O��oXtj����o]6�̵$�v9U�%4��ح�CC�̧�妯d�eOӫM�:�,d��T����4z�N��{ٴ�O5 6ʻE��ؽ1eaWƢܶ���߳�I6#��Xx��@C�h:T���)�����0y�ϝHG`X*_�ؚZ��y��`=H"7���9
�,�V�Q׆����x$a�H�#n��u�z�%]7 �4��H�^_Ł�)@��8ލ���ӥ+ڙ8*�0����|�	xv��q���� �`� i�%�&g	;O��QD��5|���uNQ���c�ؘ���^�n�s�o��v�������������6�&�����%N����Xo��~ ��Nމ<Iy��������A����W=�ϝqW5ͣ"��.C�uW'�yF+�q�;%��HxF�$_�r@�P9�oPM�󞃵�P��E5�%��o?s������F���YT��*I߽�Ǣe�Fu+[Wo�_?�X1�+�&7�9�w�F�$o,�L�n�V�66>�CMj�������VV�Ӄ`}Om�GM(�n��.�lhFe��W�O	�|���BzۤE��fvv�t'9D+']��ժ[ު�뙟�i�E��/͡�������I�_{����B?�����;b%�5�ug��PB�\s�M������	��$�E�Y����C�HH��u�Z�3�G���'�����R̍@�>��ԛ��hٰ�t�n��f�����6å�To���زǦ��p�趾=!YrчU��s�PY���i��Ebo�bl�t}Nu�6���W�c�So�,k�O:r�ܮ}��_p��涧�2G$�Gi(�z�b�ۯY
:�n���!�}M,
|�k��g��ر����ᱞ9	�qt~�$u�0�v�`���D� �T�%��ː��w�G�,8Hqe).�{�J:��������±Q�υ&}d��p���i�W���A?ƶD�xUgE8����ۧ`�0��2Ex��x��K�I{`�h�P�	���6@DȢ��-ˠw�	���ŤV����*���>K�΅��0�;+�.EB�N5�<�UAKӈ������w}L�~����IN[(Q��6���Z �#�4���w�F��������X`�iL���K:f�4�eȷ���u>�[�3�^�q���W#H�4�o�^~F\P��5���+�C>���*'�̛�M�^o��#��u�L���;r{,^�������㌂a�[��M0b�_�!����?H�Ō3��N��L����F�n[����Z2��ڑ-�zj�]&ßK;��1ˌ��/ }�^��˂���ɕz%������d���ݞW}Sd�˕tk8D�d�\\���o�e$|�>�}D�wQ�m�*`M���&%��j �-�3"�S9Ka��LN��v�ɩɞ��Ob}�^&����.���5Ch�v�g��J/����\��� L`?BFB�^5|)(N�,0���&y��ԸH�<��_��u�eW�{Κ����|����h&$D/[��+xE��Rj7���Ok$��3�,���ƫD<"W�_j�ef�%q��H8 jO�x��!2�B+Fi��o�)a�n(�.�w�53�n�fW˵�{����VT���U��@牱���[sI��C��v~�lB�� �^�=��QV[��#�.����4�a��˝�li0\��e#�[=T����7n�X�읻EΨ��������r�Ʊ�h���Xrx@��Ѓ�;��&uk�1�V��p�[�F�0���`m��F�0#�3��$�<��*;��߶1�tV{f��Y@���n$��"w���毠)jy����)��y��f�tD�R8��u�J�^��?2!������"�����T�q����{���j���kQ�@|(d�@�B"��z���f1���C��s#9	���Ds����S�f�〼�����U���f���T>uj�q+~r�iduJڬ��X��%�x�\ �YXhf�W(Y�;�nr�p(fl��1H�5��\&{ب�dP�<����)5��f�yx��R#�<�c̝[Q#l��Ll٘g���T�tZQ.��1�W�W�;�S���W��i�e|J��"�m���]���^]�[���c)��^%7�H�N�L�EA��#Ĺ�0'�X_������WFﮭ�UE���)�D���4׌������M犕�g3Mh�n���}����� 8�z�$嗢Yw�C8��{���'�:\��٥Cֹ���O��/]�,�&�k����/텗Q�@h5ܚu��z8�=��۶i��u��Q��+��_���e��a�*䨋k��9*��DV� ES�� ��u~n���5�49Z�y %��_:_46��w"\'1c��YI�Y��QR�Z��EGr���tT��B��@����o���P��Qg)��cx6�i���ة*�Igw���.c?�����.�,�>��yȐ�k�۰��^�#+����HyQ�L��^6���p�rpd��R�^��͊u7ߐ���=Rt.X	�=����@���&�Ĭ��L8Z�-��9���`C�b�>�2`
��k�x�#��ՄQ2�R��:-~�6�?*�6�5��M�(Z�6ӌ�ϸd0b�͊��c$����+����: kb�
k���Z��@A�֘J��4ѧ�(��j��*"�'�f�*<��\ڝ!3�S�f�Ԯk�2@;�u���R)p�3�m#����\��A�E\��`��NчjL4���m�'2���c�̈́�*�@�*�\W�D��bf��#��l�Ux�F�y���{��0w@	R4�A��q� ������)!�d槭!�ۖ�Da�''S�;L�|��նx�ǉ8������j�0<ieH�.:����f31��z��U��B��[��EX� N �Ǳ����v���M�����gE�4�Ige������#W8z������Yy
�^@ő6#�	ߋZb��ŕc$�`ǯ�XM�klw���o0�ڒ��NJ�^�����n{���sjڔDh�V�B̲�t��q4�����0�C���f�;~�W�KOÝ�� ;�F�Nsv���R-_�OL�y_�X��)�V�z�ȳ���ޝ2��Kb�>��>U3�e��|HK�#���P�U��ڥ�Qz��0!C��5����%D"���e@,C��@$�k!m����G�~�b��������n2�p(��cHZ}��!TZ�`ބ>w����D�*_�4���(�\_�@�B��w���by{pǾ�4�&%��O�C?������Z������ .�����t'8��D�vx^
����~��"^د�gi.'nP;�q�/VJn_z�nvV��[T~k->Hg�����-��l��$��}�#$�V���Sõ�,�n>U��"�n�;���:�]����Xp�=f1��=9c��~hsxt���͑��(G.F���:�� 3c	e���
}O�	�5��G>����o����$�U5��Z���ܣxa��	ˤ�d�����v3bgD���z�����&�E����z��c-mr�0��Q��sع��Sz:�Hӱ1sv�~:��_�j�t�=G��P��q0eGA�~��Nu]c:B�D�H\�(S�bhHE�>} �eէ�H���$�ǰ�T���63 H`��ڶG�lK�T��+;U��[�}��x|�N^`[uo	�O�ք����V�k�+@��E2� +����#X\@㙺w�`��v�?)��6T �ۣ>�7�ѥ�M?oW������G��1tS�^�hB��A��u��+�
y��,���3�����r�sx��_年s�2�
�=�����[
;�ZI�|x��8gvE����N�%���v��٠��0�AG�Dj�<;|[�$�M���J]�{[z2B�}��c�	�h�gf�MϺF\�/��%���u��y���i���C�bE�W��
ٻ��"A����}��@�����+�+e��:{C�}RS~e�.z����D�Jdb�(W~�^��u@���������#�4� I��@�$�b���T���qT_�mڶ�>7�˥��*Gd�( ��"�y0%�tU��V;��	�d�^��e�J���V'W�HВAFbêY��3�EfFUv��vĖ�۳��^؉a�P���D�r��P��&u5���ʧ}R=�j�q�Ϝ��K=�U���?�~B3k>���W��vp����z@�Τ�Þ=//ͱ�/�G��H���_ml!��Mv��B�{�[�h���r���3 ��s,���p>�i���(E���q)���i�����IFx��1����1cGs<�2kDJ�o�϶"%X3�0n&��K�Σ�3�u���<�K�m����[�5�QbIwLӨl�I[��H�h/��]����N&@����oH�1m�.b�6#�.[fxr3��I�o^������?��H>�^D ���Nof��2���ɿ��Wy��Wp��G%�P�e�M*(R	v\BS��)�Րo䑮}�G�^��k�?c�ɿ���H�4��Z�����l�D'INc칒0�c)�T�1��������*ݘ�����ʝ�
��qVJ֋ UfTE���`~�CF�
��_+UJ�2}*�ϻ��$�#�э]��3��<T��}�'K���}O���߹��3>�@C�Վ_;�dd�#h��gw�w��S�/�T@p�[Ȍ�����pKt�QiX\����:[��Ϻ�3�w��*'�#��X�놥@��EQ[~t��=Sq���lݍ˲�$_Y�A#ȇ��1"�D:�P���AoG9���ru�
V���L�:ɲ���u��Ǜ�f�ӍOӄ���ތ.�M�ܫ�Z���=��3�:M����~/��È�^�P�+Lo���U'��tP/�y�Z�=d]w�7	���|3��M@YU!��>�ƎܯlH\u{�[o�6�t~�k1;��� AJz^ҷ�~�ݿ:$��Y	F���t�����/����|]-��h4�]�p�4�pL�y���G�! �0�8)��'�@-��J:�������͑ �?g�ft����x ���H�~u X�����!�����C�_�@?ׁS����v�3o�9{4�#���+8���5k9��u�S9�X����~S�D/F������)�2���Qzec[�yG	�K���s��o���h4�$�ej`��h�(�Z/���f��f�Uä�,	3��w�l���ܺ�*��2�X���r��V�&�Q���ȕ�ݍf����6�����?���$�ws�� 7R���g��nˎM�Y���G�Ǘ��Z-�Z��e/�Qi�p�BT;�P�P�jj`��2�A�^�ox�$�k�t��%���wį��Xq/ >��.���RL�&UGG�F�{C����\g�p��>y����8It�T<�x^�i2��r �2��e��t�3�\B�}4�BS���,�@HlUH�wq������	lQ�x��s�_�t�n��3�5]jvG��6���P�����0҇BS��4;LQ�>d;7!ޜ<��k7TO�G{e���F��ς�X��w 9،�������j�%��Ф��Q±�5dh��x*��ߙh���h�va�^ا%����������>�������h��
�h�F�����c$g����NɊ�BFQ=�-)��8Y[�A+)��IГ5ä5g�,ȏ
^t����y�O���,�YG�k�����z�]Vz�J�)�vf��hc�Ψ�BF)�|��rW��D�&D���p@�L>��{�T�ɮ�J�3S��bެ�����{4�g��(F��2�)�s$�.���3<�9&����w��Kq�ߘ��1L$�i5WQ�
{pA*/�6ڀ��]�7�{n��ļ�bh��I��7gf���w���+" �Z̊�Ε�!��|�8�_a��հ�^�Q�d}�E���,����A!�k�0@fg�
\�Ё>C�դ 4e�ޗ7���|���y�*aeCY�T�P��H�T��8A�YS��|_9ã��	�L=ȳ����K)nո�{�����g�D�H<3K��gNх��D]Ԥ�wp���$�"�����̨�v���"2_�4a���������oA̙�����[�fAP��KƎЁ�$�#�?�9��ށ>&\���h�yY"~P�}m}��͡�ߐ=UJ�,AYTr+� 7K�?oLXZ!8��v0�ˎ�>�l��-�o�@ȡJ"{~���/l��3�.ޭ;HI�f��u�u��*���ң���_7Wh�,&�7$j��ŎaZ�����,E=��2l�M��`�_g�q�10a��[F���߹�J�������~��QU���෴�J���� �!��J�c�j� i� ��v�4����+�[��Tn�򟴱P1JlX���B���%
����C���4����18$mx��$b�I�xP_������S�ɫ�d/U��:�t�?K�\�O�_U#I74'�:`�3#��q�!�g�����ɂW�z��%d5������ �
��^�Bz�Σ��`�xD2BZF����BPkm27��aF3tq$�Ij�� 6�6'���e6�"���hP���S�x���庋�N!���y闸�ݜM���2N��d�o%���i�jP|����ލ�:ۧ��\���\��J���[��ԏg�sD���Mh��V�;����2�/�)r�G���b�D!VL�\g^1����]J����g�P]� ���]����op�Cή)F��m	q�E��� ���-L��[b���n���?�����[�Ѐ�
g��>�!�<��4��(���J�oMX ��o�.���=�(���G@x�z�+ɛƆL'�H��f�F�-�� g}i�64�tB`ϰ�3��Pȿ�i��s2i��a���Ј��2>��V�,}b�qI�\=W�Qg(+��r��Q~H��(5mb!��Bno�Գ�>���� q^�؃D�Q�AM�Z��%bB�^	��=&w�ۅ��Ƌ�/֥��;%�$w��"��ӪI��Sl���3H��}sdǴ�o��H��`�������`����nG?�Tw�;�Y���̛.@�}�DZt�R+z
�kn��*���T�����x&��Љ8�O��L|]>��n�Ү�ey��1������ku��ƃ��,���lj�Ԭ.�A�T�����)~���&�G뇬0��@91b�J�wJ׸�DXQ�\�:�Tt�g����-���r}�A���v�W���>Dp~I$�#�|�dBIG��K)G���S�[�WGz(�P�*\�iK���@�(�]m�[~���ڷ5����A��RA�A��hH=�ɷ�V�mRÊ��Yڐ��HA�p��Q�VtqIv_��)j\�[Z��*qG2r;�B��qV���
��4�[���u��)']�Ƭ?)5W�/���)�<�a֢��%��0��4Q�j.���>�
�e�;�W��G�k	�u�*HD��]��/��A��G&Ex�O�wg!�U���7�2Eo�l�:�Klh�k?�K��&���5�)��$ү��$�,���XUOBzho��"�Q~�~�Q�w$W콫�m�9�X�qm�U �4�^,W�SU-�?cg��&��D�g:�%����@��S^5a�Lw�������Z���L��]k�X�ޞ*|��τ�`0i�8�
���#�~��
C��j�i��M�ٲ�4���l�0
�WiMa֚�ʄ�[^}m��p6=���Ȕ�>y���>���
��z�
���2�f�.;���3_�Aܨެ����%�j�G?R�ǧ�W��ɃB�9?tE�}�ba�B|6�!��Az���A $7h�6�i��J�k(��:b>7�BBX�)�FB�I�7�M<�uУ������qg[�?�[g�F�]��)���.�,�|�ʰ�/�"�?_''2�����$K���?����I������j�c����)��[��*�9����<�$�#�i�>��w�����!���ѫw�d{��.T�;ۺ@��-o� W�ܰ&�n��l�OB;�e!_x�Y�x^�/ӆF��E�c�1;ԃ�#4 �����Epi	X�T� ���N�$��=e�i�z��� ��1�:�䪫��2U����D�#d�p�5�`k�8��шt�Q>=��~�d��ځ��!˪V}�<5(���W���J9X��g"]�aR�Et�#���MO~<0A�"LıU$�d�\�(R�.Xqc��g���Cr���V'���1��"'q�wSl@�7�j�F����c���@�E�"�% ��$�8�-#���p�alC�l�`���둇�&g���u�eQ�?z_� �q!���@��`Q4��@� )���M�����WG^�Z?T�
IOc�nu�W�G���_�5��[���T$m��l��-̟��e����˲��Ό��9y�{����^��%%7|��G��N,b<hK�^J�)żx�uN��!u�)���M(똗v���0���j@��Z�0S,��Bq�nG@Gkt`��/W`$����CAO�Z`�_�5���Q\mq9�\�<�֞aU��j�htbnF��:�+S�z%���@mPN(��睳��rtC�0RV�*�M�>.\��&��`��{��MQ�el�q��lh=���'�����&cH�s�f�/�|D����W��m�ٴ��X�����宓b@
l*�f3�F��/�oY�@�m�B����<aX@"�m�O}�h|�>;�JMޤȾH���e����\����?��tw^�K�y��E'�|����ή��lW��DǝZ�h�]Wo�vƧU��z���d�
5o3=e�gR�Ӷ]�9#�v�dAbQ�|G��)�|N��z9o������o�2��\��3Y��|f��7;A-��;%�k��̖�C��|j\�r��8{�X�1=ӷ�B3�C^n��Y8_H����*ӿFS|�<~Nz���&�_L��~�ƕX�Z+��9�cʪ=*��h�c�J�ڕ��gs����\_\�4��e~r��������oX>���:ntG�6�@Ġ��(�v��c�������l�W%�x�*��d�4���=!�y�	���Нryɠ���d4�2�/��?(��*,lv���W��\��G>σ����+j*7Sޔ`��bfw㒸hk��+��+$?�����[���٭_��\.��JbʬS����ſ�}k�­��IP�8�R0D3	��ȓ��ܞ֣� ct%�x�ua���פks:>C���j����-+" �r
�u5�(��fs���XAT>�hO��G�ƚG�����
k��7H-;������_R15���Y������b�4�mߏ�s������O���b1�^>Z�\����X_"C��l��&���6���a�n�����e:��R��h�dUT<�5���ZN��(�B(�P�TAP��׃/�W0
Rx�Qc* ��]#��,�A�,e%��S��Y�6���x����U�3�v������-�@��u] τ��ӥ/Prm�b�w�ٹW��n=�yq�Z��h�}�a�G�@G
c�=��cAu�`[��Q]i��
3� Ӧ�D TA�GIX%^�\4�>ޣ6 ���>�[��G��U��$�{�4��bd��&͉�3���ƛ��d�HSZ�TjS����A����1C�J�EM���od`�/��zڄq�8�-ls��E_��0
�l[�6�WKK����bk��s���Q�S�q"�����y'��̣H֑&=8	�S�.:�E�ʰY�~T�|�;bO����~�l��EЊ?(l��b�C�iY�5�p��[-8�K�0�$�Ξ0�Dr��G�W��pF<��pW�JO"��V�3L��p ]&���lGzh�2����z��ݗxF�:�h���r��>&�N��5�C�M�7;�y|A���EG������aKt׭�	Tn���)��=�;d��Z��Dr�i�sG����rm_X�-��5��q���BkΏY@y>�+_!�������{�3�7�ֹ�^`�w=R�������2;׸g�c�g��s�D6�B��Y��g��~S�jE�-'��Zu��{�E�h�7�)9V(�U�R���Z��K�B���$��.�Esn}��Qx��b�78W)˝�S�^QQl���6��M�my^d��F	Mt��Ѥ���Zg�V[�1�t�-�*� ����CD:O�`[F�����3�e��o�fʮ+;��!h�RC���<ԩ�r,/���axZ���q�j�A�/�΂:�5���'qdiG���kpڷk(ǈB�:�|e����T�;������M�?r1
-O1\���3��"�!�a�iY����
<�	
���U�;f�q^(��0��uz$n�Y�P��#�d��y��nI�x����zw���7x+��4�a��UL�Hǔ�G���B�'NY��{?'ǅ�瑇z��P����ctS�/@�&tvUE|)q�����(�i�-�\OT����%�Kq�1��z��ר�]Ds�a4��vk��>��
Z��<S
@֘�������T�^ y '��e��>��({6nSPr����Z^���v�b�A�C�.IQG���~�5"U�}6iƫ���좧��z\�>�B*����,�}�c��9�>K�'��,��Ͳ�)�Ve�OpT%)�M��������۫a���S���}���!�v������9�t����V��P��-��2���
d�P����!>Q��@�X���iD����������z��D�x�U`���rLhbY�j/�W^U���	\5��-�#(�H�8��q�g !\�@���[�#m7�+��:7�� ��ǆE��u�3vҸd7wxW$���ů:���� �����J5��g�[|u�h�c��
�2�N_+�@Q�����S�SZ|�Z��L�&ldxj? $�$��7<�X�H.��f�'�����h����Q�"L���7ʀY]�9��������"�Ό��)�H���ɘF�V��_]�'�K��%��W��W���0ڔ��b�=dEYD�(��i�=DٞT�_B��~l�k�i,���.H#�5�n	p�#����W�?��llh�~������JD.Ӈ%�L����; �]gǟf���mH�g�������$
�a�h����*d�U��Gp�`��[��\TT�9ű�A�)�^�C
���;0�o�ձpu��L����г��Vy��z�g�㜤N��&W�/Q\��˔ϻt�#	Ѫ� �Hwe>����r)%�	�Ry&V��8Z 5���U���I�9g)V�������T3t�V�-��`)����R�g~L������j��Ϋ�A�#"�7u���z�;����͈ٜ?��}w�@������5�'2m���v`����2"a�w�� ݟ��(F�$r�f���,j���&�����Ʊ-�����5Y�L�$D���!�VEi��� �a�2���<\`mEX{�e���x�$��QJ]��-�򈌺�vD~�輍��_F������A���\�-]�S��@�K|S?bH^/G4�.�K
a��6���0�X��OJ>�F9��B֕.�>r�x��!e�!@U�ĕ^�����-+)��**�8�N��8��ET�{@��=y�����-Ѿ2��i%�+��c,�Ȟ�)v�N�xS{u�.Vs�;�h�6�J#a�Q�`֕�@�EE'�r+�7�$i�/��!����
)=RP�ԎP+l$:�Yh�w��z��Ҟ3���0����h�i��Å��)�-uK��>Ӝ�𨇵�PG��\��ޗ4!-)+p�?H ��޷,2rTD̕!�;�(n�a!"��Zy�yO6�����OML �� ��-���7�d��-�؝�~���Q�^I��Y��MШ�/�h%[MȐdKQ��!M���(	&���Ll��e��.C�ͪqX�Gȵ"�]HK��>��=Y�w=�4웞����o��#*p)�B�X�:h��`H9���h�ުۺ��-�[�ܯ�f�C͝���@ނ�| �꣰(���-�w)��1��Tvn�
�����.w�!������z*�Ţ�h	���{C�4�������EZ\���H[%9�-5��`����
��}��g�_?�3�4�Li�[����o��k��N	�O^�w��w�"��ɩ�E+	�K"ˊ��-3G�թ��eOv��R+0�l�8��g��蝐 _�_W�!@��~�������z��%���qy��Q�����r?*!+�A�����M�E�G�z��C����䮏�S׮?�}��R��вSz�G�D��ɤ^����C�^�0����XVG�c�/tc�x�钆����Y��l���1�3�}��K�۩>� ��v�IGrc閁]m�ԐD����Y��`w��KL۔-��5@J�'�o�����8���WʍȂ�
&�����@o�O~]�_
C�l�7�͙���Δ�G�m�%��P�,Rk; ��?�Ћ�0�w��ĺ��@̪�!�pP�jR2�  =t�΋��	B�@�.i=����55�U��S�����~6��h�r����3a��a\g�}���U��4@�{Ӡ}�NB���2���{P�����'��Rf'��(��m~X�`��	����(��jF�"�E�sW�?`��+�T�!��i.'��^�̐Ve�}I�E�͘���6���ݏ������U޵6�
�jA��7��g�ۙ	&l���."��ec��v	�������9UJ���k��4�y�i*zmlH0�����r76�����,�;ͷ�W�r��Wf\3n�'-.K�s�O��qi%�}
�~�����`(�&W��S��jg����NCN�N!5?�����_H-f��u~��Nٿ���<C-O�C����8R[��:8�`�s�Yd�F}�׼�>x��M�q��Ihț�_k�H
��0�ڍl_�V��Þ�r����RG
����w6`I3���Ȯc�/C8xf�*�9����Ir�Z��^o��m��U	������T�%[�Ew��W�
��C�Ck5�����n�w��'@�mv������Θ����ػfu�n��<hvn����� ��oQt��8��v�7��f�A����\���E�::?l��Y����F�Sɠ��������6��FlRܙKу���H j��tS��G1��7���`����Nb����wP�V91�7�)�k�J�ړ�t�YI\�c'�]�����=�f�!����yB<A��R.p�9��081̭����PsM"w��O���G=<����}@98w~��b@�2�d$u�o&��wP&�x/B=$=@(��g&$��AA�<�����,:�h�a�
�4�� �dW�b=�]&��g_��T�D"�CY�ࠧu�k'����V��a�*N�O�f.�r䚩����K�"{uj*��<X��u�.?��*7юxl�%�r�Եi����;�\0\M��N�nA�j/�@;&\f5�O�{��d�ḻΦ����:��&�fDbأ�������^���}g�;��R7o�|ʂ����v���bXQ�,y��R<�ΰ�"�Ԥ"P�!m��2L-��!�S�C ��w �EN$y�95�
tV⃵'��}�T����.��S��K!p��5��*p	S�
�R�d/����h�3��&� �R��t���gU1'$ǆ}����h�/����źħ���K�@Q�]�nI|��i�7��Nw4�;����
i��-��z<!Zs�X;̘U��G�~���i��6�,�8���/��`�);��?Q�L�m
>˨���p���f��q)��"y��G�me�cQ�|*̫�07N��A�ḰħK���f5�G��Ё��|JIsUܲ�Zٓ&��C)s5@�=��o���١Oi��s�z�3#�Vy��m����b[�c ޵ 8N�^p`)�e��'�(���[�����t�0��ADj�+�ff<%����FI�1��2lU`)D���ζ������#�l �r�o�ʽ~�w�2(W�}�|��ε5��؃u9�ra��E����9M_QΞb�6,BoJs�b�n�2�jx4��� g�@�R�:KAn��Jb%m�fGj?x&�D!������%�keC���Qĺ:㕧.?a�?�	f �a�����X�������AF�˔f'������Z���}n�����F<��%��+y ��嶑T�>g���"�"rHX&c�Fc�ni��L>.6�'z�Xm�������NʨS>JX���{MmzD���0���o���%Y�Xn����͢.J��@'�gR�>��I�s m���Pͽ�Eϝo0�G4n~G�!̽��l�}��d�(Y-�ie���-FH��(PY7� ����%�ƭ���j�@�08*�,N݅D�����[��Z��n����'��U�Skx�e�We'#���$�>��@�f/Z���=rػ����RR�Cw���>��z���"��c��*��NQ���E�&���0����i��?�ի�.dރ�q�s���RUkd�;�:���Ҋ ��O�v��}-\�o�7c�[�i�'gH 
���W)�8���ad�vB��BSLv�N�/�MJK[��_RIL@���*�K��<�:��F���<s�*��y���B���$�HS�N+3B�'�ak�v$nKD%ܲ�C�G�'�$��,o;)���ɐ�T��q�zKV�pb1��aR�}�0Ŵ(�h(~YK?�2?�C��L>498�s[�=��� !��[$	������=�8��r_��j�����ԁ5���W�y�D�S�m⢔�Q�b�9���6�ӱ���AC�G�Vy���o�m:�f�fs��!��6ϔ�$[�^YL�*w$���k1��+敾 m�c�vh�6'\0�Ƞ2����#,���� 令�켾�S�-lt�K�oUv���f���D����D�����s�J�;��9x�S!IԘd�j��~~-��)B��vů��:��4�ڄ��1}кX4�Y`�ʬ����4�&y/��7���I�/;�vK��[=p/�������H5y�BI$�B����~��YR=/9��k{F���`KZ@U�DxmYs�;%�������藳�`�צ��n��`mX�8��%ѽ�f�6N�L$#(�<A���U�aF�t���#P���k��0��mN_��9�m³������{ӡ&&F�>U�T��pC"��p+.�2ep�N��Ig���Ge�ωP�[���<���9٠���A^��)&�T(nY�D��1B8ڵ�\.�^x,=���a�"���G0V���(�����yR��ظ������F&�����Y�K-No	�2mt!d��R��X�ʑ�J��E��]��Nj1~�3���=u
Rne1k�i@�����ݩ,��ę��A��=3c[f�=nWS(�
Kp��Y�=f�b����u��z,1.�m� �0�8���A�ӟp0�K��_	���\ ��.��L�GPp���� G�?��k�5N�� ��ɤBF��O�Cuױ�	�bK��X�OM��쪓v�v�=F�A1�z��W�+G$�����w�wj��7��Ɨ5�d1����G���	<�W��s�����h�5��`'�k�����4�����A�Lp��?�^,�.*���=��{���*��
jtS��x�d��K�bP���Ů[�fR�aL�y��s�j������&@���fp�>�b�[4�yƻ���F�}=z�C�$��X�T��We�1+�����&��s�����)>θh�ܛ��%2��J���6C���z%�R��0H4���l'}�����b2��q/Ռ M�@��@��MLLөH���0�)Y����Ѕ,��hY�zʌȜf��8�;�e�k���榜
W��k�yS����0�m���}��~Z���.��O7@�)XH��@�8vz�0j�S�V����2�K(�{xl�n���_��K��g�{8�_ `�o��@���H���3>�Y�_^��6��UD����ۜ�6��[
�ӣ��+�Λ{��ὅ�&΢���QM|m.��p�b��T=�!��#ձaJ��]
�+��%N��R��V|&l��ұg�u�P��Ƌː|;�������g�K�>WD�������8p�/�Nk$�wӈ47
��c�V+?F��Z̉s��rɿM~�[2� �(!?�6?R�ln辇�h4lE�`d2���h��7ʧ9I`����!����bM��'��F�w�x�H�93[���i�\��갽i�!\Q��(G�<�����#kډy�%.�n|�j�l�U���gc$�(WuQ.:6L(�mV������M�cs��&T�~�����9�6 �T0�O����G"(����I��%`������^*���mD�Ğ���G�k���؁0�4�'��\7��I������ �}�`xk�����ܕ�ͺh����ف+H��|W��/�����1T����G2����A��h8aM�{	��aV��瀼hE������U)�wP��û�Z��-��Y�%��	����J��J�y��P d��[��Ҋ#�8,:D�&�zA�f�KD8��������s1Q��Dc_�L1��e$Ѕs��(�5&��&�~�9���R{�7w?���>�^�M�V���\G+_�_�@��p}��+M�×Ka#��C��DM���� ���ΒH�y�����(ǘm�9z��g��S�8�P�|���U�^�p#6-uq�ﯢU:��Z�F�b������� c=7������T�6"Ǳ�3<�;ý��C�tgs�yG�cN��%���Q�?�%i��y���+�F������M���-�˪n��):4�HF��n]xxh�m*�*��~J�^lԣ��:~�YS�E�~� �?�<m��Z��%v	=�- ޅs*�]*'���<���f��R�15�Q���� �k~�~s����;�=�"��P�T�Ʋ[3X�>ţ{����5	�K�Cz��������^ݎ���Zzr|�TWE���u��Gk❽/�u�1�� pd�:ֹ�D�vȃ�f����J�%|]y���n̚�z��\ ��|E��{!�n*����$X��,�t�է7��/�9�ۓ��Wʛ��`�L%���~1�Zkޣ���J�^�N�u�-���Ʌ�`�F��
H��܍�V�ۄH���E~�$������u��ZJ-SPf�Ͷ�I�w6!1�?�|���/,�;��`����kd�쥕����8�p��8
f�:�~#E)����-�c�Ւ�X�-2ʍ^VA�&/а�U̩+�N����wB(�z�ǖ��S��#����Ka&��ț�;W�~�Ά�L�2!��NL�z>�(,F7.� �3Ћ�͏���*?8^���>'VQ��f�y�l@��1>Y��Z!�x�ke��v�}ܒ<��n��e(�l1�m�E2][�~�
W�9�py��+
&q���v��E�ou86M aa�<���˼t��p�S�P���:�J&��D��ؚ���V�C�U���vA*1���t�� p��ɇdj�s�\��*͙YAK��j/�Vbϊ"�4--0l�c:TÿU�J�5N~l_�؝b�l��W�uO0*%�J�qm��c��1W�T�ځ�_}�^T=!�可�����I"0��SN{��#�a����������F#ߒn�{��=tiJ�	���z�Ϧ�������.�:��l��B������i��Y�a������������j�C)��DIR�E�q�I���*M!F�Qs5;fF�efH�/�e� ��b,3��;��(Ǥp��H�ܱ��M�HWsn-�Y�#`RF���0�n��䌚��c�_�XK).i��|*�q�Y��@X.��{˜�Z�Z����-�&sh��t�IVM��`� q���k2�;�fw[��>��f*2|���j��y����ÌfKʼCep�m{�/�A!�@���Y6mf�Ai�S�&e8�3D���x��Vl&��ƚ�)�M�^Ux���m�m�VР"�N��k�+"B��Z��ۤ�3_���U��r���V����L|��ti��''����`G�L6�ϟv�j���SP�58�v2����,�\-��".(8ܓaE��D�D�_���.�,P����u�� ��5X)g�_RA��AXd��Û"�yl� ҿΡ��x|�l\-���!��4�>�^v�x{h�Oh��KN�Q����yPKQѲ�x�%�~?���{e�ƻ���j���D������8>�k���폵Νϐo���T�d�R�5¿�u~X��x_C��#�:k��G<}��-1;fA�U���'���$k�㪢-4�Se����o�b�g�KKu肴�/�g���R�����Bx�b%V�
�����!МEdӜ�_Q�5�XW)4������{_�a]�_<t���4�߮ػ�
희(�^�3QA��m}�rx��m;��_�#设�����-JYV �������i<�Uh��.���!�>�ɐժjK3_<��m�c�� �*�ZhɊ���
!�ى�K�z2�F���AkN�R�M�`?�Xx-�1^�C9�����CMn|q��%�J5 ����C��O;�(�Tr��F��Α���=�ğ�F�ot���`�:�6����U�HO�Nɶ #�X������*��p�G���7"���Fy�c�ș�� ���9�-�X���)��v��ՙ@��ѵeA����AE��A��jF,XF�4��A������"Vx|�L������+�
q������~��}����g�Vޖ��1L�{��*��a�}��c�}�3C2����E�Rs����?9�;��{S��_JDZUL|3�e��>F]n��pp��D�����뇱;�k�d���)��jY�Y��<C��U����i}(|Q$��1@c��p}=���#�oȊ��h��QlF�h��@�h��P�� ^�E\j��.3k���R���4\},�E���[����E:���W� ��P�������_�StH��s�����{����1�2����|pI#��.����.�lT�?�9���b��m-=��+��YE䑀�}vK{����=���h<��)́�p�5��l�Y0K@�9zޓ ���]���;��g{6��}�W�k��O�_�N�L:,���b�-CM	3�&�Ja��]�!�N�����<s� /.!t��_(]�2�z`�����>ڬBm�3ǟ���4�!�3�A���k��U�Nnm_�5��(.��Y0��o�C�u��Mn[m_�� ���&�՘U#`&���i�-ݖy��� x�2W�������p��*e=�������=������O�Y�P��P:��UuX�����٠�=(<;�}�~��EL\Bb��s��)�4��4+�����7G��g.?o�Kg�;�Y�J�n&����CƤ�q���1v �\���i��V�%��q�j*����Zz�p��2��)��o܅b+�&��H�hB�/��$�s2�S�|�jX�+2�{`+ꈇ�����������:��U��W�vgS�^2ŗt(r�lǃ5��8	��xV�O��ɅX��a�)w������G�|�KӼ�m�V��
Q�O+����:�̿�\�>\/[��X�ܦxSB�,�F��8��rP��{��$9�Ǫg���"�u��}�*�P���a���:K�ҽ�"�O^���[�.cs6���9m"DP߅�H��s'�b���w][6�	f�onY�{ �Ҵ���|�J�>�Hu�ú��1��M(oZ֋b���������ӧ��A��n�+���D����j�%OX����'a�
��E��IU���n�n�M�o�Z�g7S, CHke���$A���xk��)�oz"$������:U)7�V�H��|�����4�H�T�V	>��"�}�3��zz�×��'p�39>#���K����ݶ�~��3Λ�f����B;6��z�-G�wH��d��>^wwJ
TOv��s�-�=���t��[J��-J��0&}�?Mb��q�t������qY o1��?�VM��{W��|����,&6_�}�,�j�T]���.G6Ӈ-��&��QS[
���?�'�=;ѧGHg�	*����Љ�>�R�9���9��R�<�p��>n5C�F���f�3�PXul~�_�g���+qr:���/��J�4��6X7B;�3���t5{�� �X�M���K�8C��)U�"�hy��~+:�W��܅*�O6f)�u�����l|�ڽL��O��ث�?%��E��|�|�������O�)�����'�o ����b����f2���|�s��R�X�U���E���WK>��剶I��ݶ�쑱�{���:�>�v �IP��:���[����E���7��\��(��@����}�i�D��$;��V���T���&ߗZ��K!�M?@_u�쪄���i�z�(@�eT`dʗT^��\tt`ݥ��6@E�]�	ń�~����9�t�?3����f�~���¯����!H�h�f3�����2���$�m�F>�����vOd�}�Ph$�e�7�y���5 j���O�u,�����l��7T�2���S���8�Π��8�7��NN��D��2�V�eSL���c=Dζ�_e	/�M� a��l��׉v{VB!\S����E]�V��j�zq�(-���=�� eɁO�#	��g*T7��uQ�T���y��5.=�L�������D(F�kIjl��P���{O�q���vϼ޲1oe�j�~�Q��DtxA�\f.L�����FV��\zq|@�'D��mw��(~k�`�>g�n��"\7�{�����ʝ+4���$x�����Y$�Ȉ.�9��A�zR-���-���]`�)�6龒�@ڟ�o
hs ��˝6^�t	����;�e���~<���~�u}�X��t:�^�"��H:`�EPǄܜ:�*Y�K����QX�/��<Z����OH���a�NM�`[<)����m�(|�j�����"y����ݤ;.w� �f�\ʀHD��J�� eWY��l��+e�ֵ�P�V��	�vJ�;�L�H�[@�:�n����	k�e��U�)���8�]�2"��L�HdΝ� �
�������C��X2���0|����V������i݌0j~7����7b���4&�/	��GQjR��훐~h�]��4�L���_sf��D�n ����ȑ��"N �,EQ��;�M��B>7"< M�iv4��0��цQ3X�`��|��T6�.Q���,�.ߣ�=��qf�䠣�pX����LmK�|҈��4�l�ؒ�-`q�P�w���/^>fg�m_�5��Nw�&��;�h��m�y�qb��ߓ���gs�	*m��aRb���^��1-,Eq����Իw���Y�M��'��=������̚N)L8�����e�8k��m������l��V���M���q��eGB��;t�TQPj�'<��蹕�
z��Q�Ҍ��U��w:��TS������oٽ�v�9�{"��sB�q���si2��&�+�����-�z(.f�h�<�x�./[+����!aP�$�?�� /O��f�ǋ������mO&���7`p����1�Ǣ���������̪5m����$�c�v��-�[���u��p�/��ʌ25��ͯӂ���Oy79�E�`sXc���ԭ/S���ܦ#�����+�3�eGv�}�\�\�H;��}|�[�T���=���ux�R�/�-
�L��P�$<�5y�4āpܽ�x�6�
 �T��,k�z%Y�z��>�^1tl�
�8��ɧ�����y�e���փ������)hv��.R����kΉ����uE/��Yѽ�S�V��qE���y��R���ȣ����|-����H ���h����(��AtH8I�S���`÷5�VY�T�PT��LJ�|b�k͏��K��+�$���  �_����~�ª�O^I���i4*��^�5¤>�A	OUV���k>AQG���q%�K��r,�l%����Aނ��C�(�u���
�\@O��k2K���T9����7�?�D7+���}�e��\C�/91L���R0g\���Ð�&��W|��*Ƹ�v}{e6��ό$�o�QA*�uՄ�4�o4�dZ�{U�Ij����'�\�?̨�
[B�t҇�����Xi˲Ax��:N4R���9�x%��(�PqA��	_8L��F������P!l���>���B��J�Ұ li���f�b�M%o�B?C��eJ�;cy�T爏yC�����B��!�^���[��+H�C����P`eu,Ur����z�t
	�]��08���=���B���� �M"q�  �b�<������I��������k4s �Q����а7M�'�b�p��o�%8��`;Vcr�5�D���me�f��!�؆��r���w������i�1`����C1,�R:r>����ӄ��n��.�?��Z���q�H;���I��I{�xʎ�*覴ر[9��{b�9尷˹���`�W����l�ji\z�\�G���.f=Q�/S�$�v�P�&��IuN�ؒ�gYc�݆!��꽶���\mG��5��;Ǻ��1xM��Fu���c��e��B�~� f{���l�9Y���<ͭ؞m�3H�I�t3
-@@#�N�j�w����Y$�*'�u0��Iֱ��<��jx�+ى��.��>�nQKuڳ*�(��e]Y��T�1����Io�j��"��m0�ٿ��! \N�a�lo.��������d�� X���6�]��1c��2���7N��\If߅B{a
�7�fX�K���W\X0�C4��'��  ����Oغ��i�|����̎f�A�z0�#8�47^>];{�$ٚ�P�ˉ7�811B�m���Rq�	ɂ��=��M��#'��'&��E�쮉XȪ,�v�X���M_�{r�A#�X8��s��cH��KnT���oNxehT���ѳ���q{��2��7w8~�Q�6��/&{�K�H�s,{!�����y5BN'��Uq��l�1����N�uD�[�p$QV˿�l�d*��%�䐼=!�/���@U���1�lʃ�|UC���Jܓ ���X[�N��Q�-���pv����	smt�w���"��~ﯧ��Ū�d��T�`Ь_�i��N�*��/Y�����z�t���W9HWɪ�d�[9��9-������a�O´K�U��IЋZ�E���k�]!��uR�B��5䩖�}���jϾa�N��i|�}X��
i�ȫ��R�u�V���������S��fuq\��,�&��&hK��!�{�"�JH=q���3�Kz�g/Ue.��܅��2)H��*��.�D�0e��V����FrN���l��ŕ�[h|N�M�����rP ���Cێ
�
A�L��- �ӝ�m n���e#h3&�w�O�����P�
��#u��3����uy�2�(}I���~�0��=��!�*��CMǫ��y�.��F�/Y�E(soV+���[d���^Φ��z ���+�IZ�R����w�Z��|6/��Xɘ����e�k��r�y۩��$����
2�q��Q/ A��-?�dG���B2V>��S�`up�bo���C�A�i�˨̎���ǪE�S\�7��ۑ�����a�i�{����mP4b��n�C�0vHu�6��*��]/K^�[��/4c@�9�L^��g�g���G�!f�=��3;G0Xi?Q�hݥ�z��]��Nu��)y�~��1n�a�k2��eݪ�p"�b�*���� k����[����5�˛=g�HHe1a�U\˞륒��9n����zH��=� tے�4�d�z��nW�oCxV�֐:���s���M T���4�@zl( �'/��)+��E�����y~R���p�����5����~1br��;AE��K ~d��둻 #z���FPkxV���fV�2صz-(�6��kP���N����Pv�2M[n�lgN�vJY\"�X��^$U?3����|	�dv0�`sT+bV��O�x�J����dB{��+�7X�RP�K��2jY?|9��An�U�~U�4��EqNPG�E��{���Ƭ�,��"� �z`m�[� ړ'^9��I�4Y��_{*8
������4O���贼�D�t_�u�r$��VlV���b�����v9�ur~.`(��6M�?J~��O���{����}�j�ٸOd����TX�O��r�
�_���|�)�Xz�;?<�������ٝ.r�ys �Lj�(�h#YTh�K���鶫y��zQ�}�9��UD�T���uO�����s��{%<[��z{�	Hڄd��$3�"Sk���kF"�Vt�M�2�t��\[�k�\E�/T��C��ױ� �J4�4���#�y9	���4BU4���	�L�����w�8a�0�{��8�u��3:�M�!��Hn��[r�T6E�~os�V�ee�G��&)��e��:�O'�K�Î�;��a�}��͒��J�튆���+qh��m�e��U���K9KL��
o��xk�7�퉤R��l��7e��7cO�<1��@�e�p�v&#���L��ftr 2~j[ЛU@68~��Ѕ�����6G��6Ri��y_�����!�	 u|���_V�QhA��C���gW6�.3�(��k����b:�0x�y�y�ۡS;�9��GM���G����o�Ox�R�x�����J�{jR.��%��v'�۩��~�'HO<)����!'"۸QU�acu�J�vۖ7���Q�T����(��6�P	v���I�mh�A�$�L�ؖ~ ���X~ͦ�G���Ͻ��oO�i?���#���3'v��X��@��ߧ_gc�Nz�~9p�E0��ca�u��:���w�V��$9B�{��[&ݖߛWOʁ8����ע��դM�a�͛(c�5
ֈ�n�S�2�\�'�d�J�(��pK���)D��pֱHb��8�V�-d���©��1$�:!W��BA��a�-�_�6���F�[ʢ۟��W;@H�C'���P�LZ��|�{b�6��V��+e��L,Q�g���ʝ�z�$A�W����� ������^i����I,��h��UU}�\��M�3�K�k��\�*�R�{<���P�
Gc{aX�ƫ����d䗢-���x �}����E�o�3ݭ]�pM}�������5���Ԅ��^�W6���y�QP��p�[�/�S2�%e�j�����9�{��E4�����������F(�뛥���? >���ٝuR��i�Fz��e
���yt�7����,Fn.}O/�v!���q2�=Hݺ&7�(/��e�\�_A��]!���n=+̞�ǋ2�+!�Y�cT�n!:r9ì���2B0����;�k&�Bs�q��g�=�����]k&�5d�D�}VܱA���M<���
�Ħ�ܙ�hH
ӟP���y�dRd�$v9O,������!.�ݳ�㏨~�X:�ͩc���\�k��FA�˂}�������<�	�5����Q`!.#���N��dgr[�L}*�l.2S=�Q%3,`x���j�z~�u�6�O��s5�F��6�Ӵ��7����0+�XXzfs�V�t�0�D8��n�h�c�}��Ё��u��]ˮ5�]�(oH3���-��!ѭ�&��M����� I9Ɯ��A���DS��`i+�QlF��z��2�vQ��ja*�	�Q�pa�����& b�;�yp���5-��u��P#q>\�踁��^Tu%��74Jk�W>B6|AGuXET`�w��e1hg ��+��ZQ�?	h'[=J@�)�l"M�bޱ�6�٩9�;e&F_ͳ���=��u�_5����]�'QYx�8�1��\(E��utf�)�h<E`xp興�X+�2�&��^5΂����@��$���� �Q_��Iv�����[x������`�~���~ �'&��!�~3�� �
"@o�jIi7"%����#dTq��ol�Y���x� ӄ�@s*�N)���AwyC�g���1X��竕ٲe(�oL��݃:nM���7n�������#cEI���̹��7�F*��UpEi`����ZhA~�\X���R�$"'k��]��`o�R����&�8�bn �� $q��lg:��}Q�e�Ƞ��<A���0	��A��t��'���T"��}�~KDH�0&`��a� �Լ)��v4,��b1���+A�W�ި�u�|�����w�;b�@���M+y&y'C��r��n�!ZfS�kHT������4�m�3��ߴl����\G\�؍fe�P���ݮ��>���1ʛ�&��혥�\)�(�]�b �X� ����%x![�L"�K�j�<�DoC�2>u�}h]/*��S�~T�0��ʒ0�M�o���纯���sv���u��s�����_���A>�ڧ�)&<`X�����0'���ը�Ȧ��2@ۣo��5骸J�����|�T�[����>��������a3Q��F��|�C�֬/��
L��u���dKWɬ��S)�۠�nE}���� JC�Iv��H��R�H eI-�I}7�#�U��"���H.]����l�X1�m���Ɯ�#$���J�b�ZmQҥ� ��(���2�e]�&�~G(M�{��o��y�f�5o��8��q�U�5���:v�}����Fӟ����1b{:�A�aRi���,*�봰����r~���?����]�g�0?8�`�-�*�Ҫ��� �Gh�C���o�E�Q�^d6��^�#!�y���_�cTGmy�L�rS�M�ɢ�}��zۛ5�����&���)4����T���/�K �|f
�n�/z�,���!�y&S��TM�Mh��v���ڟ�L���|��e�}�PT\��ƥ2�6V��#�x�v}�,�e��ђ/���A��(���bӔ�pAm=�$K+OX��*���']��0/0:$ 2�.Ho�#�-A&M���������t��g�aV��Go�ُD*��K�����5����[��	��}��D�[K8���*�J�5��B�Q�΃޼o�y�Ip����]������`� ���q�/N��@8w�@��XjK�r�6>��Ho_����1�ZW�Gs��*���|�@���r�$b����g�t$�]��"π0A3N�.V6��L˙�")���f�{6�����d7���'��x.�q%|G��o�{��a��Ρ��3aUe\O��k��-�:��Kuq�����bk���F���4V�_�ɡ6N���m�F�׷�j1e��Y#q�@��z�ܓ</Cy��c֎�_�A�ȫpJ��+�<�B
�/�x)�� ���ř�� �`F��2D�ƈVd�����̀4J@��C����I��#(�����Q^���T�x��>�Mǒ��y���1{'�9��3S��"N, v�b,�鐀���"����`����V��&�ȉb39ir���b�#i��]� @�@�0����2�p�a���ʐ�A!v��y �H�@Y�Nv�ڠ;����>w*Cf�_i Z9�56�(�6����j��#��jwɤr�tK��5m�@HX/�	x�x�'�ﴣ	#���5+��'���֜O����??���7�qu�u�;����!r��%[-}P�7� DG���5�n>`�9�@�����"t���z՛�r����nk=��5�'s�˹�l�t<��|�WX!ƌO��!�i.���@؉Y��d�劃]�M���3Vn�զ��2�C���Ի�跬�K�xv{�j�������ۂ����:�^�k�JB��pi��_ꮼ�W�	_�.��L�3Aɨ���"[�4�
F�+ ��!�Փ�ю΂�E[����2���I�v�vħw�|�I=����ﻟ��oFm%I"<�����?V8�~�N�nr&eX�����؟7$ET���^��YИ�yCD02Z�'�5�����@z��=�u�*��zv����'x�E�����)K����F�h�������w�i@sf�z�v�j�"ߑ+Y���]��ń���$��ǭѧ��H6�R�T�9A��}ex�'X�I��/
�й�/���7m���)Pʨ/s[!�����"��^�ɺkv��uuP5�u��-R�%�����uʸ�aOui5�C垼�Q]5(��M@�o����RP�c��<6�����[aF����=y��OD%��{�d�1����k���ꨡ:��c���)/��y��̂�y�r�/��ǉ�ncF����Z�
\��p�Lc{�aґy����D#7�[O��_6���q;-4�3��!	J�!�~�L�c����U�TN/��	�Ζư�C���j):O�3�WfY.bi⎃�;�W���t| ���s
V�EP2�j�A�'�������h	<ù̩�
#��x�F�$0���V_&�c�^O�;� ��j41n N�, ��H�ÞD)k�*Besp�wOv����t��^L����ܻ��C5�:�7���l-�"lgTk��[f�_Q���Ail��g�z闹���\N�$}�ŕyǚ�Q���Y�!���܍'����Y3��ІO�^X�j�3��
%s1���o'x�8�G�g���J�B�-���k�v�D �fg�{+ �5��K�����gr��SMD� ϓ�`�q�u!�8�М�pb�ሤ���u�lI���`;�(�	�Z3X'ْ/��\�D�9A_i}�X"�b������Ż 2�uhj�3�V�,���"�e��\v�DB����U��O�y��hR��f!@�)��V����;��8��6��ib"'�
��)
zk�1[�F��R���bB�ys�Jby�>�����9R��3S�/�=��d��v~,��c,�Xx�0��c�@'f���$�z/bڥ$�B��R��G�d�����2����� Ai>���D 591�T�'&�:�`|��R�	�6<������$��ZF���6������
��b�;`Q�	���Ӳ�Y:G���*Nñ�yX�$CG]i�<T[#x����{�L5�E��NF�S>�������(;i��zme��"W�zI��#�:M�$o�F�[�}�9E��g a|�9�#�����=S��i��z�`h���B���% �(��N���R��=QfP��>٣ا�ryO�6��:
��Ph��Ӗ�_+�,U�g�|�w�'*���ӥǙ��d��_s?zzbo7p`�]�b��E�H�� ?D�\d3>��l�>K�Op��)��Y�nr�YJ��كj�r��.?UV��c/��ٿmo1��e��kD���[�S0�e�u�������>n�J닚�l)�R`��<v
a�|��4�l�p��%��C��N���!��$���#+�!L���:�\_|��Ֆ�HN���A]�H�C��0t���}U	N.�v���B�amgO�ހa,l�;Md1��l�N��"ў5�;0^��O�@���IU��;x�����܉���V�j��G���8g�����޲�
���kHD��\�,Ũ�$�X���[�����G��35�j1�q�W��� �r��P���-�	ΨPV���t֢��Є�S��8��v����lF��k��_��Y��#��Gg�:1�>�irw�Z��t�D�u��݈���!I���4��&&r����!/�b�s/^pT��]�N���d���ta����˄"�/��]���$S�L\T�=�w��QH���{����t�R��3�"uj�G@�z�r���}�Gj=mA��T�����SY�0t�δ�Ě�kG4�h����l����<�:����ѿD�r��k�G�f�J����Ry1R��+�YD ��l/�Ff?m����!�T]Δqҍ��2�ܥWG�c{���kѺ�/g��e׮w]T��<�}~)��@��k�B��Y��B���<8�6r��m5�e�ޙ�h�i�6/����f<�$�m��m��$��E���`v�"�.@/�W�C�����0ї�f�;#*_\B�E�Km�G��,N!]#k�pmiF��g^��F�#(!��j�GlG̡�	���k�R�����8��\c���nÝ$@�����������NT���P�ifhF��L���z�ecs%�`?Z���kkQk&x>�	��0eV"���)�PJ+�՘I�*��8
w���J��Io�g��>��?G�i�20iį�U>�����Їs%U��'}Y��3��+1ߔ��X���8��Y�/��bd��%hZ�D�F.�'��K��׏�%�S.@z)_��˔���<l�1y���`��Pr�r8�S��tde�q@��>f�+vϾa�
S��;=�m���������<^�-�!�r��Kn�k	���~��R?Ґ�T �vy=527	�r��!#����\�ASJe�1��]y^����I�h^�S�1j��ĸk��B%NG	Fَi7~(�iy��v����Z��XI����졊��d܋����L�� �S���M�vS��`a�4Gﻴ��	~���.���oI��2Q�|GZ�*��Rt:���w�������nk9K����Gkd��yd��#>x�nW]`�L�_B��4�e/�G�_��*z����h���'���M��&��˦��<�G��tL�_tj%"���`��%�ؙ'C���8��kg�k@� mZ9��W��#��##�( �Y�\P �FL���+�L�r���`�w��T����I���+c���)?�����r?���"\͸�w�Mk�itr�wbw1�n%�ș'��G���/�K3C�"�X�V����md� �5��E�FNٔgJg";��'	���`�*þ��Ls]{�N'0�O<�+(��W)��6а�#���e�i� �ri�=���&��PY`<�¹>��|"s���cGk,Y���.�ۏq��P]�a�s]6����PTuB֥���.q'����XZg����c��S�`��H>�O�B��S��`Ԛ�X�k;'���E<2|���=�7����`U�w�$�{]���0�0�`�5��ok�79��j���Z[f�`��yb�������Y[17)�ח�,Q�֥���S���i�X�ԉ�S���(#�~��%/��ʱ�5��@e�#�`�a!|5�5��;�8���=Z�<�ư����jT*��b1y�v2�;L&�J��Ӕ��4�AB4���������ۃ$���nN&Ki%��nB��4P��L$�+�������Y�p��@����������7CWo�r���X:DI��t��Hp�"��_ �5ǂ(���U=�7�e9��	�]v�/(9�ƈV�ܡ+���a�h\���@��i�ɍHe�"FRb@%��������p�ϼ|�S2���j�8f�߯�j�!�vÁWg��`�C�̟����d���6���������c������<j�)0s5\D�L�ibg3_)f�͕ڲ����d�Ep����1L�T�3M4ц1{H���~�EQN� �k������Y�BdwC1���f,��fm��I��m/'���`�r!�zz��_磷�L��2�Wh]M�kF�\8r�H�)��7=}{��3�`��L�Z)�l��7�>R�����`��*�˶�'�� *O�dŪi�$���&RdR��B垞2o�L<L�Z�"��p�Z���2�5�L+�H�5�~EO�1�j���Qh�O�L"&��y�Jޓ�����9���9�m��p�e0�Zdj|XX8ؿo�,���\���/b�?V۞��LQ��!��U��B��F#��V	�SLw\�E��(JW�C�ǧ�Qҽ���Q�m��H����b0�����2/����e�#Ы�Ҹu��0�x1���T���[.W�ؙwL��d2>�Z���l8U����f�9ަk�d����)U�� V�L�f��P��[I�?��_T�9��d����ڱ��+ø��>f�&���=ZJ%*x �d/��$E�-*�+Q%�4�=�n�6�6c�)�5L ��>��"�Yl�1Z&�k��Ε`�ȫ_�>J��� ��$=��U�v�y����Ǵ�����6cSo���~���ϋ�|(��n|�2Vt�A��� �i�Ψ�l�!ʱ����'��֔V4U$n�o��\?����YQ�ٙ��x9Z�J�3Hi�D�������|ᦧ|V�:{l>A��U0����Z��V��Q��n����;@3�#_0]E���R�'n�y2�P�&K����D�a�����vr�!��hօ	z'��6I�֩,�
������~��|�XA1hGGp��3&
��@39Q�8n�|oN��/+Ilm�w��yk��r�M���|I�-��V��7azـ��Dg�7����{�3��15`FdO�������|��0.�X}�8��A�2N �Z.��o4�(��X�����le�h���Z��,�U����B�e��z�i�� ໵��$^�_o�`���u�����cl:W	;�w 7�b��S�3�e%����8 ;�S�Q�ϙA�v�<�/�S���F<b(�����)�4�	�O�Y����KY�#~����b�G�b�G�k�A�Ro��áw�"3�S�DLp��ޢ�l��(,2G��zȏ�����v��&1�������'QJ|���v_��7�ɁR�h`�MgQZYt�+5��i��� ���;�V�&n�3��yzP����Q�4/��&)��gT�}Nڀ�����-Sc?z�:������s�G�h+���/�:K�U#�@d�3�>f� pȏ�loH&���v,��L���Sh!�O�3�q�ݏj�V�y/�G4����&���k��+w��=>h2�����[*7�< ��)]š� XʠU2�s��Z�/�B�;n�����Ѫ�!�\]{�cN��F��M�u/��3}Ju�������<��;��6#��*[�:/�c�wn_)���':��]���ն{Ǫ�ZMp�Q��ERJm`;ǃ�����b%����VV@�z���}~Z�fXl��Gy���a�/K�	p@�g��S@{���#Qm%X/4'l#�
�W��kau5i����j&_�x�8�-�<T5����X��%����C��e�9�sLX���{�``L̾�,�}񼪣�`�����/ФZ!����x2e8����P��*o����+�AtZF$�6NV�dsOg�t�,v�B�^�_��׃����QT���+8l�`܅Y4g���v��F,��+5%>l��#�깼��c^�^�'<����h�A>/<Zޥ,�ǁ����|Ai42�S8�v�GF{���hn�-�?\��nK���`�+�s1bg�m��1�&�6�f4X�0	Q�W��S�DY�[PČ���L��l���RY�$�Mٗ�Fu�ϕs��Kk���bg22jG�M����V�
K���EЧ�c����d�4�L�kN���w��gSV��� ���Ƞa������,g<?rh?\|�R��2:��~���H.Ws�F99�(H���9��4;b��m�&-���O��>`�_R��x?��-�,�i���� �5��Kx���!�&w/��D�$��E��OY��70�dB��E�,&�0���m�6�E�<:+�mG���lL$`�R�_:��i�	%4۪�>��ȣ$�=W~iF>�~��G�a�VXR����k� E���'Ǵ�d�=��)����z39�ܶyn�_��Ѵu����	���J)O������DD5�m�i�(<�"���/j�b��~���_!���CG=�����yN���s���!$־öŚ��i��_7���|G��ۤ ILS�Rsɸ#��B��a[�@�-b������S���;�����^T����[y��m���SE^{����2W���v��t�& /�!�W��r�D;��Li������V!u8
�ڑ&�Q��7�伸�l"�`�Yj�Z��Bs��I��lWC��?�8IR�S�$����,!\̠��۪
�����L^�M�.���뫲����x��f�hC�?�����ˬ������q�c�l�D��:W \dMi�]]�I��u"(;���3�F9�t�) 8�N|򨸡\KY�h�+D\��1*F'���[O�$O������-��:�E��6𦪐 .��=�7�^'~>t�������ZG4�&%�]4���*;��pH�^I	���gݡB�yȎ��Ȅk���:\=�T�v��Fb�R��(6WI�nR�?��Ѥ�-��gDL�@�M�t��i*�^fW^7��s6��Q�z���b'Ϲ��eץxW(��Jպ��Y�3iM/��kGJ�:\���|���l�8 9]���ʆ�<J�v��Մg��h���o�hI�����mq,��e��oב��bb�І��B�z�cD��H7;�8�Js��6��,s�������X,t���4|�u`�g��	�9�P�i�֡�� ��!�{�>���"�u���"6k]�C��O`-lT���UW�N�B�z|��He�bFK�SskBM�^1K���������"S>(�����A�C?�p���sT�l4��Ay������R剹x�h���5��w�[T�R(��2�9Z�.ҧ^0�(c�1���d΁��&�,����@+�p_����>����m�_����:�!7NV�m�t�&>�G[o�Z�a/���!�ɪ�.�\�)b<kM�@�e~�����꿛Uj���Mqz�u�I�XQ���G{��9��j
-S���sA�'�ȳ'��?]��ҋ1<�L�]g�f<�%�An��(e?0.���V��C�3��1����@)�.�1�[�aQR�s�<���4�c"c���E�gߟ�6�%�߂'�1/S#��6�D<bFo��Z�Gy�`u`����=7!GH]:��~�ds�Y��mʼ��:⩂�wX��e�I^ń����)����hǓ�(��h��ν(�R�&gS>���'����$V-%�H]�{�}�^J������2^bL���^�=2�eZr�E��hN15mNw����̄�p|C@UC�U@)5��dE�K��tr�׷q<�eȖ�d�����+�5���d��fq��I�jei��BC%�D���S�
�Q=u�����t�f�R�O,�$珏��%9*��Us�#٫�z��v��$*�,�L<Ÿ'�;��Ib��Ъw'���JRo����
�0�Fz���k�o�y�����qzO��B6��"�_3i#O�
@ �UV���˛b?��9���s��=Et�l�Q��WKcR�~	4.�c�
���sKkX�=_]a]yv	��%�u����5ӧ��*	�}k0)�����i���\�i�0�]dy:�w�|�<
���i���\V��0����y,N�G�:�&x��ρ�W�a��4v?���E3ѳ��kѝ�35���	��z�T�ʧq����
D��ɍ���5������Mp��þ�.�_�W��L�n�0\G�x�a��µ�%Fp�yj'S0H�<2SX]�J�s�W�xw�'l����=�61-o���Z&��Э�"� ��H2A��Uf����-��͞<I�B�c9��Qg�����+��.�`n�Rٚ!����W�S����K��Y��P���0g
��زI`�Z[�a�y��|g~���~����6QвgU�?�l��jC7��łn�C5���V*#�NH�)�ܳ��ܦ������("Lh��3�d�o��X�gu�[%�/L���BM�S��JL�g�bw*s�ҿ�tl�q�(�����N=���l����
�[�FQL���8=���Ծ'4h���@B,{�fH��:J�#�v�F{ە�SJ���V��,��J���)|%�#�֧�%�|ތ]�z�L�G�6�k]?��蓕����$rO�)��O��Z���؇ܒ�0�F���!�N��[�pLf�V!�c	�M��<��b*=_ ��.ϴd���\Rơ��K�DM��Ѝ�x�;��H缔S��:�v�KX���mv����^g�*���2��nb���jh�<0+���.����Cq�YT���y�^x�	�x��Nedde�߄DQ=�����-��,(�A02-�z���iȬ���?!$O�o�y=������<W��EX;73��uX�qQNH㞬����@�u����_�إ�y�:]'�#Y�=����
R��ѝ���LV,!�t �el^&�G��w�Dѷc� ;�FS'r�O4����N?����붛G����&%����Bd3O-LJucnD��֟�-|�DJ�]G>:�ӂ�~D�,#Ӟ
W%M��p���9��i�Λ���Y��e}Ť����g�M�/�`��!Ł�^�U�"��iw���ī�3�451���,,M�Q��������R 0+�.�2q�S�2����+��:���:>$�Ϊ���1N���2~�Ď������-�0�Jk(�'�Z���E�["Bŧ���IƷB��	G��p�?F*�T^�Z��(A�N�]�b�*Cy�1G{�⻮wb����UoΦڄzm52b�!��[�AW������ʧ����MK��7���ɟjXp0������D:6Y�bM�Rx�m	�����(���ƶ�+r�fb�Ą<��9�?soX��\ķ��!.Y�rs�W�9��j
v2l�Q���	�o�2I�gv��FQ+O9�V�-�:&KP�C/Xƶ���7?�
��N����q���v�Dw�i�k�W���ug5���~/�gTrB�J��� �C��('P	�a?�p(C����_ �1ڰ��K��'�V���Α�r����Úʄ�� ��t��z�#��P���a���ƒ�orɟ,U�T��/�7�4u�vy��Q��t�1���k�[�|]Р\��{�`󥒓�� �=:��L��9,���,�ז�Cg!�*i}}�&	��ʪC�k|�n�� ���;%&��.����T�0�!'F?X�>�x�+~W�/?��zI�����Zj�wm�!��q4Q6��\���h��dO[������.���������F��e���Y�A38��ۊ����Yڧ�g��Hy���O!9I�MB1z��V�_��J@a�|�sC���I����[��$�OtΒ�\G���ó9J+�t�M���������}���\=�y���Hc��,�y- �I�Z���%���'h$�VhJ��C�����$u�� �Rn��h�h��,��	˿'��������vwv��Yho����������5hP3�g⣋|̾d��t�5�m�]w.�8�7	���U����݆�s$Գc�B�z�Ә�|�eE���z:��L��zn�~a����� ��l	��Gm͙���e� 6���D2H�DW�2r�^�o������b�Ġrcm�(�P��YO����Ⱥ4>5�h�'��
k`�*�#���l):���T%*-=�(�S4�pR��?�uTv�`o3%��F5����Eyn��-@��\�w���&���rƴ��c���=����(��#S({���e��4�R��s�G�����q
p6s�ׁG���lK�˫�Ӊ����r�̨8�c�҄���3�{W:=�㝴�]US��No��)�]#߳����U�ӊ�2�B$%,�%kp�UU�+��5wemo�(��tцkJ���(�}N8ӆX���
�ڦ�4�pq����z�M��hKx�oM'��x!T��]W8�=u	��ey$��e���X��X2O�@u�'/�=�3]ʸ�S9ǘԮ���d�Mf_��2�E�1ISctx��N!�Ey(�I����QV��m?|Jc>:�˘}��Z��,F�����?��P��j�NoI�d��u��U
>��lQt�uw�k���q�t�x�sȴ΀�Ok�eHV�A��mr�&i�t��ݪ��;~!w\�k���.B&�q�mkF=(�MIM�~����6EZ���O16Æ:�ƨ� ,}4�Ƞ3��NU���r}բ J
�����`���M�l;!5 �tL�E�h�.|��V�kRې�����*�,�����K�-���*�j��6Ť��{Y5�~& 0���)��L`v�<A[D�f��F�q%�W5�ɸ,<�g�0��̨d�@k4�"���?o�j���g��|G�(M�)֏{g�As[�
��"6aA��eЂxr��ۋ`ȍ{/(R�s2�*���n��i��1%h���{����rn�]�e��_'Q�I�;@p��E�B��2w�+%��A31v����\�}D����ś�F�7��
h@Y���L4�{FNY��aoghw���My�wJp�����>4t�`Jv�O�ϖ��IeŢj��fB>U�5fC�J���=����oz
9�{l	4I�U�F6,c��:�$�폊&ܳ9T˧вKhW����l;�G���(�����P�j���"�w��6e�M��Ñ�K�_��Dj��/\(��w0/�W �6|�9&2��wΏ=�cjܑ}ytqQ)�5�ݱ��F�
Q����ϳ�	M�]p�0l��5�i3Ě�Y�qꞣ�P�/,bC���|��a��L�`��y��+��F�<79ܘa�W&El�1N���M�i��x�]S;�M{vH}+m�b4�?�BU��h��U�y?�*R��P�l���5
-<\����޻�����Y��;h��Z�=^Y��A_?:_ h�l��ǶSwF�/���"�E�?&�L���X:f�=G�Th��)�ᡀ.W��0� Sg	�.�O��U�����܌P��e}�'F�֘ź)8��R5l��Ac���"ZY��:�����p�j^ޤ�t^�u.��#��J������m�P�X��T$����<L�O���a��Wa�,����dg�OHYO7�M,\��>{%�B9qvfƘӈ9&�v�]�# V$���f@v!�I �bL�}�<��}��`4��v��3�P���MwE���?*<X���YB�<F�함ht0��]�J��H��;W2�=�NE��;�Qz:�q�]Ԅ�T�>KHL�*�4��6��"$7�c_�F�� �.[� ݾ¾/վ�	�;ڡq\�� j?f����OeI0V�� [/o̒����%d+�y��ǻ��Ә.'Q���&�\|�� Bn��r��uR�g�b��us=�'���P���2�$�A!�E�RN��A�{V�SB���,bfq����K�(H�\�drS'/��u����t�^&9m�j�x��(q{��SU����8��R�#e%��[<��oz�-*nb���v4�H4j�؍�Z�Y���A(�詅�ɀᜠ��,�('t�["i�������f�U0z��?�g���R�(ħ���A8���)�:�����8�F��"hYE*U��vy� ��IuOemQ�W�Ljl����9�(4��'9�տ�^�:�� /F����n�-�;SW0co)r.!�u��b����I;����
/!���b�
tq��l��v�3!5Mv�	@�~} ��_d�ֆ�C��5��0Ӧ� }N9^�b���9���\:�w����`�?`r��3��}//|�{�<u,�n]�[/�~�:Q�����'��s�>�ٗv�ɘN�@����9R�<�3�J��#1����m�a�G^�����Z^��?eRuT"�Q���	��
=1��A'[G�m��Ya�{�������O�X����y ������?`"5T?s_Wf4�R�^*��o*5��Ӌ�g0�e�l�!>>��o�C����bx�[�Y_KX��s��`'�/L��n�WK�n�z�1�Fg3���;o����+�+]�T�ۨ2O+�Xx�l�X���_�\�RMq�� ���a%G�hG����f�	_g�!�/v�)���H��[1�:����+}-��v���Z)��Q�PN�� ��#I�뇣����4u�~��f3K!j��I|x��7�n��n[=�3�h&�d�҂��Z�)�l2m�h/��P��%�i%ct�z��i���"s"�tB�Ű*ɛ���D�9o��W��:LF�`��^��M�Q������(:f�1A�p��?�)OQ��W��x��^+����Զ_#UZ�nw��lN!;����Tf���Id<�9趸�!�ϟK�r)��&%��Ku�%u6πq� $���Xn���P�	�Aca^O	��*oRSߠ���|�6����w���Џ5����5�:�#0�=�Fm�����^��_*����pE~�Ҭ	��2����F�8ő��H��:��{��s�S4@�(Vg���s�(�����ҭ�"����2&��JV:�C�����e*S�l�AD�@f�4qќm!��V�"�	L��U���OD��\��B\���]�2�V�do<�L���M;vU �odӎ�׬'J���9�W���q��;�6�'qn��z#?����m�Sm��׾r�w�Gß�wS���ZD+��L%y���	��C!�͎���E��k�窘+�������v%����n+�	�7�:H����.�o�vI�
S��e\��x��r�6*���$y����H��쇆���O�SBf��Қ,-z�C�/���7h����7�Н(NZ�)�}�H�u��3vJ[	�P���v��<�:4
����wuC]���=ƈ��	�ʗDY�g"���e|��������h"]yO��*k�Ԛ_8�WLq��'
�+��0zd�Յ�]ȳg�~S���"��.���5�C�K������S�8r�6/��C��ڹu�(8�`CV����Ye/������֞�}O('���%K�q��r
)�x��@8
2�(�6�<��b[�1��|Λ��#~)#��HO�;��h�U?���
��1g[�X�я��=r���e9�ď���n�]0U}�=E"�]t��T4	$���a0&�π�.���\S�/��/e*�d�?��09�����Ftjj����_��eL4r�Œ#Y�a
�h<i)�dZHk�9ɡB�N�
�eP�n��#v����x�sr�Q���#Ւ+K���E׏�t�(�$���ք/ӷ�L)Dj���o�f��s\��L��du�Pzc���M�<�+��~iL��I,����+^�L"���8s�1X�ھZ5�uO����!4��(�,M���v(�r=�XԾ?ro'�A�G�O�q�p�����}���!�KϺ^Vi>���}��|��绀=�]JU�[�ʎTΰ����j�rs���ϋ��� +���8��rұp��.V@K�WҲ�`N%�=6m?�e�9��#��+���	� ���y]���hZ<�EMy�p�Ҝ�ha
��(�EmY�}��ehY�Ce5��%:�[��J��V[_�~�X@��[��1P0�~}? }U>��:��5BϪAD��	��5�aJEW-Gw���<ѷ.q�g�֊T�&]��Ƙ�!��I�]sF���1�5^��PTH�)K�@�wU�A��&�c���-u�N+����	�n��Y�Q��	Rm`���"O���Ylx���#Ռ���Alťk �����Q��ZSʬ{@�F����<і�������u�S�]
B�AH�"����~��:�+��8��3����]Q��,JG��G�0fg��UI�k;o���OdDN���\A�3�����<^�2(��Τ�a��7++]N_j����t+)2�3��������kK�"v�,�Ԝ\l�Ca���Þ�&R������� �"��>�~�&7��v��m�'��[�r������J� �J)�zf��#wY �o,��А���7���A� ��Ă��J"@��ʍ�H���Q���q�S��$-�M�̩��	���]�i�&�5���D{lki���Ll:�@�2ZUK�a�k5K��{{
۫��XG�]	�L�����I��Z��~�D#�J��҆C<f�z��$@���"�]��Wg7����5+yZ�
�.nn��T��B(��K���o�,��	���>���lৼ���}t���J��
�ZUT��O �2U��Ͽ����:Od5b}��)<y�LU?d �ɁҳB���m�ݩ�58���!3c홼@[M�S��]�A$�X��q$�ű����6�>�=���)��������j�OC��#�����X�J�M��:M�X|��חR�BDi�2~L|^T*�eI�w�g�{�B�jg���(�ܗ�Mh�.�\�(��HIzӟ	+��`�J�I��
䠟/�p�Q���m�*w� \����ۍZj�E7�T�]Wu��"؆�������UB�r�]jX*-8ҩ��O�_��]%Wh���F����%2��ڶpW�)��?"Z�r���&�	��3���zŭ	5
�ܖ�M�Em��+�>�@��a��w�{|�9��K��:�y�_[uA+��j��G �ӕ3�h�1?�Xs����:ѽL''�R#�:��/�xk�8�ԣN�[��^G>�)N����t��$�U"��D����<췲��F�5~��'<�
��o���*A%��eVt1�/Hᨡ�/q���N�iG��J/�$�c8�r��O�a���Cp��l�������¶؍o8.�V�FXO��q�[���OV������K��W�=�ėX�������i�A.�����q��X����N;����Y�l���\x��������W��nI���Kb�i͈��Η���YEIc����ih����r��!�G���)g��p7�R��Nx2�k:�QFT����|!m�˫/�a.�$6�ej�)P�At4���{�{t�k�8yD�04�l^���i)���2���U�|}��ƃ@x����!�C	
+0���/���@k�]���GW�=�s%!EPew%�t����/8�WUc4�3"_��7���f&RU2A���N\���\%��[��3��F��U�
̚K2 �g�tkR��A���=�{��7i:凹p�yp��´��Rv��NҝJ9Z;���F�N_�&�{�����>��v�m�P�1�#�0�`�C*!�9�*�N��jA6JOn~A��~��4����SM���3~0�+	�����L�)��r���'*�;wc�`��N�JdCc��%�յ��z�ݓW�mBB7R���;IŊ��Jdq�u��ˍϞ� A�U g�l����4�_�nє�RX>����w�Q�s��Dl?U�ѷ� %�`�DBih�R��Q������P�'cG�vc��ݏ��U)r��;� z�)0���KiI��bO���7�?`$�����`��u`�e���Ň��D@P���ZG%��a�Y�i5_ioÊ��*�!���v��S*	�=_��m���l��i�x��HD�C>t�S��Z���e9��[$�̤��k���~��$!��72��W���������D�۟l+�Z�+�$@&۽=��nn�<�ͻ�_�����(��<&u�U���e_��u�LZ>F��z� w��H�̹�����>n&=l'�ޠ�K$��>hŴ�;$l���iփP�}�ī�x'���ۢ\�&Q���>������Ǜ��� �;�'����פp\�J�2���ϐ�~�PSQ[��������1���
�4�U5_���� .ǅ�>��L=���Ut`A�F���2��dc����+&��2��%�hv��2
6�4z�n��ؒ���	��1�$B�?R��g���z 4nP��[Y�ɛ1a���E�( �d�W�2A�[B�I��ӳL�:zM�͒�tai��.��ڶ]%������n�R���4%����̲NH�X�1�%��H�7�gF:�QC3�Pp�^7�AM�\�����m:�w?��|xy[h�8���%\@�4�.��ʻO/�o&��L��:�g��{^�f�T��9e�,�ҹ��>��2X "X2g ,W#��7�jh�̪��RG~����T
��+�+�.�(��]~-��,�G����ŞMZ�?E�b�����1*��#jK���2����A��`E����1�3�'�A��<��iK,څ�g��3��c���t-�e�S2U�2���d��DԌ��.��a�DT�s������N�k��Dc��;�5e�h*�K�o�]��k����̴,Jk��%6>��;�čϤ�(��!�3�ğ�1����:L���W#P�K=B�4P�E�@�3�,��hd����2�!�"�CYΡ�LI:||��q>e��,���M����
�nw����݌�ri�z����6�#;
�8(���Oz|�=��9Bk�I{�%!���a�Gش��+�!�_�	Z:dRZ !�ݑ�GӀD����M�R9�z�S���r�_��΄/t0�-�1*1&����X������qE�kd��P�1xj󇦇��Q�E���G1�z�S���i!,��3ۊH�f��8oI�h�=�x�����[�Ddə�m�;7��KW�4���� ��Rx��N{ɶ3�f*��v�!)j��=���N��!��+W�}�|��d��*��0_g"�B�\��������9�L�-8�4������wB��)�Q�� ���fr!��G�������u��y0o6\����)�C-�Uܶ�s�if~
F毾hQ��Vx�Žn�yϒ��Y<X�>�6Y�c
#{r�6@�����DIK�B�	�<r����2-��]��kYMǸ�r{���i�O*�ս���b������N�]"���m��6����-9��N�(D����U�ƛ1j�k+��Mќʄ_@���A�c�ZK �|"Aϗ	R��C�����46C�11.�>���ޜY�������r�9樣M/��/�د�k��d-�>��3P��ճc�%Il��/�<��+V �7���CP�2 �u1l�ݷ�~&׫*ن�p�7��4�ښni���5ǸQ�.O��B:���g��=?�,��j�r�"S06`D���O�#�Z��#S	²�R���(�ڔ$dpW/�{���Q��KS�L���ϙ��+7QL�ȕ�S%M+n=E7��f�le����P�u�#_�]PU��s�@�I��'��D�Ѣ�j�(��׆��z��n�,\�E��K]�=Gi�D��<ʽ��R���9K"4T���ԭ^�Qݚ>�m�~Z�����%p�V6>�ٵ*`R�eQ�'l�;��mK���j�G��Z�6>L<6�H7��ٱm�W��G1�g�%&P(;��A��57�9|D����,Ĝ���g�ɷ�y�Mw�;;�g��R�f��Cb�\Cě���,C^�;�j�dǜd�L,;��O���\�5�'� G��@ض�a�+���2D��v� 䥃oհ�>ʄ$BL�m\�'�S6s��������\�^,�}*�y(��PO�YĄ�H>����g�r���fd�\�Um� ��i �z�H��'�Y�@��5Tb�������V�[mcq���`��T�h�[ǥ�g6�U��7�S�ڏ>� Fp����`�Ak!�ߟS�w]U��5�*Ixy�~v��"l�nJ��'��=AZ��#l��b�\/�	���D��炄VE�oZ/W�Y�VkpG4FI��|a�F�l;�ד=q�Z: G����C�����T�d���%Ijz�gw�3e�%�l�Xm�3Z���m+�hf���h.�P0b���ez\[�Lͮ�~J�� T�Ν?��0�d6%.��s�Dse$��r�R߻k��`Y��aW�OU�\�%�Y+��"�9iMB8�o�
\����rrjb���C������朵l?���DeO������@���mP��i�\���=�6��#1A[�F�������[�vo��m�?P7�Q��`yD�(�'�*����x�y��i.���8[Z�*/;q�-�4�w����ₘ߻r�3ET���ou
��we66!�� �х284�A:�1�[
���c���,��Ys�R���yk�4~��WbP]Z�x����΃��)������ګX�C��g�|K�i�Q�z�.�fG#�bh�����|֫=T�g?���lsގz*t�^�f0��L���r�&`��Lަv�끔A��t1�	˖�õ&���8AY�����x�a<Z0^�l����H%�m�S�f5Uz�\�Ow�ߔkM[{PSX�/ 7�r��
$L1J9XL]=tqV
z:�ڛ�&��ρPi���bm��pg�F�1=��LR��l�/�FfO�!*�L���9�v7��rC�ɹ�b[ c�9�|@kn�a�R�O�k�I��W��*�U6���#����Crq<�e�k@$��Doe<$����\Q�Iρ����ݾ�a-�{ur���#��8*�E����9�/'��_$0�a+;����d��8�aB1+WV� 5@A�f�m���"�0�ֽ7W�y�`�kْ���,oU��ӓ����[0�u��&�'�}�u�d-d6S���;�����e��!m�nZ���GG�}��Bʋ�����xm`�"}�6Ͼz�vm8=�js �Kp�@��T��1��]�����2�+~D8�����륌./��
>�Y���n��ݝD˲���6�6����p��=W!��+�9/va&�8�	V��-�a�N�se��9M~�F���j@d��e?2@[1&��-�F�S�~�!�-^S���ǓQ`���w#�5��K��g�Mr�RN��<�r!���o�|6D�=�雒�����}����l�\���lz�]��ܒS�X���P��}�o���_��ҝH�t���nX�U�Ӗ,��l32�`���y҄� �#E9�iqO�G�1����m{��|�Ƙг!��R�T˓1�J�Fs!���M�fdP�b�% L˦zL\�'��<��~ϡ�H֭[cY���D�d]H���UWh��Ԇ7�N�\�h�C'ȜK��o��aD]�R����+� N�;A���"��3�����������F0�d��*D������
�k�s0U:�3J
�T�6�4��5�3g��6F<�[صgL��ǿ~����,����d=c@��H)�@Yi!�	<�g|ƛ�������������м�:q?�E�F�+����~e3U�k�Fț�\�����	���n-s����m���~c����U>��������-����x�	���5Rt�$z�I�:9'f�'V�Z��D?��)Q��b�pC,}~�����_�%�;�Ŝ���c��Py�veLX\K��i���DJ��M]u&N !���h��(\���̸��mª�e����,�c�T^�6Q�g��5[p�g���%��^��������J�:���I)5-�B�Ծ���g����?8z��/�Raf�O���BRϴ��$Ol%��%Nh��z&�u)$�f����ob�;mQ�Nm�����+i{�_��2u2�^�~�cL�z�'����^xq�i����e�/NwC;Jsm�D�P��@v�P�W��Z�Q'n�MA��ꚏ�T��k2p���HB����ލ�;���hke��kIļx�g`��'|8p W����\���;���� ��bJֹtU��!'�]��B��ɔmb��d� /b+~��P�k�)d`74m�|��/���~�j��:�ޓ���Ì�+�� τl'�(nC^�f�p���~��~|!��snԧT� ��{$ʾ�3�@�����xO�f X&J�=��7�'�pb����"�}�`|@.N�
����d�H���L�a�ػ���qW�L�Tq}��ae*Taj����v��H�~�{]��(����hE���>& ���=��M/^�Nxm!�Hp�i��GO��!N��C�̘��)$��M�~~�����D��#��+�̉�"���+����+�(��{'���v�B�u� >�S��Xdd >�R�1�2���\Q7D�'��@'���d���s��s0��$'�����C�������PT�N��#Bs��Si�=ݘ:��耝^��Sb�Yd�%��ڒB��a)%������L�g�����:+���2Du�Lk���hL��^d�\�,X��֐`/�Sj��"W*J<�}l'�o(!3�=7-��g�C�G`Y�t���D�����DN5�2N��_��}�Q3'G�FՍ�Җlݷ�!��<�-�#[�H�	�X�y�#].��1`������'�]&���A�8U�����b�I&�{�!߭>J-�t����F���n���t�_�%*��׎�7�.eI��ۊh�����j�^�|PAI"V�!"���ɂ9��*��5�)s�ܣ�5��Z?X#*�daz���j�4�o���m��	y�h&�{	��#�>���X��V�2�Gi�=��Vi��8���0r��C�(�"�6�sJ�M�}q�Wq���Mc�@�s!X�I��mdTՉ]��\�ֽ�a��q�ج�5,gi��"H�'�?Q��O�e���V�Ɗ�L�J)ys��w5����G�5��k��5�IJib�at��I�����c�<�\���������H�y� .�a��Z~�S��a�����j���>��2�oS?���OB ��#~oKn�߅�dz��E��)����ϵrE�ʵ�~N��!^��a�W��(0�}� �|K=ᬥ�ӆh���?+�����_�t�+�]]�K�;K}�����	I�<9y�^C�N	l�����j�E"+ɰJ�qm�3�k]0�&O_�:0�f�&��B�"f�C�a��6�N<��R��ĔN��t�D���/��Y�p�i0`�I}Θ���+󧠪�YQ��%�d�L�q����S��F�i��W"���x�Y!9x/CI�	�� 	#�o/ڱ>��M�H�]P���n3(hoL�*�,�V������m/�/x�d)��  �٫wZ������[����<��Ϳ4 �5m������x�uZ���Ṳ��ǉ#�NW�j]���E���a~l��nc������'{*�pU�k~��=���=(BRIyG�Eb�f=l+� �Ͷ����c����w3K� ����̷	�I!_Q�ǧp�#���ڗ��*��c��"bf"u��K������Ѯ�+�˶M�ƟWF�R+��"�=!?Q�)���8�~l\>��O���l/����DY��y�����w.�t����p��Ë�1V��k�s�;�7�즶�K�܉���}#gg]ݞ��D��CL�0cϒߜ������J�mB���>��tҭs'g Z�&+E ���'�1w���b���������JQ�H'R����;w����b���D�^�/��$i�x���d%�}�u�Y]8�aK?�!�:Z[�P���%s�ƪ�0��� ��׋ǔzG�jWp���3�=��$��0u�/w�'�{�,�2l����ܨ�7��~@b"?�E�����-BG,8g� O�Q@Ϛ�j��n�@�@ʦ��zuaf�[N������ȤaY��d=��TrA?+���|X�b9�IE9l����Yʄ��_���CZ-���M��ۙ;��Z���#��I��0��Ү.rS��,h6�DD$�5V�����c�m"	�*N3F���A3��6�zlʚt��sV�Ch�T��KA�b��D����di<�r��b �\��������w�k8�<Lzl��>��^��r���v�ű�&�Ű��^�i��Y���?���O��L�)����N�?V��U�Gy��f���bS�
`W&�?��Z9���[��0��D���m�&��,6��b��{��vQ�]+{ �յT�7�ᖣ�,@X?D�����e�'�3�ʹ�XNgY2x�~#khxs*
��nB(�՜�m��P4�nS:}�E}�)�.Rз�\��U?�}ʤl�$x0Q�GZQ�����U^*3�|���K�\�����J�C�ϤO'!����gk+b��ǟ%�3��\����x ���}o���2[	�����G���N��x�'9ux��?'� ���1���t%�?_�#A��g����)���C�9b��߆ny��&3� zi�],��yr?eE��C��'��,X��r�������ih`ب|1��%?^�	��]G�ʥ>SՆ���ی���E$��m���0l<�b�H�4�%� �Iľ�!�>����[)�nZ�k�*l�� ��a��;�_�:�u����̤�[�O�O~p�|oImay:,���]��'6:�VuC�wT��b���
������W����y(���uS�n7�K����u�VcC�ly�OqКY��(��}�zZC^	�{�Ieg�^��R;	���K�H����a��x,"d��&۪_^��mT���(�5`RĽ���,XCf�A��xn�9��Z��H�
Ĉ��=��[��-���4�E����@��i#a<P��H������%ȬK�5_�=Mp�����2�|�?�!�E��(%ʅ�=s? S�0̜	�վ��t#5
��KA,�E��ݰ�9\$\������S��^����@�-��,#����jG{b�#͏X��1��O�j��,���χ �'[��jZ�`�ufF�f�-.D����]�E���ѡo��OW��f�E�Rƕ��%��>s��`8m�d�I���b��������Vudw�ME0_!������\�:j��KG�TpAӈ��
�]�8�n�[���ȝ�ϧ9}wIÝ9�<��Z��e���ǟMϚʵD�&�[��{�W�54�dV��w~����s���Co�P׳b�o��	�����ɤ|seY	MS~��g��,���p�~;|pv��M�;@�yEu�fs{ЭhK�JU�zE�H�h~��
�S��$U�ʢȓĢ$V����v��f��|��tP%Q�\�I3��T�������iF�G������U�TI�J��Ow�����\��\g��y瞬��ӿWqOM�&�WNq3v�ǟ�iu���a�����7��iЏL$CM�	'A����m��P�?�X,0�k��H�8[;�=[j���q/9�����h8ޖz��a�y�߷ө��Y�Xin��8X̮�A���UK>�iI.j�*Ԇ�&_�$���^}ͻ�ꊻfn��Uj��P|	���G��f��dP��vy-e�t��ʐ_,@ޛ����t��K޺D����C
�&5�����?��#u��"_Q��L�<���ٞ��:�K�>�&y����N3E%�$1����p�(XN		�u��.�w�bHv�|�u�F��|�ӯ.������E ��:�~��F2�$�(���|�;�V�%7�T� �A���h�(��u-ȫ#�I�DY���G�w�!��n"�{.�v#����q@k�
�I<p�5t��w$�/a>�L�r�����j�u�5���p���e�������BSl��o�
�R��͏��C	@���y��mcf�Isy�'1�Q�Gw�|��6��'�F�`�,
�K��N�&o�\ԓg�0
�ɪj4`��)��^�7�����G�`�4���NNB�X�N��@�:7�L.��w�Z�װj����K�-a=�`N0哑��KA{W�����ht� ��n�6�z�P�!�g����w��
����L����,�'�K:�>̰��q�J�ԟ@��Hs�pq�O�m��n��>��݊$�mz��%���n!P5Ly��C�n�U�zvQ��=8��:3S{
�c[��aV3�tDI�����NBb�> �,Ssl� ���nr"�3��
�!q�>E���Zo7$������`��{�^H�Y���k���pND���I�wW����R)�uv���t���T48ao��\��7����0�ݰ(Tc�_ےUfQ�cvA/��]��9���l~
�J�^�}t<�������W���9��}G1��,�O�9�o7�d��R�MPh6rdj�;k���&��U�FJd�r|^y�v(B������;glؠ��Ay��,-�;E�s�O�i����o��6��	Ok�nY��c����?�9�g�4�j��64�c5 ����~�k��I�����w2��x�,��s�% A`;�����.e|Bt� Q�����mT��!A��	�����#�M$n�-^�E���,QO�
T4��z�A
t��K�q}�2qw��l���Tj��N��,r[/���X��Z&C��3�k�3������>o�	6�{��t���׺�pt�M&�'��P�+�2ǲ胍jc;������d�{Uo����/��.>�N Tpwi���覉��z�𰓨�Z2V`^(
�ָIj�c/�95,`�u͚.k_���Qb��&���S<s"@h�%��K���۠/|��5ɜ�;Z���=��Z^��V�+���½�=���	�'�ؗ���q�;���A��$���J�EHRޜAD��`*;3�#r�)�*���!��/�M�;3P]�����������Ot7y`�%��|.�T�
�
U�^�~:\ v�ߐ�.ɴ,Mt#.禕��iY�����Ӥ�tW�Ɩ~�+�mp�А��<��c"��k1f<��}���~jp����5����)��\uv�e��(	2�^��r�1���+`QE������j�ָ�-����ו�\��С��;}�E���J��)b��gI�����1�J�
�;�R��!y){%�p���P1'oHS�V����A�,}����}��,�'
g�ȧs2�x��Z�UC~U:C�B;b���2�S5J5�0�X���W>�r�ܨ�wd�ڦ���ǓP4��~B�����j��Z�~��&2�J:g �M YuR|;�V�e��	�9���[�����Dm������<�������e����/��`��6o�Q�*��,�I�.-B���������n�ưj�s#r�����v��[!�<Z/�<39%ę-4.��#Q��l�xI�;4����*Ƭ�C�����t�9�1־?����j��&�>�;qj��
���t5�>�?�'s���]1�t�-�f OwQ�d�x�\�����NV]���Φ4���Ѣs��'����R�1���%y���	5wD�0YW�z�u�rs��h�6\o�^���_�_d����(��nĺ�{��Lz�,��z�PJ���k�ޯ���N���h3�ůT��&�<I��~�5�`��ю�K̴���Vcn������	�<�s� /ͯ1�Vq�\c�M�IN*���96/�g�B_� qu��hL�҇��aα8I���:�U�b/#�GJ�kj��L\/�Z&p g�,nO�1����_��I?=b��� �n��.*hg{��N+u<��aԣ��<�>9��!�#<��&<9:d�*�CD;(��6���K��:�Af%��'� ��ꦺR+��:1���u&F��T��τ�+f	c�'�N�O?����;���M��1l@6-��C�U����Ӳ�?��B��D�|\�^���;P/�$����ӟ�lW$��GUB��s�+�U�<�R����H�8���eپ!$�S_ -a�0C���6���Ac����^��`�ͤan*+���;E��##N'z7�O���.w
�_����9_�\�Ҿm���Դ9��DSgP�F��$(��p�H��$�
��/�a2�Y�;�6��f6��������(�%�,�$�8�wdF���u�@",�PolA��,���6��O�㌪,�Jv���TMb� Xq��[7�qƛ�"`G�5X��D_8?vl��A�dA����r���]�Bk�{��.Bʁ5�b��
�7�F�D�KՇ<>�"��.����w�SZsԁ���5q�j֍YW�
�n�+��IQ��4��Zg�@��?��<���`��VPgF��D���w�66�r$,�����o�ѕ��]�i�n����q�]�:�,�s{m��'(1R�Q��oၥ�ͻP��|$� �|�D��ի���?h-Ŵ�a֎R��U�;3�o)��TG��G�i�qH�z��T�(}j�Z��<�j��g�{�G䩝� 4-p�L�\�W<� c���ʁ�B��ݣ*����G��;�=� �Jt��O�as�qi}:[O���?�F�b�<�Yftߊ�3C�2��:�IO#�ɀ��oŌ�W�v����#��EzK}�sc���&@I�x:�:�!۬�MM}������A���R��$�" �1T�-�@��姂[.��$�x3-6L 9��'��G�BF��T>�	�"��`÷��,Qe��K�Va�r[����㝻��=^>�`�ti�p磸MJ:�YC�І߬'����	�O���/�}���;�M�h��;�����(V}m�vnc�kI�/:,K�T�����͚;�L��[Ŕ�w��9́��A�C!c3C+hyK\����JL*W��r��u�,j4=�����Y߯W��ļ�U�~��B�N@�����Ay$c�_i:�iHI�H�4�f��;:];���$c�·�f��@�?^>�=���Z�$h>�υ`��\E�����o�[��@�eB*��w�!TD�{�4���B�8�Ȱiev;~R�5Փ��S��j`�7{&D���X�n�
�&^aX�Ѡ/��}4O^q���=}3�o���9K ��]���Z�����8 ص�Zz���!6�G_�0�^����C��5�ܺ-�� I|<%~8jz:�Y��I����2�H�]�tF}�հgC�]g�<Z<��W袱x	]�G��HO�˴���#0��K6Z�@���M�y륷�پФH	��' "�P��}错 )+9�6G���\�N"�Qj/ �_���k�ж��4Y2\�6������o��<��xN%����7I˯У��(r!�y�
��r�^���*���q
�����e�������p�DgJ���v|�o ��H��+!Pzb��b���T.���M�ZEeT���W�3!�g}��"G�4(�1�9����.z�����L�"ׁ,�y����n��3a�A�`���=5�3(��[6�3��˩Y�~VN9��H`�H��NDIC�����5,�����g��yN��W���3m��%͉�U�ŉ�A��^�\K�w��5�n�˳<�/�h�,/y�� ���r��qg�wҽZ�0߄�G5w���Ɓg+��^�N���g�ut�vZư�ל�C������pj>�W�R�X�����ȵ:w����D����DS�7F?./r��`J��c��6�`�n[g��/�v��$�;�F��S)f��t+j�R}J����=+&��]�/ߥ_�:R�$�h���[��h9d	�d��֍�GSUCKQ�]���NJ�	��gcRQ��Z�5��Eaf�������nψ���'3�*֯5�N,��փ$�Tʪ�z�a����m�a@��D���z�ŉ$*��-�>���&>�̓7?W�	e7)�B��}u;fSc�.!��rzԊC{m'r|rY9)�r��)x��ۃx�ܽ�_�+��難�%�?��+�>j�����0��5ׅM;���¡�HS�]Q���S��2�⟲=c��JR����2ee�E������~w�������X�i޲k���(��+Y��&0\kAj/i���v��US����h���"�ɌK�S/"":���D6�/:}g#�g�V3�z�=1��~S+*�U7�<}��߅����	%�,�Nޢ6&���o�����|z�B�Π�x���d���\��f���@O�]C������az�^�]�%��&#F>�6�R�����@���JMmx\�; ��˿*6���r�)���g/���ֿ�Q-�����Z��>y������.�a����߄�	/� ���.V�]��A{�+� �,��Ba˓���)�������IX������� �=\rz��!�q{D�|хd�t����O�)�@��������|V�|=A:��]m�Ep�d����:��|��w����Z�SR��JvގK��ᩲ��A�u�G����ZvL�|��B���S*�	R��1�*G�oa�4��c;�uf!�.�1���H'��U(d������8�n����I�MDE�-h�ď�󰔾�B[�¾�v��=��,4왡����(^d���JEA��J�O)�x54��F�7-�*��HE�=��/Ѓ�aD���C�"B�L�p����$�,��7��M��*	Z"�}4E<��=.��|�޴v�I=�h�Gs*AUvͪ�Q*�5������u�Y`^�zk�^��X����{�(�kd̟�^��p�#B;�
���;�#�|s�����h��j�����8��U1Bn}���G��������rJ��R�g�UC����g���m�c@�6xE>��B��^����=�~��	��O�+g:���w�:��Y7�D�6�V�k�7P���T���u[7\�"aY�E�"|I��%A�ʚ�/� ;l+�n�S�E<���ȱ��ǔh��
�΍"��Q��E���vv��8�#Y����ɼfwbz�\�Rޫ�9t�X���m�p��m+�������M�s�����XG�7-�$
�[�p��u)#��_�.����4����Nl��g�yN;@�+Ub�M�y>�7  <�Wik9��<���b�V�1��uj�NP��4B�����^F5K�U#6l�(���N�lO*�#�g�)�b���L�s�	�=�����9�, n��w˂WRq��Te
�w�ݿ$U�J�8yc�[���-�w2KO�4-�uW�gn�ԑ8�@�5��E����&�x=���Z 	����<=���k�N��N���A���E�� �?*�R4b��'��7�j��9��'qg^'om)���Έ�V���p쿮�d�pѠ���Ɯ�R/A�h���[?g�	M5�t�6��U�n��m��3u��7h���N����Z�%�8��J�Ⱦ�2J��I��x-I�]�of$���#E�a��/t� VUS�*�/�b�z뮗�C])�rj��t$�9�06`��-��y0���A��Z�T������oO/`ۣ�i��	6v_=�,�y~P�Y��S5z��']���P��T�k���+����x���S1y��9ÜZnd;����G���bM�1�X碚���l�1��g�	����Q�#A��N�sx���':F�񩜘	�{I{���J\�*M��I?Lm�$}��	�n�������40Z.�y.��8����ן�%�k���֬6]�n$��y�j���6�ϯ��� ���G��B���6�16B�
�������PZOE?�S�V;�M��T��.�	������c{cT�Q�|�b��X��@�(�~\e���!�QkO��N��-Ix��Iq�3��=o����@�s��L�����IUQ����H?b+5vwC�Zr�C����OZ2�M�x�f�KB�g��H�p]�^!��������������Swt9w�6u�Zp����o�ҭ�f{�YdO�y�j6����3���/锥d4�\M���Z�Ⲋ.̚�y��������ߧ婰�C*��0��rh�.Y��IO:��P�L`�jc�d�G�H�^-v����#`a�ݠS��T���&�Ne��i�?M��`#�~q��uز�?Hv�n�}�d�`W���xs���m8��Gb.�٤��=Uq��>^n�5F�7�t!G�äig;�<�f�&�������S�#����$7��q�`�G��3��K�٬�2����i�&�D��Lֳ���YG�ˑ[�RS���Y�ѡ3J�\����
��� |<�);��]>�R�X1�(A_����K�:�۟;Dͩ& �5���f#'�%l� ���T�1�4�C�^�e/r>6�fچ즭^M��twr�'ݽ�����$��B��M�5P3����(�9CD>u��4D�
�Ț�ÿm^�ț7RƲLzSCb�A���%��t�q9wO#�*�ؾ�;�b3�G�A^��\K�x�Q�A�ǥ��q�s�S��Xd�%@���yG'('��%����:�+0�|-E��(#q��f�0�����>�Υڿ�=Ґ��	�iK�ӦT�4�D�>6`g2�_dП���hԉT8r7Jr�c��b��C�M7�ui��VO-�l�z3�*U96�-�T04=.�t�B��t�V���7۱�ވ�CL��Ò=�E�e,�16���eƾNN� 1�-b�ѷ��a�y���b/�Q�KJ-��#im�����'��CiY��Ӽ�I�ތ�,����J}�"3��,�..	�4��!�!Wm�1{������W��P.h�f��ZI��4�/����Δ
j9Q:Q���7��Ԩ=��6"����%�$;Ȋ��!'~a��R�|������#'tR~�5�T����~N���iXT�-ig>��B��إ5Fj�$����t�ԇ�D�>�mz�����Bm��O	f48��d2���x��3R��T�r�q̞�~Vsx]�s�_ڊm�}ݻ�_���ǻb�v�j��i���Ӽ��,:��8/�ðz㫾��x�{�.v�N�{ =�G�u�{��V��Y�}v������]G줷�}�	C5۩R4Ɏe�y����!q�I�W2�v��5��pR�&.��@lkٳ�������O������3?�	g��>����I��8����޻���:�z��'KA�nN|r���W5U�*Z3^�.�[X���@D�I�>m��7�n����ꋿ�*q����/�rn�圞y\�u!��6h���$��w��9�ʬ���l҇�)B�/-b��^������bc�D���CkƠ��o���YXF�LwA��@\":(񣂺8��RχV���b)y��O�_LB��c����6]|f��^l������)�|]-���(�#���b#���b�xk�ѕRQg�AP��Jy�H�?}��IF+���l����v	����2�A����kU��>b��酝��_~�^&�9�31��GZ�:��Zр��1���T6U�}���%[�[c@���}�"�I��e��g�N̳L<=ߑ� ��&7�Y<�+ �+�xL�Z�6
}�M�?��a���Fj���/9��N������	�Whr�]��c4�nVhS�D 5�~ya\�?5���Q���(؝��Q�9z|����_�GU�o�����(�h�ɉ#���Q��qvE�]2L���~|�e!"��Y�X�T����?�@̕����q7��X���iq�B�Q��O�l�zPy�j��:9ߎu�6X�9���
���� �5q�t�mJ��/;��J�������y@�TRB9��2�Ӭ�d*s3���!Z&_���A= ����=H�(�N�͙�wn�u�T�m���5�˄�b�U�/���B��c�
�Tr�;�$��zQ�	�M�#�;\�Ao�8nJ_�
�xo��%5����p��_��<s�
i����Q��kh�l"ަD'���gg	u��fX�:����j?��:�ö�7�7y�u�i��NH����Q��%��@��Rt�4�]��p����1i�@�U�,e#0~_�#�!I �TPj�y�j�v��W&n��euJ?�Z�~"�m
�(�Z�dU�ti'���XoF�}��#֘f՗~�*�Y	9���"�ǿ��/ϴ��1@#��8s������}�Χ��'�(��9n�3]M�i/��yޚ
�dDw�O1�)�9�w���ϒ̛d*��~TB�&���w�+xO�}K�<���|���| ����r�K�N���.I(�#��Ds��r9�	����'�6�>��F�Ff#L>z�V��ϱ0\�9;
<R�с��3��č����3�>t��Ļ�Ɍ'P�1�Kg1S�q�|�V3�R6���oM"6��z�,^Leb9�4��;���('<}m�wN{�N��ZeE9?(�K�(Y*V>DO�AN�䳜� 璉��=��S��}�}���v��	8����Nz@�>�i2���];@�c�琮(���/���$��t�f�=�*�0+�nQo�T��~�l]�}�Z&	�g��"���z�|w;��X6<��C��$�4�^.��ˏ�{���Ί�F���,?�z�t���<A(�@�%d��N���5�j,QK�gM����۰<�Iӟʺ�AUQ;;�����8��
�/��=��\ �iR�h��0�By����;�
2{?MP��I5{���(�ׇ�NY��c��H�R�������������Tr hȉ ��.�[�jY��&�z��,����r5֐��2����}��t>�a����2B.'���H|��0'lv��p�2L�#�g�4rtWj��u����l����q�i�,���*�V-Svgs�[U�)O��Tbx�ũ�^��K�޴CIT5��ә�b���Pp�w��+[����{�*)�j���W�q ��ry�,0��*�dg�b���H0־Kh{��f��+��R�V\�6Z0g�
�(��J}<��|��)�S6��1u�p��I��]s:�R�~ez�����	��P�߸����%�+&3�Nϩ	��I(x�3��9Ɲ9V,r��]�֕}ث�ҺW{���=��S����S;�YP6+h���R5���!?��ŇG�kj��3���U`kѹ{�x^����*:--ӳ�hvz��E��9v�#]��ӝI�R��sB�M��,]�ؾ��Dv��li!L�I��m_`lNYp ���>�Mځ��dB�K������2�[� �8���͘?�Xh���}*�z�\�2��߱�Q�N�d��+�^��GF΅^�27B�����|c+�����a6�p�_�P����#^�3V�9--��lIS|*�@�5.xS;U}�Ƣu�3^Qx�:��+�U�RqX��{3�a���N��
�+?�2/�<n���y�5\>XT������\�ͱ���!Zq/�'�DzXt�ꐥ�|����[��B�7��GSE�D��FO�X�0��&�N���q�S'po�8S�w��^�\���5��
5���&h>�I�y���w�/�CX8{%z'|��i#;q@V�o8���brfM~#;ɏ)��s`!�8H(F�-���)���
�w��3��V��t�|T��ͨ�Lzc���``�)�ޅ�R��kgZn��+��'b�p�8;]�T�n���[��7&e�u����s����Ԓ1�l�*���֤B�ތt��j-l��_�7�.q�+K�Ę>�p4�U=d,�A�0�*���?!���'�Q�b�a@Z�z^([�.�T�,��+�!��c:m��]0>Fmkt�5�+�w���+Z
�=9�0�yV\�����z�ن�x��X( �	����Pu���y�`���c��Z�u|ױ�BR)V��L2�w_���V ��2��=�8��a8{!�F�@�̕�9]��:��3H^,�)�'T�ez���H��S����Z��QW�y9�ʥ���������~%T+ӭ*��I�R/�+NR��F��Q������R]������X+x�8K�������-O��*��1��@[��mf~�A�b8����߰��U�m	����6쎆�B20z�4T�-�ٖi��W��*�W���Y�K<}��!A?Y��B���<f5�>:Ohb��@�ԣk�ݤ_�3����y2ψV��.�RK�ZX��*6v��[���6���3]DZeq!⌲��Z2�KPY��}���r��E��D��H�&���4�OE$�f���ʯ��^�m=�Po����F�X%����$t�F놰�K=���z0>�7�	}gW�^sp��ø,ߡ/�ϊ�.�3�ƢB/_pWEPt������k�IH��/���zEYŏ��i�2�����ȓ�8���+�R	��R��UL��EK;���{��2��n|��6�(�����3u��i�H��+٦���ȼ��O�V���WJE�rZ<*c.�����I��bV*�y/.5������$&�ma��ǲ5�}�$����cݏ���\FiH| {=�ag�I�����R�ڻ�>�G��O�+AX��f�� o-	|YP��P���l�]�]5�d0d~�$�F��Š-zؗG����ݧd��G=��
�2^����a��o�eΒH��O�K0�֝���0]���;�)��ƴ�fi����*��N7�rN�Ds��1�+K;Ӯ�,��u,��"X�U����g2i�&��ɝc���ZmLZǢ_\���ov�s5�R,'���i{Z9���9W�[ހNì2�<寸g1?��@O�zR���,
�ew"��i��5Z+96��|6#w��j�,�M���Z��f�ց�����<���?�~������E�UM��M|���m���2�dQ��1���+b5�����P����<A�H�>:�V�z��CU#?$��.��5�3Y���P�w��ku:�3����:P^v� ��w����Jix7#�5yvݶ!��D�4��PT˯��?c�9:�V�OD� ����GpZ���ҝK�H�����	��t.���`i�κ��Z=�e�Gnur��t�C��	EwB`�06��Tl/D�w����f��5�#�t�Y�n���5LO�
Lx@�9�{y����3�nVb��i�v3�eϤ�h��
��l�[|Rs+FmI7�{G-�0��ޢ2�8����1�\b�lw���w9�\c��;�UG}���9�3���G�@�ե�(-��;y��7=����v>�?�!d����@>q��.ȩ��$T�|�ŌHL8!E�`m���:������*[5m�G�7�6���{v�p�_J�0���F�T��"5�Bƭ�i� F�uY\�{o��bb��T'W�뻟P~�.�InC��(�x�j�	�׺+��=υ��wC�ڏ�~3��#Ï,��Q�d��^��\�~<_�qvؒ�z���'�gEv>%��! �MyQ
=I�"~�L�6%��YA ��4_$\&�u�����׊ʕYȲz� �y���^���>��ddh�����,A��K�F��h� �����#?�*��xb����j�H] h��^�B|�#}Ҩ����]t��R;���ǨW����T׋ ;����e��C���rm�"� ��s��YWA{X� -�կ4h�FOU
�\��Wj%�h���!�aڲ
�]!+j��xˊ�e�s%�>B�c����ZFerR�_����]�_s'�J�?jj����>G�S}eg+e<��_ަ�)���K�!�S��&1G7�۝2��vj�#�R�Qd=�J��X�o��:�vTCo��/Wƙ~B�3����g�Z%(п�>�ЁTD5�2#P�0�2��}�VX�ge8������x|~7\70�}��)�R��3�J��o��23 ��;�*�5����;p�uB��mb���F����Sm+���n��+@�9��c���Ѿ^i4��N��=�A~�}}T_9�kB¨u��4����I��T-�A��P���"�wO�?��k�8����ϋ^y|ϮH-ȵ-ma,$S�}�z,\��
��L� ���gEp?����SO�*��R�9R��b��Q%F��qڗ��������MІ����k9��R���\����d�y��s�����aJ�"6�����9�z����[�,�mq�Ȏ��w�*��ϯ��+�^�φ�$�=��ظ�]28=ʻ��k8�qJ������W��XS]:cDܢAv�ݤgY��Z�"����� c�+�G�3�J5���E8����ܛB�\v�0�Y�Ċ��nǟ.){0�0`��9=�UF�����ُ����C2�~�왲�&I���ܔ�u��Ķ0��բ|"�hZ�T�m�?Y]�L��|a������Yl�m��x#)��y��kdz����*|f��cc���m&�n�HE�� 㰲J��ks��u����+���s �Ӽ.E!����h��rؐ���G�㶵r:o5?�7Ԉ�a��j��)����ΜZ��ܢB�����^�q/q�\��^�s�����Ya��Z$�3�g|V%�� �K-J˷J��0r�@a�rWU�u?ҕ.ef��.6	���`���@���{	����E��(8��5���K��*�� I�G<��5��_�(�!�i���#Fi�lɝ,J2W�E��8M\�%���.r2f�/E�ڈ��w���^I����+��t �E���/#(C���s�[�JP�kXw� � >�b�[�ZN+���$�a�|K���܄�X�b���uy<޲rT�5�M�q��?�8�J��3�( ��ٓ��}�����Th���0�����P�-�A�>�1|�E݅v1JH٦gB�C2e�>b���\��tl�éF��eP{�!u]7sz���U�PC�C�ac��$D���㟌ރy������ `���i
f�*V�:�jQ)��}�B�]	�_+bZ��<Y��::j:���׺?]�v`�(Q��M�����N�˞�	��o�H ��.�<����b�ITS�i�z�K�"��������(xr��H�<e�#c����j/R��䳲�� F(�Rꭂv��g|Yw܌b �˯7�z��׾~ ����-[�8�Hs����-�&�Z�L�!kx_H�|��b���@��U8��������eem�bB[�+�K��G�nk�<��"J&+U��LEB1@}���Ψ�{4��XI|����ب��Z�Sl�0��Q���~*h5���m*�9P���'� �Ge��	���S�* ߯]�t	W�C�����sG@�Ӱ#i�u�y�#D�-d 	�5�3gFt�m�񷊰��"�F/7�k�̪:�ud���(�1.�(�Y���8T�3S�����@x�lT�0���QD��=UsS�-�4�9 ��Ԙ�|)΁ۚ�o���V�*BQ�7i����J@�m~��B֖{H���9�8dVV�4�BJ��#�}T[��Lc��
{'�bh�B�Y��Ԣ�G�&u��d�i������1wxa΄�b�-���=�Ts~Є��8Sx�-#�J���s���^�9��s�AF��=���z�<I=���&�3=��?�N��k��Lh�����D���k^�	>d;��w`\�&��0F���j����eؾ #ȬV��g²�'�L�s�.�,�F'���6�i�4.�v�A���P-!��a�l��J_�F�����}��\hZ �|�$�B�v���O��Vg�y��u��- �BZ��0�6�q�A�f�?��Y=��F۟��s�|���VF�_�v
{uGb.�+�
���e��E����}�3��˟rf�����i����T�\Wұ\n�D���l����U��f`������������l���ɒF`�^W&��ٰ�h�o�E]A����	���1���Ob�B���?����g��Eq�qEM��X�̔���p���I��a$J{P���r�_�	���D��]Si��e>��A.]P�
?b����M��R�TN����s�+�|B���Pc0S��8Y
�׷�%#IT��/�5t`h]�[B9���򎥚�I�L�F$oD'#��nSr�g�����OF�x�0�����8&����N	U�އM�� c8�~��sG
EH�n��g^@+��� h=M��?�*�����TD�Y8��ьz���yT�����v�5��Sk4&��ue��<Wg�bC�N��|���q�3���(/4�n�	�+k�<��t�8u^���\���
\5��)���מ��s�7��+M�F����5%Zo��!sNY�u����o�"Q fIH�Ӵ�6�.*����ܸ�2:7���-Ο�ݸF�5T߳"Kᣒ� :�!Iҷ��~Y��� t<��?��a��W]?u�'b��c��(�ٷ�,xcC���Q����
����?��l�G����D�pT��^"D�q�OQ�8B����iP��_�tÕ�My,daV��%��*lҀ�`d��0�9����xt�&�3r�;M��*���ʞ"���>zx�.[;����]����Yp�����Y��ܕ�G����5ٯr�&'�AV�l�t���|�f�H�r�Uu:e�j|�Ȁ��v{;g�/�����X{�OeԞ� q�3nS��v
3�1�gZi[=���5Oh��5Y_��5{z���؝�z@�r&u���Z���Ȼn�Y+�����Y��@}@}/���i�̩�)}��������Dė�ٛM&}T�V�X��S�H�̨~�,E��$�������g �KT���+���b��?�X��˚���k魌!U̬�y:|y��=��r�.6������^�j�a�C1x�މ�PO��t��0���W9MoU[�;d�L�rQNF��^&�m��<,J���߼����L0S��0"���/Wg�w��M�Ze���v�,���h����w��> �����ƚå=��>�����\U��lH�ȳ(���qPõ�܄���ŀ��˭��i5���6�U���:�7��I��?��"$4�6�� �ɖ��\��@���\7-*|�J��}�B��.��3��m�n���fs�������>�!z��"²��U���z"�28��;�!���{P��"`m2<�.�������8�k�J瘑�����w�m��o2@�S��VI8��,�� �kG_lS� �F\X\��D��+"YA1�x�+���o���v��IU0�|�T�k
�y��qN+���=��V�Χ����,ڀ���wi�7�q{\m[)�v���+�S���	g&B����_-i�Ѱfb��/?�_��d'{B�yYr���""�������K�y���r�+N�o���08��%��L�	$@�'���S�&
���g=��YIg��ͬ��A�~�Q�R e���f��󌥜��%7<^wR�~����x+������1/� ��f|l	�c��F�E���	f>�7ɞx?mn�O��f�w[��R��?�)�T����
Ɔ� ��ύ���VA�m���GX��������R�0`�� O�ϪPfA��(v�9h��W��V�S>W��O���]>���wA�q�<�^���1A��n֑:�b�Z�j�L7��Ѷ�
�X��^�"��w�|8���'��qal�%( xn�>J��'�-ĝ�p8����@�;�?cH��;cs��Ɩ�+�	�[�v��j��Y��h��&i*�V<�j�`��R[�������?�D�3����2�F�}&�5��R�E�an�o�U��U���8�L�I���ƅZ���_�إ��%���P�V���_9/OsJ}_��r��f'��+O�ag�K��1���.y�W;f�:�+]c�FF� � ��bY.�>Yb��t��R5f/d�����ԳOs,�a64[�<x�0�J�-US�<�Ġ0y��7H�˻����,HR��.9�R�/6I��]U�@�MlA�G��H]Zm��zW�-�������i��8��q���3�F��T���x�{���,��;#���I�anpLd�T+q�8�W��
��(z{8���!}Fi�� �϶��bL��~�/%0����1�׻n�k��/^:������o�	�_�-�M�i����:^����E�I�f@Q���Aa�ۚ��[�=�È���E��ae7�.�!?��n����l��a�5|Ǆ#����dסs7u�������:(dR�Fer����
�w�/��L�Km��.X�u�((��&��'y�c�j��Ԝy�@bi��E/�;�L���)�X����q�FL�$�9�0��1U��-�w@#F#��$:��d���6	[��k"'/��<ƽ�ç�J��eKI{8@�\Y�����`4�%�l0��yX�oX<�R����ee���8+������Ɨ�����:R��é����5?���K��,��C��k��gL�����=]���V�#���r�z��Çt��?6-��!�ċ�QF-į���vgl�Q�y����=Úg��B<z���!����$r���Z0x�h̦�*��ZA��Y.(o,�9��"z�$8ӗwӈ���Y>n�#� �������g����Kc���C��a���er�Wǋpϓq����cp�a��Ew�"5�A�՞_�,;Uk�3��OT�=neL��9���x�M���Чj����ӛ�c���;�D'����tXC��;±�s��"%��+G��bS��,�߱[ѕ-9���!����Y �5R�m��%��U�Ms}_;꜍�*��O�߱�6���@���i9�\ܮ��$��u�'�>[�
���p!p��ۧ�ǋ	I�"�j��f�J��䦤(3l#��F7@�H�6���H�F�|��,J����{�u��!�v$*����b�_�vj� mG�&)g������Ua
��D+�_@S3v]ψ�Y���UYq���^x+M=��}�tL�+Cat�0PLCy]�ކ`Q���W�!����1X� ,}��� �p�Y]c��U|}1~}-GKx���A��PY@�ȡ�l4T��ɹa�G2A���ME�ig�q��
k���1<"%ە��V_z��3������X$�����qˏ�xjF�8�F+�̊4bW��)��m�U�
zZ|ۦ?.^~�:��f�س�w:� ge���.�ZZ��x�[�(͋vsgLfg�/�̝!���J:7p�?��~��/�5��Z�>d��E��y!YF|�����w',&R��e5�F�:=�w��	M�Syo��O/��,���������T�;����1�V���}n?����4 o3�HoǙP���c+�Zר��|�r�+ �̕#�&&vT��W'О8%�ۯ3/��M�hb8�^^�̣A��N^v�Yj	�^����鄳�@mx��ۅ����<��~���,�3S�����U(l5;2��B�U�`�ʡd�K]&������A���2-��$� v@��3� 9��gXqdA���%Ý9����������G�L3��A��^-Uʷ��9;�`Z)��{<�lUM�Bu"I��y�q|~�e�K����qjݒ^P��3��$5�h?p����]�Hh�jDM"���vod�,7L5T5λ��Ｃ	|谻��׀���]ܟܼ�g�"�';�5\/1��P����Q�k`]�`?�!�=u/?�y��y��;+5E��M�K�4���ZB��ҷ���0[�Lz�/�'}<]��8r�P��ջ��i�ಚf\ �����=�E�Aҍ �VeO��
�ppXU��{������m� o(�/�#x��̾��UӖ��@��Y����öy�c`tW��Y��ʳ�U��w���_ɫ+(�	e��%d�n[3�2�동���{�g����ˎw�����&��P��u�q�A��,��d��Ϲ����*Z�/˴#;d���a%:�@�A0�V4@󤥻�z`����'�4Q2�y�Uߗ�W����/���u���u�u+C]5�%2{�ܲ:As��n��@���t���2 �� �W�hOX���nr��h��װ�lc�[ʯ��Av�x�A'zc=ٷ+�<�錺�Q,��W ��Y��@�]h�N%}��ژJ�{��?��ڥ�u�̧�8v6~V`lt89�u*�)�����&���g�=�-��5㡱�1��)dp?%�����E����E�(X�?��;���v`4��<'%�`N�ⷫgf�m��}�e���K#(Sg�Ɏ}@]q-�9=K�_p��F�eW��_�	`P#��BOG^W%\��{S�4;���>t8u�_�܌g&�۶��˚�^ޝ '�O揎����P�IN"¿�y212@6�(d)�A���qZf���4S`q%�zt����Z�0!=�D����b�Ȝ6w�Ǹ��ٲ)��L�qyX[%�;�$��v!5%�j<���WQ�&ir���@tm���ǟ��e�syx"JGQ�*�x�d-f>O��{䁭���kɫ~H��Ӕ��*������4�t�DI�c��=V�jہ�Ӹ��#'f�62�;�OⲰ�o�%�s7�����������cFGp9����P��"Q����f��xL*������몱�AV�_uy�s�M��m2'����n���>4~��i�U�뀘��]�@CkĮr�=;��3� J����I��g9N�n������pE�t.8��[��>q����@^����)�M��]���� ������ pxG ��D��)�hL�B�M
~]��s �J�H��h��\ �)4�Z��gΙI�t"�$7��שo9��1Dr�g$^]��C(+{��ڀ V��\�DM�+6$z�5�֘<Ct���4�c���ڿv��
�^�V馃S�oIP�Ύ���K|6����3:ut����n��_������L@�(��-5�,\nv��8!ZjևC��TԥQ��a3���Tь��*%�����d���Rm������U������^3��5��>U�gO��fa����3Ҁ���+˳��=z�w���hmr�h>3�Fz�̹�
[y��X��a��a�:�Q�E�K18��u�!a�.]����U�VGv�U��S4�\����T��h�3N�B��g�m�R�X�-Q4 �P��E7K)�62j�*"(��1/��RF��}:�ji�X�]��u���0�a�>)0��3��_��(�G�tm�D^��=��c����q�E<U����`(�l+Eز��H�3��j��_6���hz���A����+XT���a���8� ��2$��Y�Z`쵯G1��|SނT��֕Ǿ0���g��sL�u�����G���U��Cr�����"�2bO��=:��YM�5�+j�L�O���kt:�H�(�
{)����cZQ�nmY��`	7�������4�F�����䗢�$�����(Ψ�#f!�a�o�g����!=�%^���T
�szXN�/��ʌ���	��̩jn��g%��dA����j	��Ќ��:.,6QzhXi����&��+�����3+{�KTxw�����k��?�P���ji�>P�Խ���;�
���ЍG���g�����C��=	\yh85�z��"�(+�����_�ۖ��.��^a��ؚ@)��tE�1w!Ē0��pr԰ه�ib��"t���@����l��M�dy�<z���:�f��~�V�A��i�;Jh`��w>��ԉHc���܏�TK������d1ꅴ4���I�f�}���|Fк	0~���J�$�� .i;`�c:��o?i�;�dT�}`��K��ĘiL\6_x߉����6��\?:�c��[?[;��p����B0����V	k��G�a�aTBy��n����$'���b����L�"(1�VP�}���G��Ϊ��D~��v�U��{��ڄ�ѐ�RQ�a�E��B��p��<��V����b���D�@/���g�����-� '5��!�2�K�� ^4��]�wo5 � fT�N�T�%˦�7*<�O�DW���|�-�`���?��x�OPW*prPSa��63 tA ����R��"�x�����"@��!�������-��.pk���毚�K��;K�]6!�3�WZ�l��;��������A�h�DV~� 0{!��tup�'-3���?H�M�-j,_��?z�n��t�OڝV~j�?Ć�ћ[�5l^"��a0q��ˆ����3�hj�t<�����z=�S'�#�õU�co%�'h,!�9-���c��&�藶rE�$Va'�L�b)�bϹ�vR$�r6[	�P�>�3VCL@���Ә
T�f�7�zVR<�2��G��`hg�]#p`�^���(Kw�6H&x�l�ˠu[΂�`J
|�;�t��� s�گɐe��9�|e�{�������W���U��x��&���x��袤����tsv�f8�xj!��v_�mg�����hX�i,Д�
�SመK���us�"�s�S�;bNn*��ޒ؃Ӂ��{�l����!�1��i�\{�?�c�6�����Xh=�����D_�d�3���U��zo�V��?Bd�eŮ�o�WB�c^��6���X�TS+���I`o���)���OY�QF�:h���a������*�\�!j�K!���y���O�f��a�Co��]V#��É^����㸧;d��5�.~]�#ނj]��.�����GA(vq	�۲��'�|��j��ҩ���ʍzյ�a2*�s��֧��9��K+7�W`�{���V�b�Ov|®'�O�dJ�G2i�|iϰ�=��8�gFc�dgZП�$�M/y�Pi	�a���H� Ą��ȑJm�1CC@�ӕ!�����*�n����"k�������m�ϣ����h���[�ӭG����n9��ᑍ��b��"�P�~Q�U���J�YdpA�ؤ�P�]l�b���tq���y��ۦR�_��C���M��F�E�����HW��J�>J��Ot۟���6]��b:D��.��6��y��`>A����BI��[��7��Y���SE��]��_U�h֙��ڑ�ڽ}�������dr�b��@��ލMQ%�_�Dtk~q��!M$.�;��U���ߏ�Vy����"k7@��j#,��t�H�iJ⤖FL���5�ڱ��CU��~l����z�x3�.H��[s��P�<u#���n��iZ����<���oL�!8�h�1;��g���qE2�ϑ7V����"ѩ�2���u��%�I8�tņ���Z�:�4Qs����J�:յ�I�'���#p �)�a�9��6q8�k�w8w`9��1Go���T��j箳�z���u*����6;��3EV�n�c�Q��ڲ��D���b�s�� F��C�4�jrt:�~��?�	����F+	v����ID��fc$ѣ�Z��p#�g�Pӎ����in\6��
�I`pV�9�]{�`�.%B���4('2|	������S��%��S���A����8���Y��z�����={��ﭳ���l�1K��w���ǋ��j���lT೮�h�j=(�7�I����ϗ(�/>�/�Y)��3���9n3�����T/� 2k'��7H�dP5E�g	FSbRd�7=�mTAڗ�_L���QI)�:�`Z��<L���-^ޣ�|�f��R�yh A�	An��yH��7��!���Se���X�
]����a�V���%�iV�ut�sR��#+�1Ef;�*J�u����\G�17�#���L���x�ɏ}�=�&|}0j@�u<��)�@�\�}��(w>_G�7�4�Bꗠ]F�c�bc�!�ɉ�kC��˘]Թ��ͪ ǲO��Q��K�D�i��ݾ ���_kT��m�_�fU�u�R��1-}k���B��l���^�*=�Ȳ+U�2��>K�ē0��&�w���^����%�Od9|wuF�*n�VAS G��K�RMё���@�C�u�o��q�� �um߫�f�	\�ҠD�J�S�F���X�H�mJ���F�?��J�)a�Oz��2��v���I�`0+T���Q4����LO���������˪H>ssA>}~f��u�"ցz�0P�P]�ه��oK'���VR��C�o� ��+�9�I@NcS��kr�oP)k�B;�62U�aK�L $O����N�� ԯ���+2�)Ȝ��oB��|��萙f`��O&[�f��e�7���mF��>\�s����<�^ ��5ZX#ha���ɘ����mdW�y/�6��_}�4n��=A�@�	�m�
�nOF`����1�d���0���Ū�4FuAcB鳴/%7���AiZ��FĦ�ĥd&�l��v�j/6�H+k~G��2�c�l���p��Cz>��B�ِ`D����Y��P�j�G�����)�Zm��`9�
5�1$��8�%o9�と��%
�6�M蓝���˓Y�I0�w4�iR�Dc����J�x���,�XǦ���-���)֡�O���K	jS\-�vb'MWv��<.4�&�V�ُ�DY+0UR�=��>)�$v�����p�|��[R`�Ά@�AY��e��'5��j�(�š	���m�|��N^S-���č �ͺ��f��c���[NYhC���}	������:_��`�;Й�ϗ�=F�K����y_f��lިi�ҬR��'�����*�/Xᆝh-��	�<���p4�n}�z璸�Έ�//U��c�G �v�����1�0�Z��T��<�>6p�����0��/&�4+H[�����k�3FG?{g�"��O.範,;�2܌5v�Q��{��]I1�j# �fO
�3�l�F�C�hh�o�ݥn����-��T���B:xJ�b�'#x���c*�bn��N���$�s�1q�G�Ծv�n�V����$C̹с�?����󿉍_���T�7��Q����z���$O���u�Z���/��#=����^ߌ]�)c���1���' (*!q7��`�_|qS�t^��j� �GJ�dPЎg�L�&�H��g�r� �fY.�^iF��^h*�y�1���q�t�m��p	�8ؤ���S���'����8\�حjL��}���	���!���!p�Lk֓��ٙǀ��.�ܓ����#�d��	�{�UDT�p����[7�X�a ���T�Q�G�����{�У�p"C$��0������r?#)�i���fQ�0��Sm�V}x�
7�y4���,����:����AyF�������N<��6>�A��Ę����Y<N¼'�2��`P
���� �u�k�ol�
\l�č��^&V��b�]f2�����h�v�(�G��i�4���p����^=!��[>�L�v�~:�75�&8�f�ގ���v׾��@mXz�͊_�� `�y3�~�ŋ��6�)!i	@�+���ht��9ލ���Kw�/�r��!�{ތ�v��m��g�)ϛ
���n�UxW���%wZ���;�-�W�C�S�MN�����7O1��W�Z�n߷l�-9��c���h�.&�؇�~<[r�Ts�����l�{��љR�ՈXI���j^@���f�'>A��k�&c)%���pFP|`�7n6�N������g�r@'l��mf��JЋ$���������sՍ���a /��Y�]��j�q��'�Հ����W=^o(�>�D��ϯ(����t:h�g���q��\�!t�ȉ�+�F�(T�����T�ߙ`Z�DOf��=Y%q�ɦ�F�x�"�H��{��@���]k���(�u�����`�]�����i�Ԉ�?rs��.�����a��W�4��C��-����,��n���������tuFI�h;K��n�IR���Nfd��'��W�	�������{�1��J���L&�,�gФW�����&|�]Ҹ/��^((����$Y/��㺓$��%��$%�r���,��<�  _�]��[�<�>����.�v:�'�
�ߋE�a���ibi��&b���b��e����y͙ȠY��'@����CV4g���>�B��{Y�cWr�^�m��}S
z��I��B�gd&�����,43�v�5h�D;���3��$��^�CmI[:J>W��Is�5z�p�}1�.��=�N#s��[&�j��1���0�e�}~O�%���.����	IZ'�3���u���VF��|3��/}��WU���Y��F''qSY�RA �U-M���s��O�hCԣn�3�D�ь*����K�����Le|Ě;�)�p%N�	?*���!
�����?�X��K�q~TӸ?�1�=V�� �ɕ�g������ňu��>4���HsϠ(,��zɶ8�K��� +��Y$0���)�¤�|_M��1������{�D{�VП+[��Lg�ܡ�a��i�kx;W�h�����D�j�@�V:%z�te#&k&.eA��Q�GR'X'��J(#;/�)ߊ��q��e:��㜎)r�*U�!-�MC�������1�;��L�����AB�YO�V-��yz���߾�<���5z��!.Κ}x�G���7�Ưӟp��\bXN��^���M+�fҙ.ڔ�Iq���-`��+���x����q�7���
�s�6c��Jv�~]23b3X��ʔ^�����)ˡ�>lzD���`ėս�z����C����>��*	���izq&�d��DY��n���z^V!9�߄�-�B�<�TN��y8+����]�N�PǨY���,{!��ArtA���� ��N٘j�]""�{��p�d7fP��,QSwv3�5��&/jݕch���9��Z0�GaU��%T"�*�d��,M�9yC��:z<��a�vP�'�Ti�&�^�b1��4�0E�wI�[c<jp���mp�#��`8EB/ު__�[G��+O�Z;Yf����*2�� ~rT��O�V{�]8S�4PQM���eD�_��J��%�@�J��u=|0p�DO[��O;_i�[�������ĺ~8�Z����]v�HcW�>f� \���ى�gM��'���&��^�a0���쯯0�����(n��q�����f��r���-�����3M��N��y�Bt4����@ň'(;D8.��xv7N�y �T�P+(R��8^Y�ٍ�`z�"|���
�O߲���E\X���t��ʹ�"���è��홤����{(���pC�'��W���B��Fx�l�EG����ٓ@[Nl��|;�6xXWVxvD@��?�_|����<���}6��5ϝ@�H����rfD/LGb����ň�ay����>;;���^L]d�8?Vսh���lNS ���1�8\�1.kb�P	Rsѿ�ZmF<��K.�n��ἫW�,�}����&�K�P���eq����_�
@rZF�Y�<�7��q/@�Wm��Hs�G�e�����ܩE�;�JL�~}]u�ז'騔�4�gC��-��ա�+t:�$4��":�u"8�?�S[��n���)�-�eH���1]g�=��(e[9�P2\������Y���T0L�n��}�$
g'�rp;�%rC�Q��I(��/m# �i6v��>s�Y�� ����*�ڣ�L��R� �P�b���Η����9ō��_=�ԻtS��J��k�j��c;ɸ�M� Հ��[b�LaK��ɔ�GЗl�t�F��9�8��2�$n(�V%�b�)���b)l���*!I.����b��W|Q���NN�Kz/�o�)Siߊ7E�C&���*6bd��y�b7�uDtR�_��8��
���?]B!�4`����2dmXVc��z5B��.k������C�_�JS��5����t�2)#���!=*���"�%@D��ԉ;�	�<��%A<6���[!t���mME��'��\���C�M���΀�V�UC�|q��������&�If#�%��A�	E1t5��ǝ���נ��'�y��l�ag����>_:WK�"c�J�8ә�;�]&k�M"'��y_�0�����m݌E�V���0g$C8rg�.)�*� P��2Ԕ���ʠ�S�_���>Reu�H������圬����|l�M<C�f��8�T3�,ZJ����dղ��A���Rz	=����Y�9t
R\W\�':I.�wgU��	d5�%�X����Ry�b��ɁO�S��>�:��~���Y�T;͇��'K�n�����Y÷����o?�dpv�f9w����jr�����6��j�=�QC�뽌ø ��\�dz���}��m�ZϛL{��n$y�wᘩh���Վ���܅��v�B�_�(�e���DG�be<1��y�������@ö�͛9�,?���>B�2[�\�����3�0b L6�x�W>�i����mHk�˜,"��X��*���%�F�=G&q':X�
�U�d�H?�Q���6�z�K?����<��N~	 	~9~�#xqw�.�Vn�j�j�橣!�<p������K��UuB7���=X*悘jR�����'
�m�� W��R�����O����2O
�Sl38?Ε �ڸW7�C��y�B����\����K��wv�������.;�=Jg��X�E��1*W+�
�]�Y�5!�	&~\oY��_@M�]/���l��,ƌ�,��A�u1���?In�J�
�9� �͇9����.-zC�b��ۏ��5��:TJv\P<Ķ*ۥ٭�-�Qz�䉋.;����r�y�y��/��!=�z.7s�G�;v�@+��E�Q�i�>;K�4�4Xx��h�Z�:HH8�,�YPu�Z	���v���fg���!(�6\Tz0Gq>����ĺ.�\��A���}��h�|�~��v����j�R*��-��30�y��#e�Q:ѹ��RPK�Uġ����x>�rNK�3��'T���K�w�i��Ug36c�Hb�7Z� ~��X��I�����(���z8t��$�w�Ҙ��-\`�<ŵ:~�úI���ݡ�5�+|���N���V�g�{>O}����Jl�Vm��M��W��WD�z0ÑjD�S���e�Ssݼ�*���JX�6��~G���`bÚlx�vh�H�Պ@�$��,��<���o���0&�-宰�F�U�}1��R>^����$*��������6�h� d��iO����Ѭa�=g7ޚ� �������v#Iԛ� ��\hC��`�#��H9Dol�����*�ɿ?�6�.	�>�9'|c��:Y���]n���ߛK������El�s�aN�s~��3��$��)���;�����k��8��.T��Q���aca$�<��Pt_`�C�'3�~}��F�&:�%�o�z��P��eR��fM�g��xWS����1��f�̃��T?��=O��2ݿ��L9CJ�򏗍��K�~�ݗ�-	�W��a�i�3��.�<_���s<��`c�E�u��l$	G�xѰ�p����D-��r7FH|^�~L"m�[:d?�*�6+���c�gVE��R��\(bzZm�� �9¢b/)�.��
���!�_މBi�?�}͢�3�T��1�r=d��I�H;��f\KjV���$�%����& ��� p+�����?�����u��1� |��A*�
�.U&_Ff[�Ks9���N9����v.����-�]<��v�{���ȩ�-Fm�Jɽ7����T�,��5�"�����Cɠ2�gP�>��8IR6�t��.O�&`�Mr6����>�P*�A�2vn�``X:�g���F���s�j��+�$H��U׬v��)<x�%��,�{�-���A���h�&S��hZ'<W �E�*'�F�*�A¼7'{0�3&Ӈ�?��ƛ�#h���U�N�:�?�p������z��Mm��q)_��ދ溂\��KZ�ϊ�� 1��2�X�f$��C�2iO!ų�W�Oȯ�*o�hz1��-[ᔹ&y����=t�c��R}ŀ±s�<;O�k`�i��f8�8� 3QE�9$vB45,�?�2}���;z���v��C*�|�"���B�hI�y{l�N2����x��1�#vBr��%U�L�6�^ �n���L��7��=�h	C5o�I�{��^�`�F�Ul*Ҷ"�)��|TT�k�p�#L��[m�ܚ�N9�&h��+AO��L/�y�;k�<om(9ؤ�(�C��5�D�1���c�����P.�ـf��dj��V�#2�m�-���9����@��ly��G;���4�X6�xtj��3hN3� T6�5_��ych�13���7��Cu��.o��f�����n&rW�e ���Kܡ���c��o���������C��|L�z�.�s�8�UGG�Ɩ´jn6�Q�&ެ�g>�Kf["u������9��l!:`�Ck�kw�)�6�uT�r� 	�^&Pݫٵ���7�G�
�[���[&�Q܌���s7�"���W��+�\�����)�����5��?��0�EC�[x\���&0���N�V�)�j)���/�{�@.��ʒ��`�K����m�4��к
���X�-{�(�5��p3��hd�!b4�S9|C�� �N��_�� ����-#��p��9�XP�u�1.���x$C���e;[�T*4�Ȝ|�:� �^����D�a���4Y�z��GRb�&��CF��Z�a��}�Pr�z�K+���,L]-W��RX'{��oa����6���U�}b��}Ӕ�+g!?)�I��@��U�G��q<$�͌ݢGC��!Blc�<���8�� �����19�|�a\~��\��*Ya5��w��Pi#hu��;H�m'Q�G��&�Ok&��o ]�������wU�p�����,�/j����F���1�Ym��\�����u|3R�U��ўG�
}�a��8\v�.�[:��sJ�`��a`a/(��o�����z)ML�!�~/OQɬ:���O����\v5��'t�\N���e�����|��)(h��~�9�y�	��m��!�n��ڝ=��4G�F��J����Y�\6P������ؚ��ȏ�D��� �(�wu(`X4��7�O!���'%'�?C�c�y��B
�Hc�q8�Ę8��.N�H�����
������J��3ψ3O��@����^����<6��ˡ��(����XT^�0�!r(��0E�M(!x܅�+�' ��&�.�W$V�3��zY�f~�}n�a]mi������\Dy�pw�qLֱ�e9�H�W���5���A�c%����.}���@�I��K�=7�z�Fud1
13�)
2\��	i[������+>�I�~�	���l���H�G� �I�u�*�*-2�r��$�YB[DS�-��֒�e	�wVTX�����n���%��m�d�2��HK�>�\����DF��]�0z����7>:��n�K��|��V*r�i�Jtp���
Vm��j���!�,��J�rXI�����4�"�DJ��Ϣ�>Ph���ҡZ��M��#�N�{��(?[>_ �R0��lUx*�m�>�;�[���r�,�@b�k��>ʘ� �,�/B
�=��">JLa�O�<SuQ>]�y��H���
���@��G�%��)1u�C�ԍxzc��X�s݋�K���R[A��[�y\u�:Czc��B�A��~��.i�p +2k����i4N��^�T��?:�R$��H��J�0�$9�4�?��]i�zі�/m���.Mݵ�>�]d�����,'7[�,A�@�Yi�7��I�'�����Ϡm`�:���6�'k6��`�&�
��kQ��L�:��!ąF���{�zew��+���7���B�66�uh~�~�-��,�j,�G{��|�������>�r\X�]�5��h�w=�I�]Y�ki���GX����ῶi�%�ճ����{��6 ]n�w����NIߟ��zVHAo�c�j�4�KO�*U��*=bJ1�Ά���pE̽.��OA�n#�� >#��� ��vO4����z�8��ܫʷa%a$�8�\�,�A�8�Q���Sί���ɳ�d��jc���\jC�o�!�?��E��ٸ�օ?��O��Gbg���:H�Y�>.������B��~`�1W��@,�;���H\¦����o�	�w=t�T6�-���j�4����U�M��F�v�K�!�&H6�>5n�!~L-�;"JN����ƣ���#�-s&1�Ȇu�`��;����HI��^7���t�Δ�5>�k�cwo|ed��EL�
�,����S��
�=ħd+R&���p3ՙ �)��1;d�t>Uo ��=R��B�2�I~FKVQ�4l�Ւ;��7�,�x�9�S	�K�w}krB�H) u44K��T̾����;�-�ƥkósƜxE�_x�tM����p�/:t��V�,�������t?�a��|��g���0W��S�s#��O�v�����Uf�7�4aT�#������a2���z�iV���w���u�ڻ���ĐC��F���_�n��8Hپ~ÿc��K�͚1�cG�$-0�,��yX�� x���ͫ0Q�6ߥ�q�����ѻa�d�R���:c1�H[I�)Zo�'O:n�Ts1o͇Lu�PD��plu2%�&k|70m��V5�LrU��`����դ����[X�n!��{���W���9�:���U{'��}�4��b")�� �T�rYY�s4��%>r[e�
�x�jg��!1�k��: �>�����S�K�%,��dw���~7�h��"×�R��P	8��׭N���Z�)�n��� �'�%3�����%μ���%?�"=�f���LLS�� ]�T�W�:�(�U�(�tx�U��pC�]�s|�����]d~�vB�X���HM�<Y�#�r�c_�<w���B�����+��C��!(�c��o�
�����i���x�/�#���2׽;gvH�}��e.J��T�eE7�� ..�bx�h�e��bZ����1�%���܀��g�K`�owv��cVyʔ����iN{l��-qO6.V0J�Z����֝�
�#�$�XȪ�[bܨ�ٕ����z	_N���B��n���ͷ��J���l�j�2&{�z��)v��'��˿��tL����3�Q���Δ�]�|��9\b&c�d���+Lxw�%_B�d�g}*�D��Oq)�Ȏ�/�r�/��_�4�ڞǝ��f̮$��S�tj�"=�Z%�E#�/�.��a�m����،i@rv����w��5_եb=�ʶǂ_Ď�J�vh�?Q!��3ږ�2�~�9w5{�_�\��/��\�\]T����rj���X����Ӓ�І��lnI������o��E_q gJ�[5C
���ũ��R�~����_t��.37|�5����݄��K����9]��!<_��xR��
��DHK0��=��D\á�Gb�M5z{�?�g3����@�o��I'���%dOoH�b�Ljpv.�@�Rl�#gf �ȌY�>ԉ�9���H�hZ�P'K�t���V�UD�ӊGB���~�HI\�S\��OE�L�
֓/d(h0��N̓?s�B�7���֚�-I��������j�sRq���� 7r@A���~�ѲMw��{�Z���z�S!J���2��?��w�VKcE���b��t��묖.�~� ��]0o#굆�oR�As ����
񁤹E��$R�ԩrl�����=�8�*�N�\T�1��eK���ih�odGy�F�i�VĠ��,�%����F�o0����Pm$y=|n��W��&�B͚��#3�έ;e2:��=�W�AĚ���l�0�P	���#@fTvc�o�$1����;�jѩ�EJ���o4�E�*6n����G�������Kq��b�
D�� �~\	y���+D8q��g���q��j��������U-r�j�����z �98	��P��12�Z�/S˿�uƎfR����%|%�>3�PL�	���#-G�^(X
�k�2��ϱ̴p ���+�L��!2_?�N
��^�z� ��;�MSE���!#��2[/3Ct	��u�������0E�j�K?l�,F٭iq2 ��;,<aIFrOb"ʔ�łb��9�ɳcj�a�| �~��k���☭�k�T��9��駽","h)eCv��YI�u�Q��1b��]�	��=�D@����eW��{ƪ\R����'�{QM䈜9ȫErr�= T ��(�?֦�Lo��^�8ttY
 F/;���
���d֠����
�eM��sLc�_=?k�S[��!P�50F'#p�d]]�H�Je^e�mq�K3kѼk5�OB2
���|)����\�R}c\aC��$|�AN@]�j�����rq�~�J`�"�-_/4�9fAz����8��\���J�h!2Rۛ�3����W%,�"����N@��e4|�2Үi�lR6�"y�w���ڣ������y���Oy�mo��|��������i��m�/�/�V�Z>3�����ݴ�����.��U ���|H������=4�!�
�F��������Ӆ6t��H�����'H���d/�����q�Z�o�A����aT��Gz��\f���؈TeKz���ȃ�}k�n���r��xy�ON�ҧ��˻(�W_4qkċq1�U!<�u�� �˧yI�ŧv�9_�Շk�1�����~r0�>	<����ﱶ��!~joY���'b��u߃㺄B��~䯖F�if�ȮvLj�g�P%G��+/�A����6:�t�n�+����i\�lB5���G���S�޻D]5��ߕ�Tϭh����DQ�]�87";p��5�$h'��M�����ߠ��-c#~��wG�fD}��)J揧�E�+*��_�-k���5�,o��}g�~"�����1)����������@�2w��˵��ŭ/�R��m�.9��7�洈����(y{@�I��Y�k%��St���:�����0��c�=����"�ϦYEWPڶlFwx�g�_��n<�K��%�Y~�.�	S�@n���(4.VA��
�<�V�a�/yC.J���\��ֵ�]�
Y��:- �y=���l�-�X)I��ĚtЇ�LR9TZۼ8|�@�o�� ?r�aj�����{�9)�r��=ȗ���`��lp%M|��`\�j1��	���X�ϭ.�+��ѽ�]-�^����p	�C�ᰥ��hQ�YWo�&�1pq��n��W��,}���/��P��|Z��s���������q�<t"��n	�7G	�3O��D��o�6�7�(g�m��g���j�c���|^ϠH��K=�B�":f�*ZĲ�v����Is#~M8I
3s�r�*+�2A`�Iz���3c���{"3=���+4ż�6(S�5�g�ӻ�ל��:-}�qm�?%��O� +���E ��Ù�Ī�;�bƣq�%�O�s��ƙ&�).�������#E�>��E�>rI��2��c��ĥqs�'Q���!Խt�Q`�f�t�9�
����S�_�7\�'龕�Y�G ?X2!�ڶ��uPO,�K:��V!�"�.�8��}�,BKs������qUK	��"�����q�Z��X '6-����	ϖR�3i����'��h�T{7ʋL�c,�#%CfD�b�s������(����<�-��G��w���Ґ¸�����9�A��*��������ARD�U'���}�Zb���m�L��i�c��}`���|�D7.J�u~�'��5���;�F�͝�����.�}��	�/3VIO��Ϛ���f���&�����oXD� ��ӷ���@0�����7n�L�Q�Bh<�k��h56bVR1��_�w��ςz��fN�-��� �:����\������H�����MA�_�׬����%�%Ag&M��h�;l��7�.΢��;�Jş�m3 �-u��7&cv[��ӟ/�^E��	;�����:݌��"�z�y��Bc�mX��u$t%7����=�p�c#"}���1V�����\[��X1�,����;���
��]M��c��/�Y@F�^� "�VsiC�gF4I'7�F��~]` ��q=
d���a���Dԫ�s��Q�q��OL��!�I  �.0����a�O��轂d�	-&�($�O'��	l�L�Σ~�&�I��3id���Ϡ�$̪+�T�M)��q,�o**��'�� 5!n���&c9c-PRKy��L`v�s����.J�^���eվ�^��U�Y�L,8_5���n&TynIh�͟p8ٔ) W���n@�I5�Nǿ��w�/e1O�BM�oޖ�ר{�?�A	f���|�<W���)2�q���F���Re���LU&>�[��H +
���?��k�֠~P��J��,[�6G���>���*5����N�1E3V�h.���3�����G�Q�vk���&��`w����? ��#H�g��f߲e�)��0��u� ؘ1N��$Y��ݿ*CA� X����{zm�������S>t^�zAU�{O�R�gh�O��d�[����1�-hx�_���0?d�D$ӽ8��=����g��3^WB �C�c���O��|H7���k�[�X�� aSȈ3D��Rc�d�ͤ���73�3
h5���f��B��${ݬ��j{�T� �lQ(�Z�&>��搐�����6�5�#�9� 8&[�#�'�R�X�J�B�so·�}r�k7���e��5i��?3�l�@�J���A����c��t{â� /���R`�.��v������$���F��0�,0�=��Ea�h���g�^��	�?��Ӷ*��s�W��l���#��F���	߫ϡ��I��.`�Y�5T���±f�̠��Ə ��C��-��eT�Y�>����Q�\�r��ao���VX���y��i؇v�B���fc�A��(]��V��-�[�kɕ���ɛ�8ac�
BW�"��8@�#G߶�����r�����)?DQ�a�=�'�BorK�Q��T�%Ip`�x#*�n8�|�{o<�Ao@ŏj�,W'�#��(3�E'�a��%<y���OO�Y�#�%�'�&{�I¾�$=���l�n����?����9���k��26����'g���G�Ȭ�~~��U�����.\٘�������s~��|�đ��~���/k4��i�I�IE��:w��h�xI.'��r��KܱLx>��|I��`�e�	�ϰ�[��xB(E�E��߆-ć���ʪoy1`!t��K,�_�24E��V������+��0�����ҧ�`X7B�Ѝ�r_K�ᔆ@��ӪY���~W��ޣ"\uNRNQ�Gഞ���p)�ņ�A� 2�&ܼ&��05�����w�?�3�_���-��w�Y���E��&b�Z'x���mȑN!54ʤ��k��W��6�B�� �7H?6������n`Vq�m��Ғ�+���<*Ayjc����Fm����'_U׳��!V2�ũ��w�o%GÀ*-�Mn�T��0K� �i��S�6ك�f��2p)��־~�e�`���V:T��+p�����:R�&)����\���f7��������Y4���%U���x�)ݷwPr�y�u��"��� 6�)e��t�b܆�OF>�+����Ü���h �����7�u���B��uWC�ǀ0?�C��q�N�&W잼����Sq�W}�|K����ٿ}�&�Hn#� �#�𬪕�'�[��b�xZ�Yc(j)F����̝E(pɦ`	�@�m}��@��s��W�η�hG��X�iq���S(j�aT���C��V�Լ�mv���(px�e�	#��S[�Q�A6�W�������i�%-�ēR�#>1�/���'��/��׆<�(!�;�D~���?��<eW��̖��>���HmG�o�Hm���m5�dE��,{�e������̡)�$������[��̀;(�$�
{7B[���=rx���R7��#��E���TV:�`��¸��bR�{h{dr��4���
�6U2{ٯCM���/����g9�	1�rQ�
��u٬�3��T^`
��Q.\��z����K9[���m��|u�Yn+�20�l
H���	�&�{A�:��	��yf��(acaMn�(�VTt�׳�
�s�>�۱�'�S���8�Ly�J���m=�|�8qd;���m	 ȉ��h�9ᒁcBRx�0�v���3HZ�����Q��m����a�\����L+=�ҋ&B�|�!l��CpJ���7D9�,��O�=��NIw-.�]R-�h��b�W�~����^�\��@8�0�ɊS��v"a��53�2ӂ=���Uyu
�P*���xvv�fm�l�!ﴽ9�+��f���`�g}u20��r�ݦ�:�@���0�S�J�#Ӥ۾UNwN!]n5A>�RF��H��M��5�ae��H1X�f7�?ZF�M�ڬ;���"�O����S6غ^����d�����֛c�_Tj���5�� �e	8���t��B�K�)�/A�Fg���t�/!��7|���M��*~/Y�J�,2��E�qNA�v>m�̇���S�`F�����6�)��ͧ�&����r׿39��<#�dxCҚ���?�Fz6��N���@�TЁ�Z��N�lU��_�M]	�ۆZ��]P=�<�Q�l+!���߭Z"[V3̴�y��%�{��ӯ	�PNy�u7�2<��Yv��+��)GW_O9�3Rҵs[eU7�jK�$|�ؘ��GZ����[�Q�����s�rWzQ�������Hbi_�?�/��ّhx:�H��!u�⌡�}6.X!Ë�bz���p����L�1J�]�1�i<�[F���QC�bc{��6=c�R�3U����3c�jÖ|�o���~wC�;Y��o�!��
U'k�|B���6R@b����4Qk�ƪ���dWo��ܺ���"�1�z�Nܘ����Gv����BJ���s���E�'�&�L�]cL�ݛ=����7ō���T����q:���RR��:�j_��;q����JJb�oٱ��%R��j��8"�*�I�P�Yi�w��|�P���KZ�k�1�{��~en��d��?R�9�.�|h]�d���_�0���- �U��l�)������u1k�}"�����{��1��X���g���w�]�#vk|�|͙��Olz7���D�Ƅ�bl����gV�k�p��Rk���^m_�<cGG�X�p�R����1-�w�e��D4�V�*+�1�Τ�=kf<���S��i��;���:���� �i��e�S�I[��l�)NA���I5���J�.��]��� ���Z֨�d�v�Ӳ`�@�k��7��=��B甋��]��1��!��e�����wS��VuP'#�'���5�'���.+��'��4�f��{OM�����'�Yc=��7/�Zc�JQ6^�a8�co9j1����g{A��r��Jj���Zv! �yǮ'^��ǿ�?|ps�>��`�TH}Jz��G]�/Ա�W���!X��1�^(B��/aN�y��,�-�;�z�L�R�90sOr�s��!0��A����X��R�w��V�z����������ȷ\m��1�\ږ�L�������s2��n��-����q=1a����e�px�~�l��L�� �"���J$�Ou�y�yvM5S'���fj4���.�����y��U�G�X�M�^f=fmK�`���9��>�$i�]`�w��.�I?	@�-YR����Xvgh�_���t������.߈�	RB.���לSٵ��г�w��F>�Z7t�r³�`[zep��?�ty&a���	�N{�D�@���fk��n�`�-�S>��N�fKcA�\{��glI�w��:߆R%�H�WK0�vw/uL�:����5qD�/� @/$"������U��+_�ᣐ�oQ�3Rp,� ������w
j���j��֠��&�d.C���� b��pƴM�g�J(�@�1�O4w�Ftl�quL,�=2��TXgĤ w_S_�yg���Ttk���D�5'����L!�<�/m�Nh�4��9�)p"d�.�;��f�?ŭ~WC���o-Bg��{�&��冥��tm�����#��B��/G���;ʩ�O�M$f�2�3���ݲ��j�8N�@�%�s�Y|W<q�����a��g
��t�)|�h�󚚍b�77v�|��%�0M�P�OB7`��z�%tꄬGA*�
�C�#������Y�_��³��$�����<֜$Ax�B%�a����#>`�GӠ������d���}c6�^�0�v�dl��#�&�09 ���zǐǪ�]��m�/}������Y��b�Rʻ'���V�f0��J�;:E=��
�gvN_��^�Q8ӠOT����W��ۇ+�e��򏡡������[�G�K��5G���0"&VƵ�Ϲ�t��A|�a<o��ћ]l� ���"��U]yaW%�[<G]�nO�+Y�PH*7�9�����\S��I��I�7�{�����W�ֲ��ޗ�')�i��1Iw%�b9BɴOZ���);�eq����#�-S�,V���.���)�����7O����f�u>���@È<j��bW+&y� �ļ����h�����)�FZ��Y;���ڇ�4Ѹ(��@�&���IZ1�x�8Rz�Y�W�D�v�K]�N����=��c
D�kF)�&sV	c|B+��{�Z����ĊˌO�����!�2̠�0�
y����=%UߺqG��>}q�9�"b�0F�Ⱦ`pS�C	O\�����=��c�N �� Jҷ!�4��)G�m��y���mڋ�
��UaW���K#�&~&��.��t�tJ��]��VL���M��[�N��~���%7���շľ����.2`�·��&gqb��u�9�����1�r�߆���0����u߰%KE��P�p=sb�����t>r��cJ��0dH����"�h�,�9?مh��6��f��4�E���Ձ��E-{�q�5�UQI����yTT?�y�T��N+h�B�v/���z���׽T1EQ��̥�˯*ѵ|�3�$`���+�sN7_�4�d�L`��֜�`0�A�#k�l zQ��O��C��i��ܙצ!8?@�1"޺�+[a/�Sf�xyܗl��E�G��/z���{�����w�%���L�;$&����O���K�� �A�n��5 �S76����.vQR�,c6&�wn��͉�}��ſ�^�j�b�H�q�샞ZNl����{���!h!����Q���n,\�ȋ���	u�>S�a8���임w�&��y�>8���ڐ!mj	z��X'� C�&s���h��+�Õ�@�)�+Pק!��.<�ѣu7�?���=˜���C���҂�"a1@*[�In܅�ê%SJ�X��fP�,��P#�Ux���V���w�������m)�7)p�۔)���xJ��;��dTto2�o�j'���9�ǍI����������d���u-��Z��J��*����ۏ.R�Y�G�O��8�{�-�ߓ'�{Q�,��闾��\$NS���E���f�Q
��Y`KI�@�+��Y�r��G\Ĉ0��鍅�gOI�1IM����U�I�#hZV�K��)K�ql��� �M����E�&��<j�蝥X�n�{�S�O���	H���m>��n$�W������u�w����	�j_�����@�K��U4h�M)ᵨ�w/���T���Q����b�h��4�&�Y�F��� "�Ҷ41G+y$6���"YAt˵�ևK"F���#��'���
���H�|�IT��\��JBe��.����i�����2�Fk�7�a!��7����7r.Q٠G�5w�e�="����C�M���hDB*:k��*ҡq�<刳�k�����^�
a�B�=��M�7������]�)Y{�Ǥ]�=T"&�����_�@���e�+�4�wU�ˊ]x7pzH{a��h�� y�ͽ�������Ǐ��eTf���I�����ɨI�M��K;}o�� V�4[g)�A�#����m;H��ޅ�H,㉏b4��V��8�9���x���Uue��r���h�q�}xpT�L=����O���7KH�'�&D�k�_A���@�Ǚ��b����ѭ��(��!.(Z��4���fXS�#C��W�	�jp�s}�a7�y L:3쟬�[?�`ĸ/��;9�Zw��'����r=�g�uo�X�	�;Џ�5a���X$�o!
c�Q��l�@u{�69n�^����`򲴞n1s 5�~ܢ�R�}����tP�|�e�#����o�+����n� �KP���}"���N�ja�U�k�^����](��@��G�s7/�޴S��*N�TU�f���6�ث�Ri_i{p,`^�m�j= �5,�n���V�z��`y~�Մ�X�/��}��A���E�^��T�����p�Oh��J�Ia`E����[�`ƴ���:v=o��Zj�zK�36uAVRy�x[TUe$�j[�O��	�2$�����V���vj��z�-�90�/�h���B�s�0��o�1�
��A��^����I��g���JlƬ@`[��[?�&-��ĥ�yZC���g�!�^3s_��9�tx=��"ue`rǶs�.�ܵ�|I��nY;vc16\l=W/Æ����TK��'R�S9��N�������RE���,�nh�����vQ�����r �V]�4j�|��D{��`�PIя�����tF����S�w��o�u��{�	��ړt��S3B���m�U�ݑ�ZQK�_ŏj��QB�o]��:��y�A� 5�+����;�ܣ�%�ͱ\��Pkze�@i����M���D���u��y�! �h��.l�b`��%3����l���W�����MBʼ�ܺ"�����V�5���a�%��� ����JE?��#��ɋ&n�7��r<ph2F��wWg�y5:m��RZ]�:K�����8v>a�M����k3�l�5�����VȘ��yc���=�a��cc�$�b0r\���y�� ��ā�]����� ���������JY?n���U�����3+&�v���u"�!AL+����[,��|h?���f 	���r���x5�+�s��lC�lBU2�g3��|�4A�*o���g��]���&ȣO#���C�CS@=4�c�A����򛻇�W�����K����)[�k/?+i��455c`}���S���K�`F%�b���V�{�\��*{�Q�����ñG�	Q�2�Y!�0�����]^%+םvbZd$C0_�jx�>��c���s�s�L��lE�n���������q��Vs�cer��|T�
�l�!�^����P�y.g'#�g�5�`�Ds½��M�0H�sQi8�l��@pUOlɒ��:�����C-f�w�w�M����%+-���N�o�k�(-�WIS4Q:֠�Nw��U���E���U����fF̞�^�]{l�����$�!��,d�����	�z�Z��KA�ܺ��R:а	tj_�eI��4�I�Y�SR����u���T�n���U�_�R�|M�#u���_���Ϊ���s��F��B�����6�<�Ɖ�&J(�g@��2r�cĭ�h�Z.Bo���zvP���IhQ=`b8g�	Tli��=e��L���:`@��?�]D���&��Yح�.*��b>"XR�� �F�c��"ǣ=Xu���g�����v��G?.��u����w��c�_|:��υc�	��)�)G`t�뵮Q!W&�!���y�%�v�]���!�מ�H|�k��%?��ѧg��ț^9�oZ�����W����Z��y��
x�\��r{�3�Y`8�A�(�RV�ɴ_J*BuҸ	�s+=����ƪeU/�m{;�4��k�]�E�B��cF����n���NSC��Dk�1�vM3�5��]%Apͯ�1�Ξ�e�������,rAqr�2�?���b�<��̀R[�]Z>�uԟ+z:� .��S4�����+�̛=����T��62TJi�9p����YSqN�:Zki�y'�|%l�׺{�^ �,����R��c�=���Pİ�;��("�:��\���hp_���5Ƣ��V/J��Zf[�+�{�T��D����N����L_7:/�6�6p���1�BVq��@�sB�_!�]h'@aF���^�C(5�#D�pLw�)�N]��AU�Q1��,'j�J[q��;�Q�Oa(�`n�ᇣ]��9��l�	0Lr���q*H�x��q͸�vm������7�hv��+2�4�=��-e��?�-ϩʨ �:���ܺ�/��E;�� �k}��=}�O�W��>{�(���_N�\K��pF���
��⿴��g�.�ƀ:�[7i�r[��k�;��j�M�= ��A��I�`�e�J��'�qwLG;�530w�� ]"���B��8��!��5�H���m��3܉Ch��nx�@?�8.O�Չ
Zt�'d|D�[��Z��F{(�t�-DS��9�ʝ����g����!!4I4���:SX���O�������]�SIJ~{��0_Q��D7$�}��49�Rz��bGo��L���0_�$f�7� �~Vч�����
��7$e=�K�A*_|D��	Kf�P"I�N�v��p�P)��ho/i��V��S�����!�fTY�C<$� Dԇx-�(į����X���MK5�����nE��Ҋ����N�i������4�J?f����މ!j�QQE@�ڞ�G���q
�=��&���ఱ��-x#b@ו�f�yB'(�\��e�v{�?�iY������\lm��Pp8�Ka�@��ץ բ�&)��Q�~CF_	y��,=�����;�Y�q���;�e��_ω��*ݙk�E9�;�w"�!�!��Z��Ķ+���E�2������[К�j%���:��_�d��Oǃ��'�(����aҘֱ�TQ�hpr�����)z�]i� �'sN�S@Z�	�s7�<�MޣAwj�s$ɢ�E�C�/z���л��U�;�V@�F	?dcV���u�����0_�f�Ѕ&&݃�t�C��V��ح�q� Ow7<����##����,�<�.p}�����>ctG��	��y *�����*��&EI���J�Ԯ樬���E0�ˮ�o��Ά�1�}�����剝���棤���^�q�f��灱[�/�����F�(�k{pB�V���HyeƓ	�������v�JЃ�T�N�=lꋬ�{:��%���D~Zz5>� ^sPP@��s�<VMfZ����2�Oa����������W���/�A��C� ��5� �ܵ�~������ʮ��օy��k4�F�T��G�I��<�0u�	����Gl\�~�2��8�����r�0�Sai���~�"A�8K��u�F�)X�5�L:��J��d.W��zsxy0~��Ε����2���D��q�s���,"���9�%�Ek�ʭX�yg�sh�-�&�����O"b�psҙ�_Q�rc~���R����K�]ԣ��>�a����!xP�v���k�es�9Gڀ"x���/����!ċ�V����NC���/�����tkf!w�d�A�i<E�9U��X��6$��
�q��)�N�漍��LM4X\餢��檄[��`�`!�n�
��+�ڰ�MIt�Z�Y�5�3�ۗ=PB}�3(	����#N��Q�ە!��,{5M)�O��]�`B9P����v߹bE�c�����Y�$/�}r�K����Eb���@��*���G��s���ymj�.�w���
�Ζ���Q�A�S"t�H�0>C��E/�]��N�is���a�;�:'ƶnN�Zo	=8�VO+���Q�J-�ͯr��������S�-·b��j#���ф��n1h��ɥ��?�je�x����o�d���gn��U��=dҼ����,�$D����7��k$\��������r@2l2��U\n�|}�\�ͽs'�l���جic��\y颣�*�Ʌ���D�P{�x��S�&�4Qj
s@�క��}�e�E����d�	g��I��N��Sab�ͤ���=u���j�+јQ* �/m�g�!1VSn�|�x�@�bڞ^K���Bk��^HhX3�����|r�(? ��iHH�̩��b�E���X��a�
��ݔ��{��dr6l;�jI�^$�_H(�Ϫ|o�'��B�q� �*:}�ܕEi������!����[���]&�F���c}��&�����mV��b�w���<��MAd��t�
-SJ�����p_��<vn����]�/���Je[��26	���D$R��}�����5���s�R�K����a�59��9v?
*�%dy���x���6؞%���g"���G��l8���`�t��W�[�#�;��e.ew0��%������nSgHBE�lĢ�(���/�&��3���x^(g��UU�5�(͡��a��g�S/�f�%-��5]f#L�B>i���U,�*0H>J��r��{�xy��B����!�ķ���̥!ڇ�:�*����;�����F��{���Y��pο^�ߏ���-@�|��v����4/8���}�7��`Ǖ�����{��#�@�:�+ ����������/�w�#=6�/5�� ���	JM��~�z@/�~�=���[���{l��c܌d\y4�X <�Y�<.)*o��Q
�:�6�!W�Az�C>Se���D,-��O�Hw���'@Q�.8�1�Ø��"���������0����¦�e���H$�h1�?�1Ȉ�ap���&�@I��D�K-���Ԟ�B2��9�Y�r��>��ڭ;Q��=a`��@E��EW������v�~�9���]a�y�a��z'����8��u��f�ۜ��ފ��;��x+*����SmߧH*w���ר��v*G�j�18(5���.V��F��梶 !�Y����-icD(�*���>��~H��4���ٖGN�#=i�;�&�þ#�h���+#�r��f��ɴ��x-ê�٠{��9�;\������ą[�9����i�7C�X(I���M2�cn�ޠ2�KҾ�
�Y&���2������$�������,�d��0`�_��� e���ϻ���>5k�h�C�3�nH%�o���X��0B�������w���nM��E�I+s	��)��$��k,eGt}��Ɗ���`1K��_ݕRF�c�c�������C%����Qٟ����F(���v���p��2( U��~I�JjA��I���H���]��&��Q9�n��?����}��-zHo���'�~�1e���������$��Y��o��6���h��e�!!p��(�~(�T��믒�'
F���Y}`������0�̜�J�.�B�q����#��X�tmy���d�D�~�s��,����
w�*�:pt^d62��܀�\(J#t�J��䙗�]�&��8ݫ�m����ۡ
�N�<S]B�~�(�^�z��� b>�ž	'g�}���5�(Y����w's��!�a�yq��B��sB/����bHdw��i��2S��Q�K�V.�H�M�A ��;Q��y�5��ޏ�g��]M҆�6%����O!-��]��"�4m^�fg6��2�*�����f���d<w�Q�+6_r����"�u6���m�%*BE�����q}�좆�	_���dO���fv<�2�C�1�87������JxH1�U�n]��CQ�H9o���S��94�	qE!��W�08 t�^]�ïTI�|��t'�z�~H�i�h�̠=� �e0�_ݻ�I���^幧�i8�z5�5�L���z��H�zֹ]l���Y֩�Ն��l+ʵ��L`�ԯ��dA�EJ�{��UM;kx��Q�\�V�,kq�tf���M����Eģ˲���J�7x��y˓��j��m^����^J����u�FM�M�Y�Pӣ��(�<���%������[}Y�B�/׊�a�LvΙ�m�f3����?ԑ�M�����V�@��3Yz��<1��C�XI:�y��/I�p����]�%B�|$���v��,�^���~�1 �1�n��j͂���1ZytT8�����)�ˡ\�.Հ���H��Esx�Iφ�������6²l��*i�{T�����u�X�(�dX���#3�� Xe�d{���]��ok�����K�Z�t��Mf}?�&��ځP����QU�����l��*���]�/)��r%�|�j��ZAÙ֝?C��P>DZ)�ﴓ�r��E�r�]�FЛ���aݯ`�$V��|G���E���ף#Q�2� �4=�x�%|$��yo��uр�E꨼��k�:,����|�2u�e���;��>�uP�E��3�u�L�\�.S��R�!ћȂP�AΌ�	�4	�RY���o��Xߩ��Z4
M�`fU�l;_��AD�Z�٘�q�{dLXs/q���3����KxA�R{m�l�$%P$7�=�.�9��E��hZ��%�Fys�=��|x�i�BlB�$�[pP}|��Wڊ/��hu�>w,\c���:6�S3��:[�ٷ�l�	�p$`�(����\ר���l�n�'%����J#���?��JȠE&_%��(����Ï�Ҥ�/�׎g�Ċ�^�5�)}��|/)����^��1����ۙ@������tx7����v�"0��$�m僽�Qَ����d��F��%����+��8S5J���m�$��*�^H۵Z��i�ɛ:g5\���d����6�8�I�c���\:o��h�*֥?x���5n������oh7��%}a�'����qd�fk'������<P�|�a<=3oi��������釱�c�a4�&6�:�l	 ����;�J8~xɸ.�֨��������dA�.�Ç0%�E��ޞ�נ�'dbʫ�\Qk�����ʣb�Rێ.:��d�!L����> ����]7�I�r��&�LK�:z�V�2''A?6Ox����..4��I����>��F���]�[`��U���t���iL�a;"kEDĴ�˛6U�K��UMN|�e���ڕ*�kTF����@12�s��g��d���4�:�H���	ERX��Ap��5}�ૈ��+Y�N�w�
���c���C���q�is6�;�%����}��&N\fE�CTY|��9�5Q�2���� ^��m�C��qJ��4���j�8�Ü,E=z��<.H�����n���pT܆t�O���.�����tZ4g!.�Xm�~��'��|�r u��ZO	KC��ɋ�e�G�a�vř�~N򕍜�_f����GM����8My��c=
���i ��@�O�X�~���"�u����x᭧f�T����8���G��&m4m	�|b����w�	�Bf<��&���YA�������H�ѯx�a����g�e���N�%8}���^l[��e�3�����  `�9#�͓:��x����{K��B�������"�&�q&���jf���j�0cwįpKՉ��K���{`	��ಠ5�|�.�5N�B�x>�8��x	���^���5������ݛ~���C�C?.4�8�[Ql�D;ۈ<�M15W��������]�r��'`@	�&i�1C�<X�zٰ��$�0Z���c�q���%9�ZF�%�M����J�ߴ:�}�,���ƤzNO\�ޯKT��D���	I�I-g���h9зG�b���!����2M3�2#g[?��ٟ���aK�g��T!N3v�4}&��p��\�~Ѓ���,4��`z�E7�A�20�L��>�N0AN��Ci����J8Z���B$�t/~m&l�6g��:b*4O��PP�GY�Ϸ`����Aw�7$ח��d@qC�M]���6o�OQM)�~7?`�<<��։�����K��;���s�u�����Յ�V\M�h�W�8���{RA��B��d&2�^�.�0V��	,O������&N� ©\ftcU�S�w�멚�EtUm���xMT��F%ħ��)��% �CT����H$ 4�5?DY��|5�Uȹ�QZ��)j|�O|�����o�e��04_e�<����KǛR�>9eV-
&$��@p�(��?gG&����ȝB���{׹+�_Q:Y��D�x���Us9[�@���� �?w����s�<�?C�h�c�rS�MtGwx��&F�92%�-{�x��x� ��9����1���HD�[��K�.98מj.�����-�2�¨oqU�__v�P�����(�c�5B��=���\�z&�� b��w�s�6�i�8F��nr���R)���abo\'�e����i�txg7a���P2�v�'3(aũ�����b�L?�����%���A8?#��<�M��5(�t�k"�+���\��\ݙJq��wCh@��f]�/����r�Y��[Z����/��g������(��gN8��
���z��K]���X�����S��$�W=q�]�GQ�zQI�q��q�q��
��PTԹzܪ�{EƔWX�#�5�Ⴈ�o�:J!��f>(��Y��?���rg'��_��j�n2�����ƶd�z�䭈�m�_g7>7Ԛ���V�Yz�_&���;K,�,x�m�`��2�.h�#f?���0�������\V�H��|�Jo�����"�J��[�4��z��U�����xu�p��t�"����Ucۘ�@�xBq�OkN���� .����ڵ���׏q���g*e�b2��>^
j�S�O�������t(?CQ��C铍zڀ�R	Z��ew'�J��`e�=�;U2<%�m���a�촛�@���^�]��L��£W�v�.2z����X��Kłd0�w4k&�)�@<�|�9'���ͅ��J��DP�H)T�1sÀ�� T#�`�m]���AڠxR#[ �|�s(�On���'+U{qP2�sx-�|���~ߪ2�-�u�±R�[�4g0�0�"���@��-lIo[�HlF)�3v(���\sKA�ބKO/�.������˿*h\���vg�R*��Cj��7�ӻ��ǿ_��'r\�V�����4�Șa�y�A����O]P��Jp��yq����*�~<��n8���KZ�K�7�¦C:B��N��X6��7����9ɫ�,s�{��e)�f�8�Y�&ur�x綥�}.��c��й�s���N����Yd?��d�e�hw�H1T�H���p*�[m�����>�G~:jS|d�H�������xx��³��zm9{a"NP��N��r3��{<q�����aM��s��B}�ș<_*�C��k*MQݒ����$;�h} n(n�$�D�/a��ӯ��?~;SP�AK��?��;~�OQ�\$`�c'+��6���َ(~U�ѹa�z�x�����b!���v�~�%ы{�����?��y���s�m�ʨ.p�"�#</ѕ��{�V���K�7� ����s�N��G��o�q%&�,���dr!�!���KBx���K�M< ��)�J��y�D�7Qa����<pw���##�%*Pcx �[����m�^�0�y��?P)���.`�\�$�P��6{��o�,��2	<p�4z���������L������>�;�VE�>v6h�.n��,NL輰�)v"�&Wf�A�24��Xm[6�Ia�O�/T3{q�x,��q=>�q�3�Ҽm1_f>�1a:FHf/8Q��8��!B���F�� I�#�!JQ��J��@��sVN������%��-G�xS����ҍ�v���2vJ&񭑗�_���7�b0��`"+��C���,�ϼ�X�DX8;�A��/�d%U�����wmN�1�='c�?�B��_�p��/:���֬��Tۇ�[���L]U�DMW�I�o��_�
&�~���_�|�17g,�����T�D�s��!�Wṁ�61����{hO��O�_5�D֙��#�}�c﷞����>���cL|�����#�0�+��@�%`�R~j�Ofͽ`W<{�����A�	1?�_�t�MƜV��ۡ�m�xf$�M�)֑�I6!�H� ���³��QC�%���w�]n�
	�_�с����Ԇ�hIE@�+�K���;֟�����Oq(a�c-��צic݉t��f�Nź�8���O�2vlW�UI��Uw�ZW����|;3��֤�&�B'���A�>n��/�^��zI~�{Rw���ܨ������I.�F�V��#Lc�3��Y�Fk��|Ӎ7�K��v^#;:Os��Wu�ڄ����_u�=;��T�OhL��Թ���������o[� �":�_��4)�cV���M��WO�Ɗ��.T���f��_�q2R�g��5^t�^ҥ����JkG�>��r��0�0�Z�����D�eM$+��%�f܌�C�t������3�y���*חa"ݏ�)O��B��>}R.���,\͉�l
�@YQ��q�ܮ�|�T�1MLҖ�N �h7�hZ7�$Ta��`� ����>�6���,oR��/�'�dOt��I4�E`J��p�xU���V�VS&��t�1���~�-���w]�%�i�ч��|�v��(Qe����0'���v��t������<#�A���q"��m���{�Nw&��O?Ȥ�ښ��ǟy�,O�G1��i͜�Ý$�b.#z����HV1��k�\ɦ��)PlU�����WقT�c�w@M6Ӗ|xh���S=�� g���k��
��ЈH��u�����r�������'��)�a�9��H�7����`ax<�<��Y���\{�����8 �$�Ɋˋ��i}���\#�R�SwW������֦ⷹc��ZL�cQA��-���<+��.�}�@�=�V�~R�iS�"��Q��ջ��ya�~�.���I���7�ޘh���e��U�G�!�OnY��}{���kdÅ)�sÀN�o�jb*;�|osC�eB��|�f�(q��X��U��� .\	�*�ٔ;.�܂��Tu�&�BD`���s����'�BgX�uy&Nf=G���7"�ؘD=�u�t�n�W{ ���Ք�tB�s�4PU�:�(�����Wa2�';|}�.cʺ8,�MG�)Ӳc-̾���Zwa�B� CF�J���:��#PC���Np����<,��f�} ��4��G�*༇��H�|k�-�}l�a$?m��4pƘ"(
�A�x}��P��k�_8!��/�*̾�ZM��H�(ˆ!�y���E��"�:0�=i�՘7�������$xA9G��qB��=�0���b�"�=���Ff�`�l>�ᝈb���'٥�W���?K��:uH�t�q:���Cb�P�
�H��w�z��VՋ���N����X	I�2tK�g(``�|�I>p�~��wJ�s�0C�>��y5�}n'�X@3��޿#�a�� Ᏸ5�I�Hp�h`r�D&��(Kʳ��	�o�J?������q��\��>(������?���t�U�d�Rh�o��ۣ�V*
��QI^��4Ix�c�N�R>���'ݦ���u�D�\��h���Kg@QC't��X�oMBZ�D+�t� U��,�IX���o�-��	��e®�Kr�-{���%la��Si%�.���4��{7���$��~vK�Q�zcn7�1�m��g1S���;�⌖�,��z�v6G2�	?��Je��J��g}��0w�_�~_1�ڂ]5=s	i�!Tuj�>��/���XI�!�h#�{uqN|�o
,d�� 7��9���K\�p�>��4f���+w��,��ؠ�AG�X	�e�3t;>������/�w �of���n��kl�Li���vt_}���%���PE�C�h��H�n�5G��EE�F���wt.Ce�SyE �.0����^N���xB���,�V"���8 ���t��2���f�C($ud���fW�yFrgW^H�/�Ͻ�a]f�"�U��F.Ǯ�;O�dA�E�U:s�uFJ�{[�Q�5�P W](� ������� (�o��7���;� <�.��Sz�Am�[a@Iͻt�Xk�;m������u� C/U�s#D�6�u��l�X�re����0�4���a#��,��|5�<�*i-��p�ΰ�^(*�v�;׍,N��_W�L�ʞ3��[�m��7�2>�J RoV�Z����j��(|��U��,��^f�:���pˊi�Dɗ!S�[�����{iME��]�\1oHiּ8 �2e��8d�@��"�NdM��_� s�)�dܤ�L%�P�!K��ZB}R���?yP��Nlp��u�1�(�i�싍�i"���tI�-+SȴtR�y�K�M:������9q�x�'SߤƎ������GK�����#D���tɱH�1W@��:n5D�8��(Vf&�3+M��E�k����DTPV��ی��x8��BA27��jL)X����Zx�eHM�Ad��5����-<�Vu�Yv?'�`��-�Y� 
�Bb\�����)|�1�sD�
�

R�
���&���(�	g ����H6=ac�����~"��	y@J��=ȁ/\����f �� %T��D������BHtϳ�X�(`�-Fܢw�m�6���({�/<z��l>���7��ʡ���4�{��hȮ�sTF�K$�=)Emgu�!��;�L�7Ώ�����<������˩�n���FVY�i\������Z1D� )�ȌtNG�Q����Z��G���4Ԓ�ϏZ(J���G ߵ�+����k�\�I�k��ܪpT��R���gddG��O$2i ��{�Q�����J�Ҧ{�%܈Ay�ဥn�)�u���A.+$�=^SG9.�n�W1#|1v�`c69���$V�4���)z��bU�w�V�����e��lm=��mr?�~���>U�9�0��l�� ~��'hHQ����6�[��<������Z�O�Q:(�o�O�c�N��e/V�:1���(�CT��ݘ=����I"��aۋ�3l[P���P[�'��ͪ>�JO(����� �[M�9[�`^|%�X[(߀�N�;$�%o���8ʤ�[pW�,�8x��)�TŅ��5L�h �H�y9��~�LM�U�︕�+�zD�:m<�Q�0�˪�4��[��.Ɩ�%��n����n���#i�h����,���Y�E�U�����F( &�\�i�FB~�a)k�8oӳY�$p�g?��Ձ�^|�, g�L$ю>�E%"�}v@#<q�ɷ���R}���d<tg�	��y�L"(�Y�FijWK����A�g(�^4��n�~�9���S#g2�SY��KZ����iӵ�K�KCs��$+�Mj1���m-��#�s�0����(5mh��"('���3ᬖ�?\��8��0 ������B���|G_;R!v�����F�n� ��$�	�;L߰���jf�G��H�)7���w�v��y�������c�i��N�&ip��e].�ڧ/�@V��U�\j��\8�\#���)R>|��[j����h�8?+�t�X5 z��s|	* �E@���{����Q~�O�����%�-�/*�|��_˕�%���E�&��m�Nj�e���3I�'T��PzՅ>�c��|�����R9|��!B���Zh`!�a�$׸��Z!x�J?re;z=��.���K��q����M$~��b��l�y߈o��F������+�`�.���E�B��XC�䩄��@����y�F�חE/�d�5bn�i�@%�n@����a5r��Hο�D��׏����1P����
�,�ȃ�R�X��_ܢ�eS������Q����^���� I�5b"\���O�^�~�ǽ��d}պ*+�*�;� QX�c��0h���Q�)J�(w|�� D����ڼ��ԙ��4-8��b��}�{h1.�#�,�/E!,�*�k�}~Y(?t�V]�bN.��=|��+R�q���i�M���&5B2��؏]���vk��Q2��ژf��G���l��hu�?�I����C�Im�7<�������Ԟ�T�d��l�rh�� ���t��yd?i���S���Jv�����=��1�[L!���Z����x�I�f~?1`�&	F�X�:�U7r�Ė���)t�pf�:`�d��h�7����d�EG�`�*��0��PL���>p��	��Ca1���'8Ĥ4��<&5B?u����v�p�\�S"�u�NX1�;LXp\�fSPUӂ|�2�B�8����@Ҽ���J�$���;Me�3��<�b��D�a�]^�|�	d3P�B
��'���yn"�U�!��'���J�����-���>��H����~]ޟH�߳ݺ$N������%��v�6|��,8���J���o}��������0�z������{���+?�g7�[�6��S�)��]R�ϗ��"��Xkx]�r窱W9s3��`�����a_9��Q[��	�IV�Q,�g
Q�H����:��ى�h�U��+�U�f�i$���t�p�d� D�G�򁋭���-I�$e�?��<�#`�<��{�c����14O�<^B��t�s�e*���S\�qXG����U?ݓ���l�9���2��{C� L�Ʀc{r����\�h�K]�����[3����B{���b����"}f�v:%gl{l���D�/�ux�H�-�D���A�·o��:��Ks����#�����گI���sP�Dkl��ϓRH9���o�i iI�����f+�W�#N޶��[Wٽ��X�4W���^�Es
B�Z��kؼj]�JD.QfwT�7�QЦ�zڬ=t�ٹ�0����.��{Z����j�41L'#�Xj�pw�1��A��J�=c����,�^]�8����%^���۸5l[|���R�ŌM����{�F�洈6[�PU�}0^��Sdn@���ŻV�Z�X�0����G��C��{��%,���������JOq�V��gUY4��U@�z��(��'�ح?Vh�Vɉ���B��rptN4��	��O��ID��4C��;*ט���������rˑϠ�M��Bo
l����,�L����M�L�M�#���,}Uk�c��d\�,�;Z ���1Җϱ�9��Y/��,"��f+䦱�=��"m�C&8ΐc������wW�P��.�P��2<D��I��� شc�u#֬,�>�=9s�P��o֒R�6���z��sji���y�X�oq���/��>_ W؇���M�$�w�X(�?�_�;vo��0�2�����ܢ��\�;p%WƝŴ�"i�� 4T�u�UO���|�{ϬJ�tm���r�.��l���L�f4�������]�#���%�GO��␽-���4����� ���woNI%�D�k��)�g������(�����a�� J��5��l�����@e�����)Zj�n����q�|[w�>�>_3蹟����o{Ѐ}>𘴍��cE`*����ρ�>À������r�hxe�}+^iق.�V l�#��>�w�k��lj�DR��rs;���R
�,��䛡�ɔ��VBj��-æ0c�'�ÑJ\�Q����f�|=���eǳ�����8�b�PEڱ�߹P&v}������UFF��\�q�6X:2 �G�#1��uKIĔ0�~�uL%)�l
y�+@�F�'��%�: ��4�6B��V?7`�,Qߐ�b�ﯕ?�"�����	���L�{����6A/<]{(��PQ �T.9�Zf�uQNKL-�l��`��|wﲍ->[W컾�yL ��a���y���K'萫_��Y_��<i*�\�/9��bY��+��-V��g��譜ӭa����n?�Y�ݫr��U�Q<�N�Է��w��%�W����܋�B�"(n�(+$Rt%`�R��g���(�c��G�A*�}"j�?[�rY$OA��S7O���GlbJ��W�,'�"�ȅ��b������-xܜ6��AN^�0k,��[�D�_8�݇p�y��Q����.��RP���'� .U����:u�)�@�ih8`CH!��Z���׾'U�;�ꦜa�5�c�$���h��;x@�M���]�K��.�;H/d�6��O2�,�?�a��ӵ�J\	{o��X���u ,��鮞���
t�����l��F9*ׅh��P ���`d��5TNPRr�d !���F�:��a����4��e�|��a��R0F���fE9�[��Vm�^��{ӗ��Q��g��0�����46�
�׳�;�o�T�,E��q(�_l�Q�Έ���k�A�x�Mu��9sbSD�� ��}�&M$�bs������C������>��<�1�R�A������\�����+X�e��;���y��%��j����D���*ͼd�?A��r◹����a���hRYiU3�=�u��)R��2�(C)�ZD��{g����R�ذ��Ժ/5�ᘃ��e	�@c�=y䙯�&��p�x�y�p�J��M�����^��ko��b���Q�1H@p�3	�y�3;�8=�HL���(���dv0�g-��X�p�ˢ^�M/��)����8+�UKGs*�+�褃g��)���v8�����*!Ӵ�@|��G띹��j��Zj/���h�q��2N�V$j�k�O�uU��fǡ2���O��Ն:|��D��J�)U��r��J��R���W�M)�^)5! w}�K�CB�S�G)��� �� n�y(_@�;����Nݾ*O��?@;k�{NA��\B�^W#��Z�
A�V��A�`���[�>�
���e��woK(��!��&��ɰ�ߪ�M:6�ů����#	�b����	�E?�u:���"��'�g�ȇ�a4�$������a�O��9���)�i�%a/A�����\��|�*N�G%+���|�j
�
q��w�vTDu�y�0I�Ϣ�J��+$���F�6�)��$�KHOH������IWr�ׄ/���Ոj��.-���e�!m�	J���V:�Ա&A�7-��ĸ[G���=2O�fȎ��P�{���1)��}��n���G��Q7�{g�`J�.7LZ@�������fgdwKM��?��7�m��;��E����z�b�&��ČS^y��I���gs��{��"d��2����+�	��`�t��E���U��
�LE$�?���:��t�D�W�Ztozu����2�y.�{G�>���*�?��-��S��1@�͇f;��ĄIų)���j��$(�ђX����rԙ���������)�n��5�{�fr�z���Y�(�����V��� 4e��@|�=�=1�2�����=ʢ.��ӊ�xwe���ɜ��@Ïi�d��;�e[��\�;.3j6����M�hxZ�ՅzMf櫴`)�(���n@�-�K�e�U{�)$�Q�х��.H"�f��*i�ge�����~�l�Z	Ch���X%Ѓ�w����" �������Wm|�4�D�
�dJ�TQ����;F�d-�K�&;._G��J �<���c�Y�i`�g�k�i��@�''����d�������D+ba�������Y5R�uKw��(�j����rw�O��\%�����&��0�,bq�H��#�/y��E�+q�"^c��B\ժ�"0'�aw��ʄ��W�ɚ����.زDCA���c	v������1ГN��kof���Ƈ3�����2QpZ�i3Si��E�7��
��B��!󞉡�PKiz�2���f��|�}1��N�b?�.Y8 A��
���E���/�3�����!?�Ma��=��@�n��|�!��e�哂�j|�H��>$������������>�H���B��=�y?�����D��e�Cݎ�f�����Q�4%���S?� �+��VP@(�$��&R�ǈ��կfN�R�F� �8����V7!�qJ��[R�ã8��1��Z=]�>\�eĝ�+�0_n��~w���|k��U R&s�)��6�K9��t֖i\7�r�}���ǒ�> �]�&<^@E�.ʾ�Ń'��
��ڥw6#�'cc��;c�X^����YN�B׈��͝K]���#@'�g��*�!����Ќ��I�R
U>q4�b�J
�75��<[�ɎT�����P��v�q�����W���d)cX}�/<,"gO�{�X�@! H#�KI���t%�D�v�.hPKD�����_����0V�L�4n������ZTZ�sr��U�a\B̈}9��g�f��|�RL�@ՠޘ��N�&�������%8�2�d?d�nJrD���H��8�M�+{�j�R�rħ�K�ZR�>#�ĕ�oZ�5�Y}r�"���Z�:��������w\���#ح&��S*��-�"���+4zs��f����U�O��\��~�z#2���ص���?ݽ#}v~:�H�_�p�;������� c7�b���@�!�rhM�\�*�
���^t+��K%�U:�V���$#Nv��n&�I��1��Nj}]g�GNP˖��I��ܧ�R��;(��к_�Ǖ�F	��9ϛ��\��Y��Xh�75�$fWL��' �����֔ڜ��e�����$rP��>g{��F(bN�1k��������p]�j��>9xP0�H��Ǣ0 ��+]��	D����q� E�Z4QW�'��������dc���a��WCd!.d��a��V�7ry�f�|9*�4�I��&��V�\i�#0�j@?H���(�"ͱ�T����;�7� E�*S�l�x0p�=Z�����4�
U�f�A3¥�pXB�gI���n�:�����1�G�כ'�o�{���%Z�@s�(FDA�[�y���]*{_��c�Kd53��fR�.;���@�Kjz��Ϳ�˰�?��d2�ܤ��&ȏ1��\���AW _�Q��NW�9�����X�$Gyr����X�[GSc���_���`2�iq�0�!����0�D�)�F�U��@�G]SZ� (�O��ɫ(�OH��긅8�[�Ȗ�G������Q1�� � ��Z��w�4px���^��
�?�-j��e��f���v��q�	%��[
@� 1܃�_�au��3N^mڗ��b(c�P��3��Q1#�S��	��&�w�� .�n�����NZ�UT2b�%�k+Ӷj�V�����	?6Cd� �Ug�Ll�}Ť�n�5���
��rUn�_
�g��e���F9�M��A��n$� ���1�kc�h(�^H��y���.��>s��rW3R@����#'�z"�R-���ˎ�j?)G6�)�U�>�G�x�<rH�7~m�O}������e��g���L6v��n(�I����]�G� @���߆�>Z��ym����>�?��V�;q�$���e��W��a<��d�v��:N#�dyb����,r�z�V�]�EF��;�^ɵ�2yg�Tf�4�)Vn-�������(�A�\ƍA]h�{`xV b_-<�I�d���ʴ�]M��ĭמsߦ �{�
���\i���/���F0U�֤���=|�K���$��Pm���l��ȉ�K�S"UJjB'X�Z�퇝��׍��An!�!����0��Uˌ�����B��~�z�0��-��eв�8�ⱊ�T��EC��[=�K����N�bI���n9-�'6�- ���kS��P+�c.�͖�?�o3>go��^���:�j��'�kfMY�χ�egA>5���5���9ژ�:�s���M���K"	������͞��O)D�)�E��Q��<J����V�N:v�������N.��gB��K����R�U�$�t�y�R�|JO���I��p��*�;W�%����Oi�����}p�}JW�I�����ǣ�%&6pЃ��ꀕ6Y�8�Rr������G�2������o�tM���ڿ4�y��P�E���ʹ��xoF��H�����P�8s�ө�Јv��,��)� eQ��4B�}������`\
F��������>Ĝ�c��Kf��7�7�)ŏ��.�OeSBZ���}�.�:=v��ȃy���j�s�W���Լcϝ^��vl��D��I��e�Z����X�c}^�F �Q�؊r8��['$>|ϥ�,�E'غY���)'p�[Ꙇq�H��a�9�y*P.ֵ�/����ua{tH�F����(�y�_���d=+�=_5�!K	�} ެ%����0wyWW����2?4W'"������YX��u»Dutv�(�!J@HJ�4$�4��۟���nY�{ �R�C�ޓ�����$p����?xj�����=lH8�D 0��
��3�0�b��F�^߷HP�(}�.Zg���XHS�N�1B�˴��Gθ~�{23�����}�aS�r����"�EQ��i$���A�S��_��Lxm�~۩�L-,���ƍ� ��M?��`> �x�y�҈����=^�O�b�:��-c��;kY,2��_��c'�Ӻ�~c�~ ���&�!H�5|�GyM<����0v�c2���*l]���6�7���)�Rm_ ���2�.8��]h�p25�K ���mb��'����ѥZ��V������FS�Kp��#�|`��
WU�OAyD�w�E���!�o��7{G�f債~�S9��/U���o�������ʸ頞\�f���wK���lش0s�ma �|�B^�P��d�~&�(Џu��`�QP���[�Id/�Kw���m�q�בSv�jA�RI�&:�0�ty$B�=˽Y�L �Ec�+���U�g<B�+��!5�@���*+L��ow��4�zdejV
��ԏa�����o�Ϡ��s�J&��ֳǺw�x{ۑg���uk�G>��W���#s��P�D�L����$>��9�ݰ�&Q��XV�r�q�&�V	�Y�Ж�e���������u��Q^���h"�*�RzA��b��˯�ό'X'�yg7�q�}�����IE �!6r�=]��e2�M��{����I�m�2�m] )��4���xc��t�F���A�ޫ�ynW���A��:K�)�p&��`��xR)���9�=x�
�9A���١�"IOv����"y����<�ߌ�&M8���戆�[i�=�}v�[���9�:e��V�t�5췎C��pYqMcp�t����l��)yr�@�$����$��h�hWj����s�H5�x�߉����6����@7K �֫�#8Rd��C���ș��>���A��]�Q�J��*.8�>4e^:�愸�����b/;_�vej@*�0O4t�G�֭GU�߽\`��P0�nӤk�L�yD������'q=��`�����o�}Uh��m�/,Un3�@��<��eƠ����zʕ��О-�_Ke~Y�|�|��������#�Qvt~g읕�5e&PS�ՃyT�G�CdG?�t� �[cv�k��ZI�HYѲT���^���Ɨﶰ����QD~�i}r�=uS0�w�g�}w�z�=;u����~M���uh%�]�s~j06�,�8�qHvz9�F��l-ŏ�U�h:��+DihȬ�8�h9�MF�sRb>g pl?ܒb��!Dҁ��(g�&�D�5�CT�X����[��3��GP���BgIӘ��<p��\TQC��ڄ�35�NX�  ���������'�V�t�י�3wŒ܄3����$�6Ĥ�g]��﹣�y���J��}�����EK>�����''��r�c5��U���r|Z�HG���G���?�G�N!�>%�|�)3�e�%�~��b�4&�@i�вd��v�T��#�q2ɏ������{�wJ�z�<&�/�~Ph��/�Hc���MPJ�A�*_ �`�%��X�)8u?��	 ��pWV�G��'��H̝���h*���mйb@�%���ϙ��5�g�Qt4ٲT��;��[n�}�;��ŖG�Z���W���k(�_������ל��f�6 k��u!Q�:���f��6�����"��Ց�:����L���� ͟3+��2C\�1��5��!4�W6Z���`��B$�BI$&Ah����"��=�����nrf�����ye�Y�N8Y<�7�T��g�ssA��cJ��N" ��Pڵ��!�<�{�_IRZҴ=�A�,cOzHV���'�ۊ��C韣8&;|f����@���!R/>�h��lc�τ�F�=����_Y������Jz� �7�U��z@F�ιjx��!���E�w]�0�˛�v��V���G-���.��P4A{�ϧLT�c��
��� �`�p�@>8ݶӘ�oNS%T���7�ٺ���s����X2e�p`���� -�PAD�n�}�z��(�}N�(*��k�?�+A�岡��*�6kP4נOY���a�>e�q\����?NX3�X0L��G�-Z��yǯD��e����,��;j)��SA��6zW�!���u
Ƣ�Z�գ�S���{����L���L��!���r�� �ě���_\�oT�s1�u�����&h�@�/5D�j��s�P6�<#�ǢJF���$�Q�������4y���ה�t �Z˿SuBC���\�̈́����:�eys���Um��kq|���=��X�G�
�?}bv��(u��3�������Z�Z���.-�w�Pl1�c�A����Z
�%lmG����l���qZ�H��m�9�9���-�-�ځz�rp]�8��K}�O�����p,�P���6�BVK'c�
���,��bG%u�]��8�Ld�c{� b����?�mj�	[���·����O��QM�Rt헭��*��a��V킫\0j���b�?&>^�4�e�dc�g��T)9�1�D8�V���F����I�\��5�hyiX7S���u�'��?m��h�"<5�s@��$YJ+fg^�z�5�1S2�U�V�5�o����%ȵ�O)cQ�~����Y�3��rA��E�|�d<��}-0ϻ��V�.e�4���<H��,$Zt���~җ��@W��sWʨ�7�;&yD�⩇>��j���܈�L ��R���b=5�dT��\�.���B�)�i{=W�����Ɋ����>b_�'M0ٖV�s&c(�M�Ѓ����v�S0#�ݭ�{:r��':��]N�p	H���S|*nXG��I�6�V�&�� ��C�J#G�R	����<U}a)����kh����փ��"��%q���C ;��O�T|��M$���97�C���q�π�s:��S^_�K?��n ��,*8�m��g�8�<?��+��K�Ap��p��8;���FL�o����$e+Nk�Oքa��v 	E2�`�Y ��[��8K�y�U�ZN�b~!���^�L�vY�L�+{��F%�=H�Z�`~�0%�RyGV[������M�(m�I�[�c���	�X-���ve���F�y:y�u�{����n�����3��DV`"����u(8�N��S�WŰ�1���`J��^�Ь](���`��(�\��'�wM:���#���to���F�g��{�b�"��m��7��QR�}=���g&�blz�,�h��:���k�\[����uqT����.}�:���]�C��uS�H��9�G"��[~3,� Z���M��AKK�ԍw3��w��o M�iZ���t��4,VkJ�O�_�����jU�+Ej�������H�-p���|���&A��K�&l��m�n��C�p,;�f$(��K��l6�?����u~:@�����J2No�$�ڵ�N �p�����*��MK��)|��(���#*	����0rߘ���"m��e�)����ꂊ��q�s�8�?8��cA4�-�TD�F��z��;��#�8�_���d�@��)�ˏ>Pb|s�)���J&��t���4�� BK��g�����nҺo'�b�`���م]֟ �����܁��� ~K{�ƀp��a���͏��M���FH�f�� ��_�H
ek��OT^�&	�(Mb{՞5ox�/�؁�Sq��q���_=��sR?2�ꐧҥwt,�I�5K���L:�
�Ȱ��-�̭���w#$~�__=��Z� D����r��H�*�v�V>ٛ5�'�|~�)�o!�'����B�=��M�#��^�/�`���zfH=9�B��O�~nA�q@ �;o?,޲O*�e5D��\����Mp�T��Ϩkn��-�SWRT��4P��l���=*(��o�#��H���w{�#��R�BD+�)㜱�Q��G��o40 `���ˣ?Ć9}���i����)`���MY����T�0�Q�{��1�h(
zV /r&q�����&jeME���,KZJ��	�X��&�3�Q焝.N����q�Fўl���6�8#����R����GYl�%������5�m��#�g� ��iqkp�z��Т��x|�Z:����	x�9y`��9�V(�EZ~����Qy�������P�`�e��	��y:���s�'|�5��"c�����:���Q<�7׈M��vK^a6�'K']KK���<�RK��`�`((��(Y�l���b%����h�ҡav�Q�X�;�U]�+�+��D�]�\��o�V���*v\� ݼ����:�z.]�D�F���ԣ�GVi�'6��m�~Nk�X�Sɸ�0`�
f��t)AX�<l������j�kA'��4�����L��o�œ����=�@w������q� �m�1-$8f&p{ٙ32���9��^�,P�fA��{0��Ѳd	�+Y��[�{n��r��C��t�A[v8F��6 ٕZ
k�������ƿ̃��9!�����[J� �Õ�ՙ�n�+8ɭ��%��Ht���O���U3���2�|���x��ߥ��F�uh�0��G'�L�8ݢ}�Z��
������ȩ�L�6ܫ����)��P%.��+<J��^��\u��f�W��5_��?^�� ��8�ʅh����T�<�71��6���Juc����G�_1��u���������i�&�	Kqѷ�	A��o����4�.3�#�.Pj\8Z�)e��������8ڠ��9z>�G$H�_TE��E�3��׶����Iǿ���D��T#�p]0Ԏ2n��.�~׳; �J��h�f��dp#�I���O�&s��m!�At��H�ep��i�����<aI�2tJ����ߓ� Sg043�6��7���y{��<U�o�wT��Fv�j��G�]A ����(�%��=A{T��{vP3�׼�]х��}��3�BD^���ݰ���w~��.��:�R]��ԫr�mݤח0���n����-)�� O��⣌��� �S1��-������c$QN���s��A~�+��}���sAP`��){D��I8����2�n��}���C�/�j�B�o[3_�~u��F�߿H�b�R�y�J�-��ww��8'�k��۫XD⒂txu��JPsU�(Z�gGV����J�6 �����W$�	8���)���[���5������{��zތٵ��*��(L��8W/
=���:���V��j�][�R�j!\L�a�<ҷTb]TF�͂�UeQ�ѱ7
қL�hu��y�����w�A��@�،�:����No]������w����T<3>��=�#�l��x[�/e�EBǖ�~���>��ڽ���p����b/�YR��+ے-�N��AJ�C�/y�A�wAo*�;�x%Z������o~ӌ�G�_ ��{*T�m�E=�@YՔ)5�U0n���.N�0}�.���-Ęs�A�h�ƻ��8�)LB��>A��G%���&�V���/��8����� ޗ7�@�T� zެ3�,��h��瓺�O�.�GpdSW���G�q��o��'�;�4���_��i�]�~;����ܚ��A/w [����/�l(o�HG�T���Ey�k���5|�ƬK�`�V�=��P��4��~��}y���1�$�.z��n�`�5
����rb\`��B0�0�|��0��	4��"=��&���_�5cA0Ӣ����Y����s��e
�)�`[�h 
Q�!����[EI�'M<0kz�:��'f��F�5�I*Ţ�%l)6ŘS��ˊ���4�C���g��)�7s2�/��xW�v�A�|J���Q*�4(�l^�"��u�^���{����#����(�!yjm�%�g��?A�b���7* @�p"r`����A7�4'Q@�t�6)g8����O�s^E��0�������1G��xF��j�>�Y�$7+�X���U��u#�n�_ϴ��av
sQK����o�?O�y_4��u���K�5B��d�Υ����� Ԧ+jT��ɓ{-��m\N����Q��v�)����i Z������aK��Wؑ~M4�������i&%c���c�I,�U��� ܓŘ)D��YL`QZ�s��7��\�}A�����z��[�>�����C�p�]�-'�nN/l�Qk�"��q�����lw	�˪��D�S��w΋����RRʑ��y蒔 ��-G�B�To�\C���	���M�Y���v9�"(<���ǷuS���A� VH�z��W~U���B�s��i�ӏ��
R	�]�w�pA������=�5��Ͼynv,dn�T�دv�ɔ����e8s�7�nj3a������ײl����V�d�+:k��ES*V$f�O�{a�X��-�1���Ց�QN_� /;��E��N����L�����ţwR@BV6���y����M+@� Z�eG%�t�!�=?�>^;�vu�`K*��2/t�������<�ƌ�X�����e����ѵ�ַM�u���A��f�
�q��� �G�*���P�J��� ��ո93/R���v��_���f	4�OR���*?.o���aW��.\Y�¼�:N��>�Lf	I<����d�+8TPmv�[�	��jg�ռ�>j\LZ<���t��G��95FHt���*T��j.^�*?`�_��S�షEx~��!.�sx�Bܫq�.�������n�.�+�z݂�����Y���N�#B��~R��`�Ŀ����W�e�G��y*"�+�`co!���HOw�G��H>y����9�w`x-�a�!Eo�rd<�}bh�~&��$�a9��p���ק+i��{��M5��*�$�~t�m~5��QKjpᛲ��l��o�fk�~-��Y�ё��O�㏣?��W��񒥏O�aj�^]bw@O�4�r�����z�ge�4��ۍ�3o����:�����*�@jBj���-$ߏ�2��?u�v3��l���@�
%����֫!�>��s��
ʘ�N�}�ک�2��ٳ���;p���߉��<�ne%�\7��[���'t�Lh��I��~,8	V��l�͌J�K[�+�l���'�q����Hp���hVM7�ܱD��c��8�@�S��p�:�`8���r��s�Qh<H1Y��
|���"[��+����n� (���^�˜��z�^�v@Eާb���P��S��.�J�1a�r������'��I�Sk���Py���}/1s9���F����V��\��s�E�.�#9�6�?��f8����]��/��uME��Y��Iz��� �$C�
�ˆ�'������LcI_'�M9�
2�3�݄e7=M��ͥ|%�%����7��Fe^��n���=E��=2�E%NM���u �A�~k��0|'�g����1l.$
S�
��G��Y�R�Y�(��@'tP^E�  �c�,B5N�~��!܍,`��,&�U��O<R)��φ7����$��/$��UE}Viތ���V�q'AVh �}��C�d�~�Μ٢�O��S�yA��a8i	�k�[;b"N��	��	ivAϊ�W�z���b\8����R���	���+�Y���1�И��L�
�gkkܦ��,Ņ  a�m���E�]�����X9s!pe�h��@�0�]2�68c�ɪ���}.�"����x�Rj@��S |D����rڨ�o<�H�'�� ��-�\�Eb���b�����-�N�<�َ���mΧ0[
��Ia���+ML�t��+<���]`���	mŹ6u���
D.�\�R.ߦ��T���;��P5L�v��1����r K�*��+�M!)�w������?�� ��w��Hº����`��;�:Eb�"L���G�H^t_�'�'"+H0+����a�kR;��18Y��;�
J�W�h}�\$i_�3�a}� �:�������[6
�ܘ���
m��6�r��]��!uu�RE���]��͛��(虆B�4�s7�YeH�b��\�hb֝��{�]SG��`���F]fv'>j
��Tc_Z%y���V*�%v�7e�����ֽ��2���3�X���B��m�Hր��cE�d�űU�	w(� E.��kVS�N�=BsF��{���%s��`j[G�ᛝ��K�xp=�H��@V�!t�s��0�Wk�3�������V�.�4S1�"��2B���� �O7��Y7"*[KH;
��My���w8}k�U���ǰ97VR�Z�!3�����C&�(w��+�YR6�	���%�?u�u]��3���rteW�u�2=�ڔ0�X-\�D(��u��YL�U���?O�Ѡn]s�1P���">qcs�6������a�$~y��3��ٸ%˓<����1|����	�2m�q䢙F�-%�AG�S?���l��ξ�R�+�9d6�A{Ӛ�\�P�� ��wgl��|ݚ\�CE�Ȋ̢{b��v��u"����p4���x�g-�Qn������0u�3:�}@ًF�7V�^��mC�z?�@>��r�h��S�M�	{ ���� `��C�e�.�A����wA�`U�Qu�O�J�w�ŏ�:V�a��i���Yn��;�x�ֶ�T��I��(��B�=�,��4W�<�^�ߦ��$�~�pa�K�ٛ���ב��Y1Ɔ'���Mv�e�t������K,&�P��,)Kcđ�ڼ�g\��ϟ���,Y�"���C�"���v_�e���g�7�_	��쉝�\� ���C�%�ߧ�f�շ��3�dJ����bM%�|�ڨ�+���.��Si��p[9OR�����3�~'E��V�l��[%}K[
�!˅��۷a��B�0��KpZ��a��f*͗����K����� ��Ռĕ���є��l 5� w� \�ޔ���X&"RԾ��9 ��W�'q��a`��/�١0g�⊂	[���oUH�9/����I�xB-J��X��l� �\��T���J�r���GƋ�!<�s�[ v�/h'z�dk�ҫFD���2����'z��p��k��M$��fd�=Z�m�Ur���t�҇+��Ҕd�]������7m���U��|����C��i_q�r�n��kA��	�"-��Q㦔�6�nCz��t�����0�k���J�N9j�i�ѧ��nٍ7\DA�ׂ��4�D�L`��p�	#����l�I1���c�/R�g3��,��$<�زa��¾l��v+�SK�� �d���&=�	�U#��nۮUQ��T��*���hR��������No�`����)p3ܔ6L��ψ�+�g0MXDegRydD[b�?�3��_��X�Pp���8����]���<ʲ�����i�.�j���񕔘;p�UrK�Z���k���F�<c[�?�K֕�9�Rڳ�䝲��_�V����ͪ蘆BM�JxFJ�&Bwb-̐�8)]Q^\[��w�DXV�*��Z�^���`�3���ࡐ??Sn^J�	�<�4��8q��c��j�?�gB��j�YN���d�Mr7s�sIex�Hc��򫫻qi���֝Vx����m?���?�ܖY�P� o��f�)l;_ĺ�&���ٚ�E�T��F�u/Dh}�n�e6�,}B��#�t�P�Q"���|���S��G_�.�c� �awC���m��ӽ��1�9�Q?����Q�!Cm��-,"d7i+�j�o�{Of�[����H������a���ί�F�(�x:��Ԇ*-n�'��̻7��@��K�d�23�5�t��鸗����/4q��	�>���9�</�2`4yGPu�o�Hw�������4A�1�pk�Q��B-vnw�3 �g=oF��kJO�Ə?���)&��/`�NHx�3�Ijc$��$�j]K���m�<ʴ���e����}LZ�?0��+n�t��^�Dΰ=?����a�ك������t�%E����vB�O��9"lR(aXp�������&x���\���γT&��s�DV���?R��$�ڬ^}��A�K�(�1NJU+i��!E�A���Va�˽�;��d���띟eߝV4ֿK:i���Z�2�b�D3B����(I�K���$,�_�B��):5��?�'4�/��k�)1o�����?.2�o%a��T�6��M��^�ō�����&��A�X����gw�CrFuo�.U�"���D&�C��v*�sd��=С ewT`�Qj1O\!�����[͒���d���[f�����~[�e����5t����Y����B܃bƒG� C3�zЄgT����t�Pc��h�)&e�p�"##�{ߟ�Ap(�U�S/��A: �EF�beg�S���Qk{M��ńw�⩘����4η�JB�8x���#bCo)��歄����g� W͒��������R�O,|0��N�0zu�RJ�ēɃ�*��j CQY��)ܦR�r����>-�	q�?��yA�C��(6��7��ƗiiBO��VJ�I<����2�(X��
ad*5�����ffҦ��穄�2�����A@����r�7c5k8Cu]u(�*E�f��6}WH���Ժe����蜧 �ܹ����v��)-�/��T��&����=��E���x[��+[�GWft�ot
���k��6l�������u����ij���0ʴ����IJk���=fM�釅" �O6�����*��A�/<a>`�'�ؠx0�'��6�3(��u�1_�^�S�T�A�ڷ�9xl�B("U�o�����>��,i����i�'�X�y���X��B�9���u4�d��S_��M����L���
�S�K f���;d{���&ˏa��A��?#�T��p�/-� kxe1fw�̴�#迉S�<�x��D+?1 %Fgo@_)h3&�C��m���;Z�[��~ۋ���w��G���-Fܒ�3M��?�eڥ�mWfݕzMq<�,���������+�z�N�QL��{sW�#-�
�n��I�51�'��'Z���Ķɿ���� �q5���fF����h�x�zd�2j�!�.P�nz��z�< �pF·����aOІ?�#P�����4t���)S���� �m�p���,L��#I�R��'>1#>r�~�VD�����a��U��Q� �}�"��p�O��ј�7r1M�Fk�eM���X@���K�O����P�g�ی7ȂB"��l�iD���AS䒌�y.��p���so�!�yh�`�-�v���4A�/���ʽpF��>��)��N��%�i�#�"��b�c;�gY�S�w��=iH�bi|a�6�lFG��Єu���xT�1��KM���[ci�4}R�6�hW�o�G�G�	�KY���12`��'z�.(DB8���D��Z�t��+B�6Ur�۽�b��j�]鬊;\U���-$+w>��QMn��9�
H��|1�	ȼ���=���0��'��C���s�lp�C��o^��;J��mOBo��&p{t��Z-Y
}�ގ��/��q��9$�*\���aW�t�D�\ݷZi�bg� ��y�����%����)��v����0�t͛cP1����1'�W2˶�ӆw�C���|��<��*9<W���[��Wum��[���8�x��Į]�;9�Y�*k���U=l��?�f��!�w�t<OO��$��m����N>�_]c����-��x�C\�m�eĹ2 {=��W�Z��q�u8��|&��Q&B��`eM�)�G=���{�@�}����k��5����J{5���UU�DW4� D�% ��=���(�5�0nu�N�����Bt���}J?Q{H��K�ƶ*}�}	�ҁ�;�I9��S:��f���J"�\�;�S7
�EY��D�6d���\�z��
f)3�p�M�cu��h���J�(R+���!צ ����L�x�^.Êq�p�n!TuF ޕ���kC�z�ZG��a�e��)�&=�Z�%�y	���6+�}^���m��vߞ�?��?c,*�3�9��6�c&t������Jz�M��}~foo�����
ͤ�:��u��P�)v����>զD&�Y�Y٦8L�55�J���og(��鮢	�=��+��G�iQG���y���$5C*��5�i]�/���X��Q��tח�D��V;o5#�{؃Κ#�*��E-�qޯ~�Z��N�k[�8���}�ь�9ɲ#,�V���c�x�:#��7��c6��#`��k���˂.,Q݂�lr���μ�]Gh
�D��v+�*p���"T-�S��8��@�1] �-���垊���T1��t���'IN��a��^� S׉ɗ#��C��=��(- ���5%�/Aز�I9j�y$�-�~�Y��H2t�Z�>Pf�2�B�փP��nx܄6j	��<d3Q^���L;��'�����Z�\�4��y�rB����[j�4��1vUT�h��ē�j��ņ��]�{-E�I�;^Pz��Z��H�Wӝ�VpFey�Z��Mp��h�4�L�W��Uo}#��-Ư�WX�P���7h�9^xlmXv��S��;��=E�����}vU8(�d�i�~i����~)u�w:$)�}_�o��Gu�<^҂,���5bTY��q��=�b���%�N�����XF�iqƁe�d�S/��x��ήL���uY�� ��|���[%I��d� x G�?�j�v��o��A]ъ�K��0�z]�H�?@����� +l��V-C���-��0a���O"m_\���W�
�R��v/�.lr� )�㟴'k+�j����Ӌ��U�2�	�` �^��Ή�Ul�
-s�TD6Y��0r%�Q�#/��. �T5�y�yo��(0�TvS~`N���W	!���8���f5/�Ak��,g�͢��%v�-��`2N��C�VZ]�B * 3_����m��k�Xأ������:��*w:7�<���]�@�{3xhȼM��d���7±A�,��y���3x-Թ?��2��s�e�Ӗ�W���>�RC�Tbpb����(��E���K+���N�ОU	�5x�c���M,V��5`��W�\�x�,����m|�;�O?p�7��}Ne'�;%���(�M�E�;�f�ϯCs�56j�r5�E�5�,տ�������2�gRb�w�0�I��ƥ@_l��ug���1S��<��Qq�xLv�0���Ԋyˍ�5��~ɜ�[ ;'Hye3��{C�H؞���3xw�Z�22�C��/�H�6��ǭ�k"���Q���h�vx_��60!��3��="5HX~3�o[�0��<M'�� Y �y��sO{ݶI��#H�Hxߏ��)��V�&Q��1׬���8*��A���&x���uD���Gξ-�7�mA����;1��:D�B��Y���npkJ.P�8`&���!�/0����_��ú�,A���`�xm0��T�M����.�ď6>�p�G��`
!���X�v~���C���B�?��j��P�IC�5E�ذ��6��zw?n'����$`6_n7Α�pP�a�M��J��L�̖�r���D_5���f����*�`˂�R]_��73�l�c�
��^6T>��&�68
2� �jЍ�+W]�>�y�x�(G��tAO]�I�����rs��s�������#xH�\�a=u9�b�2�ΐ��CB�JL[�H�\�����sx�Ϻ�P�C�X?�4ݪ��FU�|�c=�5�##eq�>�Y�J�l<�����(?��2���'3����V��W���O�e�7�5�}JR���^/����}b�c9�V
V]s��=W��=R�;sٮ	��똬_�G�T���uw�v6%h�ix�>�ǉK���H�����.֧w�'�����{��U}Bl�V$ʑ�ё��⁰vi��]�كnZ�hYj����[Lȁ!�I2q��_�e�\H����[�<"�ߢ��!�Z��rE_����<�C��T)!�0^�ⳟ�ˋ#�1��ײ���ɿBQ�jM8@�H�݂��LÊ�N鵩"k8�0#��˧=2���E�� �����b�d���H�N����)7��
������	I����Exh3��k���`Ԝ[�H�*Њ�K���)��!딙g1 �X�㸃*�Tb�LQ�ޫ��F[�U�1񸶓��fX�it���}�+�&�`�9
Z;�m�͑GPIܸrB���7S�
}S�'�S��S����ƍ+1��ǉU�O��2��q�s�_�Ɇ�\��t�ꗶ�L	#Q��&+1���%|`����˗����^�~�,2UrH,�����Эy���sŰ� ��KO�КDGY@O�\���0ym�$�u��܆=�TC��5��k�Q��t����S���k���SiI
�J -5��9�n�	�q"�	�O��­�w2X3�6���Y}�E�Ӂ��ܟ���-Gj'q�I�X���  ���^J0�|C��bK�=��m�`�	3������e�(��rp��W*/�4��2�!��<S����t��n\tv�~M�����ef�۬.Xy@���*��6v[��o�u�:%c�ů��c��X0�A�ݴ"��#=��	���n[�)��06�m��4�/�V�V��[�Jg�4y��*�z���@j�Z�[�D����nS�»^D��e�_o���;!)`�0�x$?yuif�"V���n�agr����0�� �H�������`o�|X�l�;��2AUW\���oC`��ۨ:qMFJ�
�`�7-��*�;`��m�&x0��R\�fh~�O�X}����iÂ=�V�l˙>��`N�*{��פ�<� � �
i׵Իa)_����N�3B�g8@f-��.x�3!��?��׼�[#��&��� J?��Y/�@����s)�.p;vLR<���hhoB�Y��Y��H�"��a��=�q��Q�'�V�]�7둑�]��@8J���TL��3NS�E�%��Ҝ�b�`�	�.3PZH�P�#Im�Rl�c ����Qe��&5tƃ�����.��P�`��91�j�*1[���	��H�\��+����^�Cp�
�Y��9�ȏ��@�9!�j߅���
��]l��r���@O	��2>货-&P�4`����ԙ����Ǣ[j����`Y�R:U6!5������\��D�.�&$u��!jt�Dr�ȳ��ߏn���VW�V�U(����,jO�G2B�|SsG���/��̉Ƃw�k��<n	c���7K�`�oP���T���xh|���EA���ۡi!S�TrE��QPL�N�ũ�`ז���ꀀ���=W8o���2 L�)Bn�������BIK�`����
7�ԅ���P7y�3y���==k?h��Q�vO����+��g��Ȋg�d�V�J��0-���mB�T��qgK?��F:�U�Ma��16'�:����&:)��>y,��5S�P��Ki`n ���:��)�� �ߠ�Yd�����A#a��g,�=���\1�W3�ڗ�'�nK�d~�#�33����C�y*n0�³-��R�r�|�(�s�f�\
n&�]#Z�%�a�G���t�y��A�$�w��m�����{��Ê�`�m��5��FP���U�z)�����*��+?�lЗG�q��x4z��W��ݻY���bӖb�5����Ӥt3�K�d���v�Z�k�l�t^0R����􃭲��$�k�c\�`Ȝ!QP�/�J�i"�)�̕���pN�7r�$�� �6�Y��Zx���!s���"Es����{����?]:ʇu��SQp��c�n'�8`(� �ο��E�ڧ��V��t.$�J�X���1�o��.��c�	am�c��DͰ�hw��%��p6�*��F���<�j���qM�q���$$�[�~�H���Pqf�U1�+�0��	��F�H2�`�	�!H;,ٕ��G��'�|x~N#0�g��Xf+6=]�Ik8�.M�#TG�P���wNPidsBL�6C�-��~@Qj5���>SIKg5X�%=j��R�Qg�!d\�"�p��=5��^�]5K�G�����~�N�;R]޸�4����m�~��M��98C�
�U���(�C���:p,V����VD�8��j��1�"���ƻ�uG
2���9��{����f�@���D{��Ⱥ��^2zf!��7�+��3f�Nndb&��8���T����^�(���"��`;��Oۧ������q$�q�ռr��x���e�jⴣ����\	=�ųEm�͛vU��b.����fM�e��v'#X�@�)����U��h�F'�0����pƲ��+� �_�%�T�w� -��'�Y$�"@0w=*��<A.L���V~�:�r�%�\�*�r_kF1���R-����;(���+$�	�z2����RD���˷�9��҇Uq8D�:}iٸ����������gς�a�m�	�`ß�C~��A�eOleV籄z�`S�oDO���>V�U@�|�9��p��TV[��OxT�'������J�Q���  \EL�s!_��,A�^w������b�ޟ�1�j	�_\�p�+u�W�?��]y/P�"۵\���1OQ$/�\RdݲK�fYd`�p�g��CW8H�;}�l�C҂�Fʕ�hq��yX��P����v;o�wX��hkT�s���rD�2�тF~��ڿr�*���f��|��li��x��1Ҍ	f>"�|��vb����n�ԒU��k8<oloO!�ha���Wl�;����4��*R�Έ�d��涱1�#�T�w	��O�����V����I^홛��]�@�ka��mX�
�N����5��3{��ٽ�6!��i�۶�ZP��ۈCP���Mx�� T'� D�����>�T͙0�S���=���^��]���i�{��B�ɑ��(�����U����4��\o0���T�F`�5��d���n��}��0� d7�N�ǣ�����s�����4��@άDL�4'f%*[���T@����˖��	a�-�Z�
5/��Ǫ��0j�,���͟�C�7�E	
w��c�S���}��-���R�*�ʒb?F��Ӛ�J�﹖]�K�`���p���L޹G�)�É	êshg�ġ �	���{�ubL3K��I�B��da[Zw�7~�~�	���� s�H�c ��As�����c�z �d\Po�ߠU'�q�v���ݖ׬������s!7�D���a}�"��|��Ί��i�d�xޠ�`��&V�u����B��.P�+u������F��[�[��W�ი�V�5h�qs�;�{��n��ɰ���u����_�!!c�u����˲�F):�%���O�Q5I ���G��N��Q��ތ��@�@���[��s�^L���3	�����˒�ÔO�Bﭿ�����l1�%��������O�u+74�꫚{�x�p���?��\T �h�{�
�pw���  G������]�<<ީ�a�+e�nn�S^ ���[�׈U��">:�5�Ϗ9l������V;�к��' yc��@�Q^u��_���ك�ۯ%��C��F��̀e�#�ݝ��B�T$[%�o&���'1OP�^ s��U%Cш�]_�Q��y�t�
�=�y*��x�Àj�`�9���� ���:tr7�7/a�r�����R[�x~p��r�8��6���@�E����T!�-L��v� ���i^R�vʈ�. ���EZ��c5�j&��;�B4����y����l%X)F�;%(x&��
F��=�Ӭֹ�ܝ�Z��#C(�κxG��7a����{c��"�M1)�V��NOuyP��Q�n���j��r��o�,�1>���ୋ����4�zu�9v�HȐx�T��BF��;�l�]Z����������� o��`buv]��#
ބ�pE����_����(�z�˺��{��������Lˢ�\i�ћ��<�&�#�k3r�LX�>��:!V;�K�K\�a�$Ճ`��Ԉh#,��5R�G6�S!G+{�k��	��/R�Y.�,zƛQw���s�C�������e,��5V�XsF�
9����W�W,�i�t�����򨮧�g��Uo6��v1ee��f���<��@����yVV�uy���Z�)(v�B��u�1c�AH	u׋J��ŵ��� ,왕���}$��I'�q����'Б�TO&� �<�z�a/P���w����dfZ7$��|����Ƨ�|*��� ��\�%È�N�y�Y.���:��s�U��j���;�^#���#�CM�.�n����V��:aY<oCڠ[}��4�$\x��U����<�1;�2�⤑��D$��E]�ڴ�Z]a����Ü[���jOO��O�������K���?�#�T�&��yr��Wy��2H߹�?�CA��s˖�v;=Z7��r)s����%��n��;7v5���L|�.ZN�k��1�q��Nl���ͷy�Y���.��P[{�ʝ�l�h#��z�y�>:��{L@�N�l~W�u;���F~��9��k PaҸb	?����������,��I�}]�>�%����j<�tQ���CmF�׊���Pf����t�8�o�m���x�+h���$^K��PI�q�|&�U�:������ƟDf;��/���in��C���w��`s���%~���A8�L!���5vG�
�u�鎩� KLm�j`A��y���Ɍ6@��YAIҤI�d�W�OQ�gx�u���~����GX��I�!�x�����p4۳���X�X.�`��i�e��~��D!���ܖ+���J�P��@Z�����1lL]� -s�xyT0S�\T�Y��0�i^��|!s��N���u�ݮo�~e�Ά	e�&7,	��:��`��.mC���Ky�N(U"����ǣRD�!qc"h�� �w7�0-dj��l����>�&6��5�e�TW��-'���̖J���G^8��2n� ��EyIg8�^R���=.t��ĖGV�Y4��Z����|T�)���
{��;
���k�l�>�|�������(K�����k�d��J�v;3{���Ȁ(y��(.l�d�O~%)�r�E1�����|��f��8	��`�[�nP��Z�j�"D��0Ӯh?�`�Dz��A���h'�yű�g�ſ3���u�?o�y[�O�B����M����aWu�����1IY��Ft8/p��`Fێ���a��B����x�6��kIzٷ����������'��qj	�D�Ųs{h���!����e�2u)w"��ʈ���	��r�J;�!��^т�Q-�c�0�>�d����C��b�0i׈>tۤxꚕ�nBd��U0"�ն�yXr]#�Y��� Z�0V�w��r	H࡛�\>5[l��)P�ha�;�n[��Z/xb�<⬵o��9��x-��]�Nh���eP(�FM��qK恳��j\��N7���A��8\Hic����z79����W�<z���+&��,��S���4�m�4�F��Z6��W���f^UU��:��d������䫮�p��Z51]jC�B���x�s��4��g	�
������������8��k�!�:
�@�F��#5$'�L֯W^�~Y���-�s2�(�Lo���#��/�(�IP��zb�z�����\Ж\hAc�BPhES��:t�Ԉ�{Ys���Y��,�ӿv�z�Pޖ��u(�_�!�����Uh��ΰL# �X)ڬ�	>��Q��}'��&��W�)w��B�ܱ���{���eG�ծ^���Pc�Е�r6�NH*'�/�ᢵ�B[���z��m��xH9+-᪔�ܚ����<�6�g��PS1s�,���@|>W.°�������|C���K@p[�hk�1) �-X�>,�#`�C,�����өUR�/eLl��8hh�kpP�<aq$�|"������؎���*x}DIi@��y���>-�~;Mǃ>�Kj�g�&�!A��R�ͮ�n����!��K#��ԋ�>+�$�i�mhY��{�M2�@ϰF��UD��F4k�ZF�B@ ��<ri�������I�~�u�(�6�/=ȎS=\R��2��[�{�����	��0�k���C�ᙺ���4������祢�Tf�V�)���Ũ�F����+���\�R ��L�\h��H����.C�U��yT׷��/��t�<�e4���[����"��Ϭ��ɇB�j4�'�=��x�-�X�ܛ.�ˈ7��4���m��ܮ5�l_a8(m��o�פ �A��8?	]�]F�d_��xz��+;��#H��DU?YO�G� ���)a�I�C��s쑃B��g�Ʌ)F�����6�����5qy��:N�r�,,RҎb����I�R�^�y���%�\�����%���h����ϙ����r�X�d�w��4�Ov(\�\��YM����f�'�������}�^=.�h�!dϸ�|o��]���9�M������.6����%٠4�HȻ�1C9���!Č��Ф��%lOݕ�B���7�$<�ޘ.�n
Kgp5���V��!��66E��xqv�7��H�
�@�{�QהV�=�ܩ�#r�L���x�����}���yvr�2*<��R5�Vk\��WpC,�����=�̔��1֏��(-��[���۾��T���H���jhպ��[�k�+�O_��N����.�L6L�9#���&>ᠽ�Pa�!A�Eo���_�����3����A�2�ǧ)s.� m�&�t����i$~�.-h9���s���w��b�1|gP>l���;<�B�'�ݯ ���QN}M��e�8;\+��9J����C���9��$1�Z&,eA�U~�iX���9R��1��q&@���Y{6��C�i�x#� e���x'2wk0�]��Tg��p����գ�XvC�y�9��\h6��[���)��7��F��z5�� �w�|yT5�.O~4�=��0��b-�d�C��Q��������l��:8�{QGx/2�����>'��5�iW��A_�y��hѽ%��E3׾��L�7�_�丰\�)�$nY��{��?��u���3GQ6q���be�x�H�3�f�n�^l�$J�*��7�!��*whQXy6,�dxm��b�]�ʰ�3\7*j�Y��j������F#aV�t�EY
�4�@�B�_��/����Ta<��;^-$������&<<u���q.r}w�9�������8����S?�{D�(����0������5@V��V�ۼ�n�ɳ�(�2D[�8R{n�8g�nځ��	�R�6��o��ŕ}��V���aeB�Qymr��3�&�&�+t�Tdl�(�^�ĈvE�*VM*y9�r?|�?�:�^em2�t���M��q_���Z�e���4a����m������e�Sù�c���8�Q�f;�#�������/���Û��eK�aNw�ׅm�q��Ix�y�$1oLB:���2���������_�c_
NZ��¨�(�
I�<�4�f<�*w8��{h�ϊQ��3�9 x�	�P����CA��b��n���CD�10I���~0l�����5��i���A �_��Dńn-��;�R+V���hG��1	e6���b@q�񾆜"���9����1��co�#��$��#��ç� ey�ny��Iq\���K1plԀFN����Fp�����hyg݋U���m��c��_�=~a;ۯ�/��8�*y��AB�/)H�o��F����u~���,K���U6��P�nXvZJ,J^];"�Xꬸ.����&�����nt�C�y�MBa�s��� �`��S�i���j<'�ʶC�C ��&���s��`�/�C�sο�x����k;�'C%pيf�nm�q;�J��!�h��w)^ s?���2��V��(��{k�X\|o2�͌��v+���
���G���&G����O�3cS+�nrk��8HL �q�O�G�"� ��Q-|���L��k"�����s��SE�/�ĸ�Lܖ���,�a'��"D.�f��O^$�6#�����#���hDk���7��J?���J�?}Eá��c��P�D}��R����_�W�1`	~�N-D�4Gو���ݚD��z�_��W�+<;����d�^�����7�r:��S��#Ԥ��s0e�ɀ��8ExdF��NcRdX�
U���?�#�O�*=�!i��x�o��8�����ƔU����p�V�=V*wU��,��Ql&� CMo3�� ��O�q�q¾���^�.�}�FS�Mg���*9�B�(�ɱ�%�W4Q�xU�N��_f��iOu	چ����&�@�Tr�;��+޺� |E5yh�B�lW\�G��¯�~�gDEy��[@�&�vD��͎'��Pz8�x���а���#A����U ����CÈ��ů��!�QM$Ӎ�TR�����r��5|5�HR]�g���w��������`^U�)�^��3qg7��H�DBE�3�P7��Ԑ ���C��������û�xh�~�˰�͆�\������ʯL�+FRٜ�:N���W�k�xٝRp ��UmY�"���5�-*~�U�����G������&���g>��c{Cғ}�~��H�c�wI�*(��@gOUN*=�2���L�^��. x��P�tj�K��c~m"��f�˸����O�_h��Μ���)ד���b�=8�<;�]�,�:�>t�$#�A��B���q���_�à]e�_�c�lV���?.�զ�L������y�雉�qt.���*7������i=Ȇs��_[ <7/�4���)J�cs�Ǚh�6y]t&c�+]��4e��[d �2k�Ӝ�]*#�
��_h�zʖ���tN����W��Q�(���w4����P�B����{�D�����dSfM��l���/q����jU~8� %L�Ţ���D���\�yHa+�p��r��|X�7�U�׀=8a��I����0�2ď?4j���R��%�x#_j./yD������ݔ� 0b{�c����Vd����5���Ki��9�DC�y��0�U�/��������w�U���cE�`�/��C���:~6����M�Xk�(���n��^6�gM8�D5k42����,i![�8[?#�4W���}���$kj�E�a��Y�S&	���ť�x9[@d�(ԘY�4�n��c>v����ݴ�8��_UF-H�W��i����}���N�S�W"pҙ�;1m6r3Ti�����]�c�ǌh4s�����7�K��i�|���n�H�H8���W�ajq�^�f�����!����%Z��:�����Ҵ����S�㡡2��2_b٧^Ox�d6��2>���L'��Lک��x:jR"��v��7]4�Nz?�W?@��W�d��/+���q�I��A����ihz�l'1��4�Kyz�Z<σa��O��"^�])RŴ�="��~t����4"�.Dplf�2&S�!M�op֠;&�ה"�::�K�fr���+ܠ��zd#%��w,�B��A)�;(D�YP��vJ�0�h�����O�߬}P�p����7���u=ʠC�H��[q��h�Чw_��yGR}�a���-q����l����A~p�ٕ���ۣZ
�7g�~�Y���?�_Q~	�W��5��O�V�?S@u��q��n�Q��$��F�͜�V��\{lV����pc�l�?�9`06��ӍGr�<ΩO�v�ԟ�㣯�y���>ڟms�B.�;�s�}j��]�J�Z�Y魽� ;�lc�z���Rۍw���ޯ�1ϯ�Y]ݧ���T������g؝`��f� �I2:q�cm�0f�!���D��P�'��vf"��p)�"$�pఒ�E�*ځՕG�WS/�̱D%ɍovd#t&���E�ܼ�ξ�f�U@_�*�`�<�R�̪�W���t"E�`���&^3��+�S�b�r��&:��ta>c@��ȭ�:k�b1,5_l~c��?co�&�du�&��d�A��(�������6f&SwU�h�ToS�h(q��Z��@��E4�@N_m���e�_�"�>-�w6����V��=s±ܼ�{fp2��K'��"&�I"wZO��˯���2t�6Cɐ��i�v�u0��j��r/nɤ��J��v]>��i(�ګ=�¤�k�"�.IJ��q�87��vHkQ"3�2���lM�}<8��JV�E�O	&"�Lވ�?�\����w����Q�GPn�TR��b�Bls�{���s������Y(]���o�����tR��nT72�_���W,���?�t�G���}鵟���2Ŭ�rX7��Ɵ+x#č��3-�+��,���D �O(�!�:J��*�}u����zmZ@,�zČ��QVP��j��#�?�q�����9>�7����H����@�=�T����zb�,��i�7�:�Ɨ�o<ݢ���(����
���Y�Z�#�Q6�)賀��pes���Z�'�UYFH,Ao��?����=���ێt$X'�0�R�b0�k����'N%�7��!�Rq^ޱy��w(�H����T9D�0�qF�l���C[s�!C�T�n#�Z;�P(�쎪�fĔ[I��ѐ��H����K0�p�eb�In���#��8I!C�:��"d�q��K�K8�#L�*�@r�`Sy����<g9�\�����rm�E�\��.u6i��,�+gu��D[��a6[X2QV��=�*�J�C$eB#���|�N�2�K��I��o桔lk���{�rE��=F6&-D��5��Zkn���q�����H[g��4��GG�2���pKFä�xeEgY��q��I�[���H,����T�'�1�%W���pJ9���Z�G�W��)��j�Gb�~ +�d�o����;'����c�'��1��_:W�Xנ!l�Ԣ 	�~
8TH��W�Ǆ%m�#���G7�C���8e�lv��P�W�nh�L��9��Z�P���m�$!��Xy�ЛiM��_�Qt�cyG�^�[0b�� ��툶~��q!����P�U�ď�������Hέ����x���#�Z}�u�r�r-�[cDW?w3>�׃2�� /���.��\�ԑ�fץAu3�z�����݊�c��D"��������[��P.(Z���14͹���$�n�t=�ᇃ�ͬ��fb�	��V���gn�]
���~��������(��g�9�C=�+\��?��G������3m�6�[t��:��S#�ekŇ�� �ֲ[�Wvc5MRZ���5	�9G�1J��m�mz�7���{ӍRmf�sȮW���e��GyK&BqQZr���ۜrxH�K�T#���q�HHi�(Rw�H��o�)��9bkkN�p��y$���� a�(*�"+	����s�d���MgO������1h�����x�t�%O�S<Leͭ�¢��w��.��A�crN���]��ĥ��c���1)�\>�EY���� �Semi���b����T��-S��|(r�t�$�Œ����2�����	��7=�\��1Z�L����U'&����V~W$,g>:�em���Pj"�Ȕ���ә^���v~��������J=���*������F��{��� �1����P=
������>�g��e�k'[y���0��l�B;<$��>,&���RzAS���<���i���}b�Ӷ+��D�Td��_�'�!{�2\�=��S8�@5�0�9.~ɶ ����۶�A�w��]H�W~�_sY^4����w�����3>�=�Es�$r��,�T�{�&q>�T�Bn�/}��rŘ?������0���и#�D8�ԕ�YwqHk�aN����`u^�j��03s��U��ݍ��~m�0���M.��<�$%�jڏT0d�e���)T55�)�(��(����sB��Fh�R�h}���
B��:�������d�*�U��e�q���4o��W����
I�!x1 iቊ�����5��T`a)�xc��0k����ֆ�L�+|�5[hQZ@/�=�s�P)[�}/����|�\���c��b〬�*��D��8#C��Պ#���w+>?��{�H&R � Ɓպ���q��5(L���*�����2���CrO��з��I]C��~&��0|�'{"�q����0����d~��)x��ڻ�	������m[������y���,vV�7saQ��Q$Vl+2PV�����n��8���989�O����#��Ǒ�����?U�Z�o��f0��JqְJ7T&%�^����*����U���d��c�o�f����;����ÍJ�d�p��"q��`�yM0���^>b�p�t�5��`?��ړ��Rt�����۾�	V����\|���d��
6�������{�`-�+f4����`^�l7>��� ����d����+s%]����Z0.=��L-�F�;\�|q��O��w����ɧᗌ�@�r����!�����_�K�XE�ү�ƛ�*�n;Ʊ^}�H�#��N�o�-�ǹ�q\���������I��P]_&��s���&�s�c/�JCєd��b� �����袚�L��#u|S\I:&(}E=�����Ȣ?������/n:|Y��h��'G6�?D�D�?�o���|2��bΪ�?�t7�LY��1������E	��ci�F��{s7U7ް��w=�bv[��\0�aW�HU�����1��w����������!�'F��8$�O2�^��4���H"Q��� ����! �k��J�E˺G���Ҁք��$jA>��_�e�:�������QIA�3�Z�I�{:(�{d-�@~/��]���\�0RF؄@��]0cۅ嗙vB�K�|�[����������� ��?�y�MO����޲�[�2+�VY]�)��H�MwV���	��3<)3Y�����|�\4��E%�6qٮ6�ե=[6	�{M�rsԋh�5W������|�����Òsv���f��m0�i�]�d��R sƫ]{,3i~�*Ɲ�kr�J��j�c���
R0����u��R�F1�x&��f쀡6?�a%�s���i��a�><.#<��@E����Ҟ=7�KJa��n>�N��i?��X��~�������B�1Q�O����C�"����\��T�J���!̹H�.���s&~"�y&
(~筶mtՀ�\����"w
��X�0���Ru?�y����ʖ��Ձ��DLA��?݄�`VQ`��b�pϏM�c2'��,��[`�ѣr�\��4q4bb�4�Mh�(q£ڦ+�!��1���f�bIf��ל�^�7N��kgCg2d��������l�<��ᒳ8e�g��
n�r}���YB� ���觭X�����d�M�����q e8Hzl>�:9��Na2F�0s���a�@=v}bB�ۿi��@4r��)t`c^l����{�=�g�AΗډNM@���A��g���Z@�nM�G� ������#8œ$�BCj��6\Qš�������;Ok*X��a�t�;;�����~b_z�J~ҍ8t�����3!�Z�֞;�],� @�(z��F>���= �Ȇ�8J}�7�?\�[�Z�˔"���{�=ӝj[����OsuW	�Ys�o}Az�O�����ɖ���c?�jy^��Ր@Z�K�q��"`������]��L�H���̓�>#ƖM�ԇt3�9��������!�����A��4 �O����mؿuy�%���#�N���.e�?0wx��� %�ې�����z*� �z:����jQ3�oGdD�ʖR�#	�{9�t��WN�z��?��(_��'�0,j��UG�!{s0�ݎmy��v��lɁ�=�)1��\K#�ė�Lm&��ď���r����%�D$��M�GI�I�[_T?�
�4���*����<꿢 �+�^P�g�O,���Y4���OQ�����h��!����w|��͑<?�~���;�H{ĩ[�u�k+(�kO�5GkV�4��K���L��k+s�R�K��ܺ���+Ĭ�9C��$K���!�.]o7w��t��V�K�t��7�zW����7L�q{?�Ɵc4t(�.h��U��|������
��̏D'F���̛���v�jj���2��er��3q��P]��TD^�L��K� S�׵7��S`w��D���0���]��|>luծ��(qn��{B�5�x�����P�ue'$/e�� z�3BC��S*%���yP�GH�$>zT$U��Y���ƣB��3�>�*Ԥ�懁*�;Pqt��P�Tm3O�O� F�QKl���ø�1�I�Kl�)e���f5M�Y3g@C����zi��}��ϴT�N}d��:;`�+�׵�����������o�5t{#d��M�G"��
"X���\���P� ��L_>`���}T�1���ԡH;�����7rX9���k�&�D�����4�X������tn�v�r;�����k5��>�-�}Y��6��~����t�I���ן�؊��ϥZ��������D�Q,���M�P�D�����p�#�˘�{_Ю��89_|cd�zXP���@��/"��9�rʏ"xtSѹ����aJ���(�����x��R��|q���
/G��}a��ߠA�B���U{�E84
t��7�*��Ky�:�JX�4�w�����/���l`6]�I)�'��c�a)�J�M�6�
bn[�zt���SR�!?L�b��_k.M�o� !�m_�T!�VL���ں� �ۨ�PkD	�娀\y=�:�-Eta,�1����Ro:��Sױ7h�@�*���U�]f)u:�81�
�j[�%[K���v�-�W|��1�\�~�M����\:��	 +�s����`-�y��K��H�)�lәڴ�]���(\�Z}ɏ�Q�υ{~���Ѱ?�p9	`A<Fn;�U���R���6��LǪw�Rt1W���L5�N�q���6@B!���)wf����Iu:��B#nTs��re
����(���4j�'��e'.�,!&��\�%���ߴ�*��/�>nڲH40���>��� %w�՝>� �2(U�,��l��=vh�x���^�GIj$V��c�d9N�����1��>� ����/�����/�-�k��*C�!��a�Riצ� �>�����I�J���O�9�/��jb�c�TM�����;��&�e���Kp�N��;��Jpe\�.��ͫ�pobqw�D-��˚���2�� ��5�~��h�re����
���G4[��M%/,�ʫ�_%��B'φ��R�MX m-��[�u�>es�**S��d?F�͖�6cP���&��כ��p�f���E �u{J;�$)�Cߐ���n�.�-GU�p�`�j3��G�$,�r���������� �L�^%D���l�Xy��]�����y~�ޜ��
� �e���9$93��Z�nrm���lg�6��}��ӠsR�	��,���~v�J>��B_�ҡ(��ݢ��U^Չ����9S�?�Q����(�����sѓ��S�)6��z��c���X�6��
��O3� � �R���o��4u��a<2���ˎ͏�kOդ6���6B/�}���2HL'?��?���cĲxt)hp(]���- ��1�b�m�0{	,|ɯ��P}����y�Of��Þ�|:��M�5��=�dj"82Y�KT�6� ��84M;=W���3򟛡��F��"��'�<Ȕ}j�Y��n�1�xU�8|n��	=������}9/���	J� � �Ȅ�UFQs��À�o��3r3���|5�yU'��D��x�B���F��jB�|���a{c"Y�i��T�*�^�ֵH�t���z�q�Z��s�3�f,�?�dƺ�Nvu�����ْ���vݢ��&?�L�r�/����X�%��6���8�=�<zw?�m?v[�W��U���ac2u��ξ�m׊��	��W�����`��9T�q�昐 ��k�_\ݨp�[����Z�hó5�Y�:������HC�Z���T�GZ ��fk���}��Pw��p'��<���/l����X�A��{���Y-�H�C9ݔ=���j�8`�Ȏ����J��.�\����]@�vwN�UԫO��e`W|�&*Q��*��>��h�yoZ�:2�A���Ⱥ�z�3�^/� Ʒ�ae�@E��ռ۝�u�����F���t��A��ME#���J���=��d`�yvr8D�w���:,R�K!��R9;&�t��&���jN��e��N��~�D�2���^$�HԽ#��ve߯K%W�43��L
I�+*��(�)��c�
���������g�H�^B�~j$	;[x�p�?j�}�cX�~wQ�}������[m�[�ZƸ�9���ll�14}!L���,����m�2��,y��<�#)|��րnon�/x�x0(�b�`�
3_g!���t^���3�����m�x� �[d'ӓq�?�4DG�q���Ntmڋ�>`qJ��D�!�Y�XV��d\��'�у��`/��푬͈�ky��Z�����?�8�4�8�����_�����s1��\�s`^����!��~��f�n�ڄp�[������7��5�̊R,�X �H�¬����U�c+F�:g`�ᯐ-�L̡��q4���]�ۯ���۩0�����`j纒Dk�PPp:�%j�¥��Q`�H�B$)Z��Z =k����C�8
�4�7�驖<�|�&�	-����Q������\��Nx�ѥV{/�=�C��ܥ�C��ٺ���U�)W4	]A��L��
~w��&��@�v}��c�N�&vx���*�|�&�T�O�9��}WWtEa��Y���^U�<�ε��X�?�(9v��cf��
�cHb�'�)�bZ=@����
�<�X�������xc[��ԓ������M<+M�Ǯ�W���d R)L)���7t��� ���;dS�wی��!u���ˋ�'S7];io��t��vV(p.,�ո=��I,N���}|/iXaq�S�����������$�����Rt��pY`oaD����[!��N��h(|�=3@��0�\�\&~uT��r*�{��n������>D�7�N�}�'C�����jz��"����|-4�/,�E��`�l�B�5��:��j�G���-�����2*�:��(�x@Hjf��G����H=����Z1�p��Kبl3%�3rd�Ý�#8U|���W	�x�?���f�KJ��&��*��A0�+���+Co�������]DTő��ˊ�d���A�.��-�Y���Q��c��ԇU-��*��&*%���`8������+/�6��C���_�>>b=V�w��w����s��P�^4k+�3W��$m��WNu�mT4e���e��\���ͪ�e��ϴ��@��yL=�[���ҙ��5!��I1և�[��:Bu��L��rW��`d��]���im�}%�/PI��3Bi�_Q�|��N��6�L}�x��ǲ��֧��m4/�N4`D��1R�]���sI�l��=F�EQ�������RĦQ\��&�����D�4M��`]p[���G���g����"Z5�sp)d���}��ڬN�+tR<}4���bu&@�{����	�zA���N�h&G�����X�ˁ�P����&:�_�j��h~�3j�z;r�]֣/Ib��K��`G,}�,���������,�v��h����1�~�y_���� ��s��>W�gm��d�
:�'����E]�L�����p<�t;7E�#��*�2�G�K��-���U�����}/7�j��~�,m0�KD ~�L�/�_�v����&�j�3$�'o��ԭ){�o�;��|�r+�%�	0b>\��u�4϶�dE��*�S��y�X\{��E7���*+.5��<�©�u�E^���%��:R���+���u�]��g�`���E1-#ʮS���F�2�������\!��$�i�#Jn�.!Q����<���U�E&���M�:����eC�J�+�yV1�xU٤��*��y*Mݛ�9�f*�g�^Ȗ�RN�%aJ�J"�Ŕ�1*�s6��Z�Kg÷���.�����E��ivp>�YM��q��(�Gz�f�F*�G�mZ�;��W�b�-�,CL~�׋r%CR=�/(%B_�K�?{ג�$��BN��|��������~ii����e�̙ɞ������c��!��ߋ��gF8�Ҭ�g[Q�O0��hf:đ����*�^��-�y��S_�rB
�V�Bo���[++-�كԃ+�u�݄aa�.:\��*IF?i%wP��f: ��ٞ�~|3���Gg/Ϩm<
�ev���i��� U����!ҺL�&��&�Q�Bm�#g�2m�t}��Xzf�BT\�ߋ$Dqނ��mࢬ^���I����g�*�%���U�&>��.��G2H*�_�.FD�4n{�k�3�y>�L�ȧ��	�3�M�P�;n	t͑�[��!�&! V�T�9���P���B�r�4F�]-�S�^}O�NK��s(��aT�e@�7,��	������nb��bE�:5y�Z*ֆ	i��\�a��qe7�cgd�kjR�{��Y}�U�Ԡ���Dp�S�I�a>O,H���%�|Y�\��#��7.��J|z��Gm�ջ��FQYwd���2L�a+x��0�oyxT�"����b��-��5m*�����ksFS�
z\f}��Eӏ��)5XhI*�3H��6���m#h� '``��Se��n�ç���1�f�O, ����fg�e��o淪v������j�I�0 �yS��z��d�	��趪�����@�r���.�0K�%�Ḃ!����F���;B.�Vڑo��^K���H�)�Ԡ�&��{,YN�7���A��t�:i����}>zt�؝0��	�74+�E`��2R���#�d��C.5���^h���u^�������*���!j�9؊U�ֽRFm���3k_������:'`����K+���2���0b�����a--h?��]���*`9��4�Q^_�A�A�|~�ǐ��(�Pa�����	�w7{-f+'-';δ�|[�|6{�J��8�C�g��Y+a>)#��|��.'������΀�'87��n8�an�2�2�]B	,A�ҩ��-���(�#��!^�"��-�����g�:�m�g؀�N~�F�͞^ђ)������L�R/��z���U�-��j�~g��-qUe��l�54�[����:�`a������b�B���u�����|��î�a��9�F�S;�5�wk�c��Z�^�Ԙ$�d�K���u�2*`oٴ;~��W&t��E��%ȟE�9�!�a�7�ܤQ3#�D��uNJz����{��i���$	)��2�iO�'��΋�?��Ő-8�����g}%�P!��)�����B��bJ^B�����3��B��ډ͊o�7�n[�p�
=���4�����x�<��0�Cw�E�"!�o�Y2N�=�a)6+y�o�(���^Y��Y��x�6�F20��lآ�އ^�̄HC�BL
p�S�|m/�Ű�b�9=��^���,
 zm����kYV��w���Aa=�@���30�����xϙ��UD_^m�`1�L �S?f���n�Ò�s
cI�kW�P�cȶ�зzK�v3��jqM|����W��O$
�Em���I�^�-��%��f��)��7M�j!�Tg��O]���O�aG^�3�~�F�qEQ�;�&�M�����s��4�n���_��쑲x��g6#��쟖�j�X=��=Ŏ��_q�X;Т�$���f��⛇���vcJo��Uϕ��K��*��m�
�'�т�S	���e��0�JL�?z��gd;=e[��̠���`P��p�y^DL�I�M'5W�����k��qs�� �3�4_�NOT�H��EO��S��b�x�To����l颋XH�v�?���fF���|XQ�� ב,�GǞ�>Mǖ�u��`����>!	x_��Z��7�ꚂAW{	��/JG.��b/ܬ�N���o�Z�~�"��ʻ��BtK�����kJ��k�% �9U8W^�D��ڞI�a�R Y��*�)�-܈0Idr�C�4���qf��tId�䙛�F3&�!YZ'�~�lI��9�h��� ,y�p�(AMu^������r�Yy��*���`bk�{�B27�����F�S�Sl�
_}�:��%Uk��"��˂k2:Jj��/6UC�l���~+f�5��m��F��.� ��ت�}�ΐ;zy�-(JQ�ŵ�~�������$},xW�|�<S�b�'!����F7@G��j>P~\�����ⶵ�_�"�d�2pk`f��_'��#��H`,BуK�m@��~��?O1����_�+I<�x�	z���͋K�ʦ�?��c+���#������r2w�1ٛ�;��=�d��SXnp�A)�[�o�����_?��+�`Ν4z5�2J��q^K�)d�;Ž����
}�M�t�ӭ>�6m�
���ȯQ�?�m��5��j����Mᥴ�z��]{��{�+�EP���c���Z0B1��c���!ǵ8y1匨�(��۷@H{HR"PP����G}�j�x w8i\��+�4u1�4�ѻv�:��FY�>����M%�l��?�;!DH4b��g٤�KP�'�����4L��j��îƒ��$}��5W�t=�tW'�������oRݧ��Q?���7�,�z��&��M�b�J�hV��ycU�#� X�����A6��� �p�%u�Y+P��ڡ��7Ӕ��"�Y�3�x(K�Ԓ;XyP98��a�����x���.�<�!�6�m�@��k�����+p*.�/ˉ�r��1�����O\nx�-����	�E�y��:�F��eN��Y�����e �..+�b-<�Ѹ#�m�i�Z�.TŰ� �a�*�?��%���ȍb8�bT�2u)�Gm�Źe2�(g�"��a>g����z�X�f����$�[��<+��	b���n����$�[]����Z�h�g�K�#�/%�l"������nd���4�|�m��]���%�#؀���f	^���_)̗�@��,b&��MM�$��� �!\Sϖ�ऌ����A0l�� ��,��ad���4F�;EEi5������a���9��<���鵜�lxZN�:o���+T��xPJB(�C��9>`l:�AaU�s��n�"���X����.K�=�՚��ׁd��A���~7u&~I�~f`(\F���ɚ�X��~�\ܫ|>�r��0B�W�Z���[����>�j��S�=͌��Rg(�=�?aUr���t@�c�eW�O!�g�dݫ>��Dn[u ܦG��!=(���>.�D�1c���+��"�����ZA���>�-���OX�ٹ�c�B���pE}���z� �|h��Гgp0�-)�M�t���#�{$~cw롆�����#�B��V�Uoм�g[bfm�bm�*ׄ�����@����� ��͞���.��٨��cR���.��Cʷ���<�5��6���x> �]��T9��w�E���J�������N��k�L�"/��e������5=�76'�e��U��|�*#=�e�W@�aU��]��D�V>���Hd*MbvL؀�/�O��7��3�4Hf���>�)���(Du�筏�UA>: �����k����%1�M���ѲOM��cBD�Y�	9���軲�3P�]����E`f���mr#��@�qJ?��� H��p]N�-kx{��X����:ru��ZJ~�\�LO��M;��处�:�{�]W��.6{�A�P���a?濊m�>�6>"V����TN���B:Ĺ��W��l��ǭ:A�;�#�e*����F�*"N�̛>�x��3�e�����Y��,d�ԒH���=�NA�t?�]���<�ϮG|����J�m�6l��3��b���R@!��׼�ޥ�w)�>�m�����z�xL98O�����W*�٭�������곶륢�ϔ���8<`HxC�*!�6����y�Io?��R�ږV�g��n���ϤO&�3.��
�gl���@���(*t{k`�r�x�Sf%ص�SEK>�#'���>�h��ЈU�g�ܶ�  ��8䆹�����$�8|��խs[�R�'���|���	�� O�!�9�� ���m��<h��]���pu�E���9�
��'��Q�I�ݐ�>��Q�w.�aR���5��~q�*�<��+����u�U�Ox첳Vr����5yc.�$/d��S�.:[�zZ�J̦��7t�K�_N*��%�2���>��v��0ݍ'�4^�`#C7�y����ݼ�P��	N�w3[})�P�#�'AZ3+��#�5a��U������w����;����8w��%0S\ ���iݗz�`��֫���2�����F��Fi�JiHŲO���kr�.�,��}�2]}W�bw+��@�����m�LݳM����bx�xE�-�$q�{w�-�rN��~�Ч���{,2�
C6�!��������i���Q*�T�hY��G!�t��k"3 O�ұy]��O$��C��1$ �J�=C��z�M+@���k�v�;�4���C��R5_�N��n���a�dC8�Գ6�JՒhQ��_�bP��U5(��XΞ[��7��ވ�V�G`�������n�T߿o�I��r��`�F4�⣌��Ґx>.���xr,z��x�uY%��)bQes�.:�{�x��b���mJ�#,/g�ѹrNʍ=F�ǉ����S�'}�ِ��v�����	�0�u�o��x���VN��a>���������m��rF��g�!�X��iDevIc;����נѲ���k!(�1X��o<��Y6�Q�˘�X���A;02k��/*7p6"��0��zC>�W�R<ѳ�`�T���K�S�g!���jӴ���_"�R��ַk0���{�C�QP�"p"���IE���T�����t�\�ܯ[���᛼Ĕ�&��f8�_����u%}�+@��0/��U���Y�����9�dn���?g��R�0�z!kE�2��4�.!� <(�5@�&CE6�"�#�E"��- _����>b�Wg%�o2�lzr��>_��f\��:�p�L���-(�d@�\beɖ�f>�';a�z|�(�ş�^����< ��i/`�=wl+ �H�Cf�?�[}P��ܖ��H����[�/1�z�GjK��K��F���s�j?|婤�D�[�&~�2��e�i}/+/x�>KD�F˼z�t�I���M�^�XJm��R�ur%��,#/?G������K^�5�ߨ�C껝oJS�nJx�8S���aK�0��I�VY��=�u�z.%:_��m�������e/FTk�.�q���T@{�.:Pސd�� �㟤M�f�uw��!G7V�))��B�O���z	*[@�a����#�C�8g�����<�qyx<�V���?�ᵄYR��>�������x5ˑ�ofΤC�f��V=��ZO^�V� aY9���j�1>2K��*�F&�� ����ƅ���h���R�;�����>�ُ+�w��t��'�7�����3܌>��9@<5�qm)��y�&�/�R�U.O1]�\!�e�W"�JN�^kHĴ*��e��r��>Ld*�Z�N=t���T-Ͱ�{�p�|����G�Y��Q��`O���|��{�(t�o���ڻoÎ����H  ��GsT�o��$(I����J]^��Z�m�&�����6Ce�;���N��8O�xD���X(�X8G�cO�9��a�u<��?=d`����W���f�sCP��ȡ�+\a,GNu�������Ӯ����
+�/�oV��dU����G�=-Q%�(����ͽ�v�%����Y�/��h�(��[l=)���?���Xs}LGgm��/L #�	L՜ϖ�ag[71���^���1|L�����d��� ��0�s�>�4.d���C��I@�75U���<�91�󝋋���c�z��p<)�!�G�G�A�m/XH��)��>7���!�&x�X�,}���-���9���}3�4^i%5��^�58�6uQ*�X����"����#fn��#�J}%c8H?�t�ێł���Wl��,*n4�K���M�%�+��n$?���� �޾`4{�<�@� ;EQKy�-"G�6���'��5�#����W�=���P��ً�<&�����t9��aR�F���4j�-Z����KP��*3�k [���9�X�/emn뚦�܈4�"�0�������;�d���p��5��x���☛��? �S�f�vq �(Î���?�o���E�����"�+=�C	=�{w��V�!�y>P���b*��y�_�j"=\lgY���BB/?O���ʧHbÕ��|�Nf��3>s�V�77������lT6��W�<�x�]ϯ�������	��p�<���y�@���Ֆ$����D�ðy�R�D���HH��:NG��zH!X�}6�H{)��v�V���9@���f�t�@�zo=��)Ɔ���M������NK��B�=ί���Bo#i�R]�e׳���"t�y��ܓ4��%�U�Oz�_@P+>\jD�J�Wr�#��7 ���J	פE4W��0�|ҟ?n�����������d�J��E�E����
� ,ǛrW�-Ad�}��F���E:��o`�3��YK!������m��������$KX��ܑw�..H�������^��ֶݭyR�P�r�Ӊ�^���׽M����z��O��=շ����<o��G-��C?�������S�1�c]�~:+L�pᶕ��Y�o�*�rI,J �P#������t9)��y��z� #��llD\���P75@�=�l���KR��y�C�G.W=ZVtj2T����hw.���+C}�8C����=m�\ݤ��g�4�K�xbz���)��*�iX�æ��6V#����L=ܚ5Q?���xl�������/	u��ǛR��Ô}n�����,�R�dQ�{1I��Ranp5��a�@�g��h�f=������K-��v�Z���V���br�.�#O�`�.y~��%���Qh�0�d��I���A�7�f}`!�["����p�,^(���}��kV3����Yd��R,L�h�㬐;L�^",���N'(�.���j��Ȣ���,��9�8�ϟQ�o����n��<�) �e��$�C�VA�+��G�x>�jL��&xǾ�T�Zʆ⌋�#��N#��t��`+hskE�F������[VO!h��F�� ��ap�;n:�G��iJŶ���;9�&���o�Z��p�x�a�I6@�i�q���2;�_�"�;��=(Z�ÖV��Z�, |�T�-�9��I��Έާ:�d5$�� ��,J�-qz��H�#�-������B�<����v@Z�7Y��liy�ش�KS�A�d�9�����KZ�� �B���*�r['s�đ�|�g�ԡ�g�3Vgs�_� ��K�7�=ێ�
�>bے"پp��<�tu�_wln[��bCđ4�i���)�[M�lX[��A��D�֜���)]l+	���3��$~ QY�z>	����4��mZ��*����s�^V�����(����͈�:�EW�I�Ǜ@f����[�fu����ɎU�@tZ�K��vKy�fF�R̶��sI8ɷe^�i�S���dU���-_S�6i�y�����Ϛ��!>�Yu�z�}s��{����w)�����͡�N� �M	�)�
��7�76W{L抻ak��6��f�q�4W_���!�W�� ���sc-�P�(��I᝘��&I.q7�ؾ;�����%��`�Ӡ���2�mJQ���"q���D[��1�I�Lġ�|Ĝ�����+�I;16�r.�0�v�g9bV.����<�Ȧ	�{!j��f��J����V=ؗY��1�f��2y��XG�֍2K$a�y�̹�ʕ/J�4���K�rZ����!���XL�3W����Jؑ_�J춁���H	��z�]��ו"�Rpu�~�CY�pld�\�rH�m��� H6�mw<�V^�rU�/zō'��UK>�J��L\3��)~��p�R0J�$\�$�[qx~�>ȀhBv����ș1 )_�������3�6�K�Ϸ�՘�Ń��}�Q|�T*k�Jq��W�c�<2�8��=�"ֈ%�����g��IƑ�O6
s�u�7��W] �`�u-�~J����<��}���c�psY��}�B�b��	�X������I�\�Ԫ��|e���w
�On���uj*&s4,i��h[b]����L��m�,H���
�-�i�J����ϸY_�-�c�\�%k�S=������f坶:1��R�����؀�"J��A��N}�P�����h�IG'�>Fш�O�&<P��bj6�����j�Ҽ>J��JURON>f�^�c���zJJ�dOr8XP��f��%��!��m?[��_����ϮQ�n��`�/�2]\��t
As5'N?������f��#QS�Ā����CC�7D ��$}�X�V�L�q`�C�:҈���<*��`08>�B�T����S��ƈ�����Ų���6�0��nMx`�Yit?���� ��bȯ8�ᔥ��y�'�:-�<�~�������5�R����ǭ��ó�ѩ2�P
Y��0�y|@����$ܨ㒱��N��z!������mV������<؇w�@�R�ؑ���V�,��vk�Dܘ�n_�h�I52X���/�s��5"c�kg�Bs��ގ��N���>����F���i�~�A|��M�Q�1�<Y�f�*��[/��'�ܯQ�~U�'_��� �	
��·8�7� �8J�5$V��&@��� ?%ũ�`�������T�2���;�A?�E�������4z~C�����S��2���#)���Hi�(~V?y��e��v��ʰ��H�~���(�^�Ӿ��R�h�`�8�K��ހ��7J+g-?��[�CJ8�dU�5^��)bc�8��vb"�u��"o��%�S�����O�k+�]u�{/N��~�5'L�f�^.�Ԝ�וTF��]a����#�Y�/_�����5�*�>r�U���B\����t?.��	(B���᫕;�Z�P��kD���m\��W܏�;�Y��[������^�҉�8�}�c��(��g��'@m��� %`'�4
j��|���IZh 1��1WW�;�����J�eO�Q���4 �����Aȿ\�V<���i"-7  �� S�V5N�2@4YZLs����<=U�����k������+���ɷsv<�����MY폤k��]�#x����cp��j���ΰi��)�TC46�嶫�I����,��y�GK-#H�yy ����`�]�;=iweNNݒ����߱�V�*9w���{�Ex��7��I_-k��-����s��)��ܗ��uy
(A�$���W_�����c�=ѝ�s�	��.C-�Y�$�ѡ��.^M���O������wZ����-�d���
q�b�Yc���nyz ;��n�aζ��,޵���,'� �l�ෲ0!���K��gE���NF5w� �L�9�o?���A2ӴkoP��B�k��xka��̢{?"yզ��)�� Mg����[���F�(}y�i�'�#9��<f�� t�x��\m??�)o��d�p�d�/�[i{�4TU `[8�~� E2��*'Ԗ��
�c|�}s��s�h8|�>�w��Κn8{�T}����I��/�s[L���F�VH�������F�n�z���k�DH6oɆ�8�Sޔ�N������R�����/Q�5F��L�lAO����	��ÂkC=�y?Y��{O��έ�V"h��ƺz��e�%H�9�A/�rx~n��-"���ܚ��]�(34u��SI�bk|S[%�L^d${���hY�m���$������n�ʘ�@q�h	�(�S��"�4� -��d��D��N ����0+�F�B%4%��?��~��	\������G��,�����|��A36-EhUHuH�͈��[*�Վ�S<(_P�X{��{t�o�9�� ^C��ھ�&Ho1��{R@��xZR��2�@v��^�o'�/��H���A��js����0���8+{s���@���45灢�7$���U�f���t�W8�Բ'"�N� �t�:i5��[�0�2!8#��?kݺ��I��g�L���[Ԓ{}8���,A!t�L�2c�l���8��]��vWq$p���/#x�%ێ�ջ��!n2� �;\�ħ����,l���I)��g�/��������m\�[���`���U�R�*����dǭJN���s	�g�.��g��K�T�7��.��R�N��`�d��pl*��Jj��`wj��������$; K�(8*%��XҼ���HLȿM�P%Ty���a��/0���� �qw�rN��\�Ƃ�Z��x�eY�v�������
Gb76����/�4Ο[�ڼ��Qs|[��$^a�E��ޢs��i^�<׈��#v/��؛�z6��ֶ��i�z�2r�m���T��C�~�vK'���"�9.n�&C:�[�F?>�Z�Se0 ,f�G** ;@k7<�zhdu,[�id�#Qh����^��S=�D�(�AXp�����-�̢��o��9'��������To՜�}���(idž���k�>'�����? ��k؂~�5nc���F�8��Q�s�'������.��ڌ~_m��04fk�6�U�OS@�F`L^h��<�����rɥ�O��^������Y��o'�t;ƶ~��Q��֑q����(C�7<� �h��-�XU�Ϛ����G�0������#θ�����~\�`��޵��ZR�?B��I3�)t�c�Es4�al,2�Ch'���M�+�q��

�o�V(1����K��tF����:�r����@�8�Ö�eũ��#��:+���#����0��z=H�&n�e��&����2B[^j$�_+�V7gl�Ѓo��CR�Ʊ�j�����ZF�2�Y�{TW��?�ӗ�%2�����K��K�� �i`���~�_���g.Q.�Ś�4dKS31xy8� ��؋H>�xR;x�
�U��f���IH�l_��m����D��ĉ'��:���y@v ��Ý���?�U�Mi*��D�0��W��l4�:�����G�����k����7�&�U���+R��D�d�9�<})ٰ{{f}uڒp�r�d�uV�QP�˙6go&zt�ED�E��B��әWo���@��b>�$%���Y[ҼD'Y#�1�p�>y؀��)�}���d�K�s�A<���~iWn��r=1qb`J�B2�:F;���Pc��}T�)�Z�6aC�pRLH�����Im����~�n��r>?�{�t�p=>u�j��EҬ.�Ɍ,&�)���&M�"�;��
c*�*Ί��WW��$>񱅮�A�	ݪ��tJ���GXk{�)�_��T��UcC�!1���&'�t ��;֙vܓ��vAyzl�ճ=�ށ�c��U��64J��=ZMnG[���kL�hX�J<?��|RXS?���:?�8��v?F!$-�'V�TȬJmu�!dW�%�Cb �|�'ص��{H�3�j2�5�0�5�|����<�ݘ�гQ{)��%�t���TK��v��D����c����zd�u��/S'���6S=�u��U��y��z-�㍯h|�c���>oO�Dt?:�PJ�����3����[_�U�+Ǟ�#�I�=�jc<DקN=�#3�=}~ �ƹ� �|,�3A3M.U��$^�<!ok��5���p[��g�ڷ�h���xqa��gALKꕥ�E�����i��>7J���g��z����]��������Yc��\2���3y�D�q�Ǥ �I�+U��aՓFȂ3K�i��m�~Bp��t=٠�t�9`�K,���e�����\���2 �0��*�yO��
Ph�\�U�Ex�#z�� �/��
��������+�A�]�|Ā�r�(kPgu�k� �R�Ą�C_%8��0�?ۜ�g��"�-sJ��)&2�K�I�ΝE��3t��<���L��uj�6�&<������=gp��.b�'y�c��NM�'i��I6J�O��p��̩d>��̙e*G2�v���=a���3�B�V��'L隉�+��x�|Ghl_/��J�����������3.]Ta1ba�l�b	&+"��p`��3�b�&ޫ�MX�Q ��]�VZ�/�:��$��AE��@T��#,zq���1?�y���=[�s��������SBZ�W!���͋�~nH*�?�sR`����<"�%g�%Ҋ��U�*���˵�/��o4��[�u�?�j��rr0�s���3�?��|����� H^&�8�,u�i�Wy��?9bw�c$�
Y>(FW���`�x&�׍Yӿ�Q=����rR[�M��
\�cجU$�S�7�G����!^�}������-�r]��1�;���n����8�/@Ӌ`���"b��[���o�v�D���8�T��&����A�	uh��t�Z�V2Rf�Y��ľ��/\;*�r�W�ɐ.��%@]�H"E���u��i�͑��5,�!_
�������q涉N�8n+�5�	�����Q=z�EW'U47�vu�0�_YDǣ�LE�{	��r%K2)O"��JtUC�Pe�RԌ_}/v��}�~%��s�"~2	�{��E�'O���Z��z1Mo�ڸ!�w����\�_�?�(�qh�]��k���	L�)g�{�a�'�-�ߖ�'p�4G�J<�Kh��+JT�p���1��kG/���v��y3��~)[?�`Q,&�A��uq/7?5�![�
���4�S�H�O�ܝѱT��w����[�'�����"8��-K!�6[����+�e���jmY��󰲇�a��{EFbG�%:]����.v��d���뇲.��A-���<@�����2<���k$��᧨O�ccD���I��wa��0���נ��&�G4o��^�>2ut�8H��@Z�!�����GB ��S��Fk�$� y�M��]S������f\�Rգ5cϗEƮ�ߩ�p�%�{��h�M=��>v�w�$���潶�����m��G7�L���|ѻW�]�{y��q���W���֐����� �w�x4t�SK?�Hu��Ar;m�=�!��g^EHZ7rmCߨ�. -T�Ў�u)7o��u6�bF��UR�+����Y���X�'�]�z�K+ơ=�v����*
��o���\t�&W���H*u���!�}5�U���J��1�</��Ed&�(�0��࿹����Ԃ�-n�,$e�y!-x���Z	d�0��4�ʑ%7Qn���Wx�/�'x|D��#��O-��j�+�����H�=�Ä��$��~ � ?P�#���"��1�#f���NU������n�E��3�џ�J.�[�dk� {������|�x�L$��(�j�����ZH���O�d�)ӆq����2�`3Z��-צ�t(�FX���G��c�Jy�+ �ݨ�){F�r]�2���?�n%<�rٳB�?�,���xs�mA�k��$fkv�zG'IR��?Y5���H+[F��}�����*������p�u�1��G"Ļ��^�g�A\������)����L�q���6��\��@@h���J{�NuY{p6/�]`i�oa��1 ~RąKXpH��3Nvi]%l�0"���b5�ul��~�˵����!�s�Lq�J��]n�Z��%��Յ�˝(��'�2���*��%�|K��߈̴�ZIR��"����tZ}�Ҟ�q)�<���[&ٸ�|�x!N�ݛ��3���@ȱ-�l+���G|3h���#��$��CAw����n���5�Uʨ]9�K�X�r��ܙ� 7���>U����}����Y�լNHx�#?88����7[�K�`��9z�/-�g���ӥ�:6�c��7.���)*�}�Wu�Ybݸ�ߒ����t�a�~�25^�
�����[�')�JQ�����	śǑ�tz��K����\�6	��(����]�XQ<7J��$��E48��s$�4����jiȭ��>R����>ed8j��@�m��3?���g�_� ��
d��W��t���Ǽԟ,(�eբ��0\�Kf� ኴ��v`ȏ�[�z���,��W>$ ^
Z\o�@�,h看P�S4"r��PG��E�'js^�{��:��&av^�I�K�P�S��¦�� �ސ
��4'��B_�W"Ԧ�=��NH�fe�&��R#��c��>�C�JnL�����.9-M9k�?ꄳ���p�Yp)���՟g�d
2r�{��"��-�@h������<�IJ��a��ƴl*�NN�I��G�Ҫ�w��K��B"���~DZ1�c�>�<@�S9קK�M&�8��b�N,��v^g �J�[A����p(��=�m��~/ڦ}GJ�b<�:5X�7�v��j���dY8�=�q �H�hɮ���� �qd�Xo	(�Uk��^T�u��
B�6��<B��ĭ��Y�&����Yɚ���:��(,��f�"�����Vܰ�YB�s8������O�j,3>�SeC?^هx؊�8h7RA�Q&M[��
�#�kTGP��¿�+h��2m&������0�j )p��GO�|~P`ݿƢy^y��VdJ���a�p�r�ΙA�c��G<z�ۃ���i,t��I����+Z*��R���ǽk;��lhq�[6�
�
��C_c%R�wv�_
�[��z��h����2ިq�V���Sq�ͤ3�q~�[�f�ɭ(pU��\1t�1�-Ir��r��,��F�ڢfs�j�b��&e:T߀ZquL��2�(���bR�ue����(O|�����J!CL�W�!�{S�C�L��)��=����<�� *.	�C])�.�Ə�#��i�jX=���ɽ�X| c�T��Ln�,5^tƊ���ӿ��.��l?�����e�b:�r�1�����I>�\l�k$��M�1�w7Cct1Z��$Y� `d�|�ci�4�^��t��ҶB���	T�>[8O"��)5� |x���GK����`�x������	+������F����j�̣7��w�:L�B�~a:�2��ޑ8��L��s׃Ҙ
�}�k����T|��R|��~R�n��f��^<2��`��L���Zƣe�C�ʆ2<L6}s�$�t^�=-���߅���{�C��T{����|[Cc�	n{��'pA��s�{x�vor��H��#\yk9k�GĈ�Ɍ�u������~5&�^��\c�a���'}zKƮ}U��Ǎ�֭`6ֳ'T��RT�]��>����E�r�É��N�O}��7�o �c�!�/��|�>|���I#�N	�>vJU�,�92W�y�P0�~#��)�Op�g��Dk ׳�媙��G1��PNx!�]��%�=�Y���. �4@"��Fn_9�](�Ϲ�)7u��F�R�, <;WZ�U]\�u��)5����e��&7;�7��6�+��5jAkm��F+;��������{�B�\�'�1�YT3�4����]E�Z�������Z;�.~N�D�-[�����\�GRPs3G�O��aC�!���KB@���u?o3�~����;C1z�7s7�A�A;���?�:�ħ��nS6����2u�B1o���n�=�[��s��Uu�{����)�àj{1�1�Y���l�	W�5���l�@;�_��`���trW<��.�Q�u�W:��΢m�{��Ut��4d���� V��h��4��Sԣ�,x%��nn.�&�:�o�>�;�m{ C����,h���.PYǌ���.dN?`z�X����b�E�m.GA�T�&Mj W;�_�,!1�#P�����A�I�}��M���XQ3",��K�?Q?7\4	Ӕ|��ʣx�1��p�5�G�xb�&SBT�=��:��qĜ�iL�7���kmo��j�_x�E73=��g7�Tk��2�Vל��gh�=Ql�
�͖��G��d5�!�<bQ���m���%��s��D3�oN�˷�:bSu���a��nL�����AM_��aB ��Hl��)ur��,z�pb�w{��TJm]��w�8�v�5(��f(h#\����N	ʍ�0Y�W%�Oc�. �������ղ��-5�>*r�r�ADFv�����L���M	�āf<���Y�DI��v���	x���g$��7���ΠҚvS�I��*������--'��-�K��>H�`�����}���J���6����S�����,��A���!��_��6%�Q��?U;�	��L^���zW���b/�'�.1����
QZ�y���μ|�;�3m%��8խ,�D�5J��ٸԯ!�v���CWm��C2*M�����1��si����ס���C��x�U;&��Z<Lëo%z��:�8S�P�@5��[��uY]�j6���_�U`xY� NL�&��.R�L�`��A*��Rn�V��oُ�OX�3�v����W�n�`vτ�C26��N쉆$A��q�kw@��%�����f� M�ؗ"�b�a��H?D��y}~�ǐ�<����:�߶�$[���ad8�-;<;���Sn�>��D��*��#vJx2mI����+{�������o�Aw�/Ϳ�p.*�*�@�(Ci��7�k-n]�L��duu��W�>��v��7�Hx�s���]$u�V%w+uW�Hq�m�gLc2�U�wx�1�7������p���/<C��߸tU��
U���M܀����Nv�w��� ���u�u���G491%��sŽ	�_	x�|X��q�]��Zޅ݌��������v��V,�]ۤ	^��s�y�EN�h׏L�I�$�Jm�.b����!hr������Rޕ�S:4������WMȎ?rN��_��=#&���ϣ�&0M���iu
�E	l(u��Xn`�P�����plNiK�%�͂�����=��i	o�s3�g�4�*�	ՓKw�s��y�Ql+�$�;�:�R�=���r�z�:������U�9I�u�p|���ɔT�q�i���V���p��#U�mj��!��D�>/V뀽l�4D�3��
k��É)�����e%����U蘾ȫ<$���{��Tz8�T���6fDQ�@4�v�#���L�ro��ѓ,��I;@�+����9�'��v8j�R�h8o� �?�,[d�o
O�׼�4%�`r�п���=�tFJرOE����z��g�\`�덴ƚ�yٯ�|��~>]T<��TZmB��������
�gX�9�e~�o_��PH�J5z��Wn����h�-��^3��qi�jБ�S��L'В��8�a����$X5˞?!�{Igt0"w�\�������@]s�h"0����g�tq��L�����9��z���/�
c�8r39��(p~�arJI~2@u�F��+^A�W/m��v��_�5�ư^U�M�O��4�],3�څ��bu�>�����Ԗ[��j�,(^�|�JDNͣY�������������N��a�'�����|h]i����E����3�=�Be,"�?�1�0B̜Q���:6�	Z�����+f*��1���~�� �ЋϵT+qĨ�,%3�Hr���>��v����X'+�^� �Lq��$���c@X�����
,��Ñf~i��F{�6rke���;�3�9��1P��՗���9�%p�סd� F6�hG"_�/c�m��[eR@�����(�f� n��4�X��_~���>�C��|��Ό熨{���Y������������>g�Q2��xe��P��o[Q"z������`L���Ɣ�oK���j��Z'U���,s�CN�Wt#Ƚ�����?"�rrQ� pU,���j˩V@ȥ��f9�r}�m�!\|�Xͦ�8��k���DF��F� n��2/��q��OӐ`���uY�(�۴R��pw��5Z�bbͲk��u�~:n��N+Z�%���䖉�_��F��X*��IU�+�|E��{��*��aڷ�"�h|W.~�}ǥr�ʖ�����Iq��8�'{�1,|�/u� F�6�_q����nv�L��`�Gh"�F�T ҃����~հ�*v��\�(�aP�P�~6 X��9�Q����4J}��w�Ak2@I�w�T��>,��ډ-�Xڥ|6u���9�X}Z�9Sh�_���DY7��;��"�qW�	�zv��ճ+����'�@��V��ja�0�7��G$��ѨSB�q ^=�Tx�t�@A�-@mY���٥W�M�$5�n�?�4�6�gG8m�{���l�"�� ���@��nW�$�y��Z�@©b�르���D��N)-�F�j0R��Q
d�m[7�����Y,�2Q���9�[O�h�0Ԅo��*�i,W-�AT���������YZ�۴����ؾ���S��OPN`���@�`�6V�Pc�s�@�ǟ\�=�f�p��/t�]M�6h�,�o�Z t�08Cc�⧩yY��Oc�HM���z�8!��
��78]Q��0��wXCL`r�&�~ĉ���l���l&����ߓ0�f84ȹ]y�a�s�R|�&긭�WX�(+D?���
��ѵ�_���]`++�n�n��W��Y�ݚ�������n,pj,�&��j|*`�����wNF�rE�9ݐJsG��f>Qt��I�XC���K�/U�.��,��d@/���N���qa����ci++-�;8�~�d��<Qn��-�.�w	��c���`P�L����+1Yb�Y��=Y<)��pwv��o��b�K;�6��tLɁ��:3:NwmIn����:ր��8BȞe����Xe<K���WJ7�qT�z�����mo
����HE��'��W�ȅЃ������w*��.���)�]~��g����9�3J�����2D��hC�c�P�r�n�a�}�;�c�jWO�0�~�65�*�@�"�U�d��BV�R���r���E4Ԙ,�<���Dr��)��J9=�~: ��kJx��=���ʯ��mI	�^�P>E7��5pO����a�<��O:ifψD�d���p�ljZ��s���y��D��ea�ЙZ��`%Z�'�>�E�~p��dfg�W�G��$n�'�FW��=�,��lQ|t[*KkB<���E�pb>/Jm5v�W�\^m�6�Τ`��'5��a������CN�	����z`U�����-���!�����/���M�RB;��Y����(p aY�ߝIĈ�ӆd�s�+�s՟���Po$Z��\35+8��*v�8�����ɏ�^D^$�ݗ����Z�9)w���%f�� ��H�17���jՅKޟ�%U���KT�)F��5	�F���|�sֈ���+ L���o�|I��^�e��?��Qm��W�(VzX0�sx(�)|������I�H�=0��y���T�R�zK��l�0��o98TӮ����s��S"7ِ �#�$��lƜ嘢eD��)=zс�=�m?������ic�<�s��'�-��,�W&vr��Rt4�%���l��,!`B���}'�H�I����F�)_&��j�ެ�e@I�"���=Q1�TȠ����T�#r�!��Xɖ�	ಋ���7�q=��x��&���Q�n!�	a����J�}���y�~3G�L����d�F�}��k�5 ���A���Bi��ۼ"%*�
������S�c�k�M�K��D�i��Ʉ</Q栫^! �����R�A�;/��1͒Ǌ�0�I�d��ru�8G�J1�T/�&�����}q[����R��6m9�X];�o��ze���C�A� ( 2"��0>Z'�b��"��WD��ѵ�%
�����:��<�7:;�#�Vo.R�?�/��C��r{7�U������%���-w*9�U��:oD�mm	���a=�3� c�W�-К%�h�^�q쟕��
�S�^Q˩�R��л���>_����JJ�ITn��"p5�\[xᘶ���G�!Λ6q�wQ��>�D�;�v�:$���hIBi�}l��a�#����Mj+y��v��'Yq�2U��I����u�d��]瞤ob7� ~�����,�����'B�f�:m�4����i*S�qW�\�-�����Ȇ��&X�G��Ԙ��T����=�t+դ��<������� �����	�t�{K����"ju/�L���wX{d�t�W���=���ፌ�@������	�$e�DoQ��^KFZ�)Z��k�xpÔ|�9s+�(�$L��ܾ��U]�H�k�hf桋�f9,�?D�{q��Q��}W�)z�ޔ�7������,�L�a�׵4�2PD�)����n�
�N�$K��Z�E�[��������O>�0���
n�@����	(1\�N�)�㩫rQ��"�S
@F]�����Rb�#�\A~@0�R�LK�\(C^�����4��������	1��/��^�7,n�cF~����Gi禤�h�o޴>�թ���B�w��j�C���Xq��ZϽtʉ��#�%żx��CZ_���f_e���%u�f2�3�~�Ô��g�g��|g��<n�!��J�~d�rR�9���c���f&І-���_�� 4�;E��,�[�v0�r��~I{-��V��˄�X�2�S��+�Q `O'�g�{y�t"��̻Z]�;����S�����v%�B�ﾳH�-�z���`t��#\L���H\�PϨ!��kA5��11�}E��� �G0hQ�P�o��(]��d������?z��e����;���:[5J^E[ C��P߻�����S�i�O�\őRe#]Z�}dL鶷����
өʮ�9TW����d�\�Yk��1t��g�b�J�����"�kk���xϧaz��S¼��	i���J	�w���u�QjT̂,uDn~*raP�����1�Q�7��k�=��2f�G��Q��X|�x��л�7l\�� )O��?�p����a��l�Йl�槁�-�iO��U��J�\Cs������*G��$�DUF�{ȕ�5zkC���Q׹��)���q�Ma���.a�eL��Z+2e�o�m�y�ۯ��{���`q��(�#��i�2J����~�\���jJ�I5-	.�}3i3|�c�/'T��B�2��qO��{�Oʫ�E�ċk�Q,'u������73\5����r���5J|��?7,r��*T��M\nt�i�~M~�a)��st)B?Uȍ/�jy�j�~0X�z�������М[�VM�E'y�CF�����������D������'Z���M/������U�s�e�O]��.�r���"�e|>vX��:��*�	�1�I���L����H Ohl�\s��}|1\h�e�Gs���7_u@�pA":r���:�[P�3f8;��䱌1=��1���N��ºc�H�;�)��Y3��!�gp�R1��	U����P�$ ���7+��^e'�Z��5mh�7� �g��l���9Q�����#E����C��Ӗ���먫Kq���߮���׷Z�b�Hu��y ��Ă�R�
A/Y��,o���`�3jW󦀣��@�Q�_FE!���Oy"��etwh:)ϕ�o�bV��T[j���$���MY&R�e&�SN�.��
��<�.��P�ݙ���Y/4�̴Ğ.,aRJ�i��S����#�V�������y���[���o�\��{����/�jMY��Di��}� 3�*?ϊP�W���n6��X�7"3yۗ%OV*���u����[k�%?��R����]�']��s���:3����o��)KJ�a�Tn�P��$�5����-D�Sh�#;<ɶZ��Y��|��1(]�ߝ���T'P������ZJޯ�q�=i�ɺ����wX7�Gi��oS���*�����~d8(6z�,��(W������ooѩ���W�.w_�e��̰������8%�f��`���A���L=u �3�(��a��yq�=y�P�)j�|��.w�T�n�p
�~N\*Y�/$�*nV����������A}+8�7�+�,��2^0[�p���Β$"�Q�-z=$u^����&q��u_Z��ؓg1�'� KXe��T��ok��xHb�~�,ą$3�W�Y��s6)1�ߕ�Z�����u����?��W��Q����*\��)yXEH���T��S<F�(�=���\��w�x�8U�g�Og�o�.�j��?�=IpAn�g�i0�ɼU�E�T3��%�m�.h#�&Z��UR� P�}�R��S���o ��xSwP��G�l�,ӗ�:��P���+��[�Sz��<ּΨ�:U��E��ܮ��*��2US��R� �Ǧ��*RU#�W[��]�� r(ć�"�Y����	.���M築���6��FR�B��ݑ�>�'t40����˪�D���9B�Tb��g��P��Z�W�SkǱf�a���w��rk����"��^��8��kcٓt�����}+�s��@��w��w):iRѿ[�� t�rE���
�2&�C��t	`�Hr#)��!�iՀސ����he�I+T��xS\�Q^�~1p�79��?�	���܋�Oq�pHBdm�NwP�5�$C݄9�X���j ���$�*��	Â���Bރ��P�����צ���fS{	`�ҶV֦��w�xbJ�?w��ɇ��_[�6��E��XER���V}de?m])d�T&���{+M�FGO0㢻�>��pڝ�/����pMjX�6W���ݗ�jА�����O�ӗ��E�N��
;Ř"�!���Ȃҗ}��g�^�Bd �s����0o%,rQ')Ť'����<a�]s;w�" H�)&�"Wq2_��uKi/�@vyTfG	=�7��+~#�R�-~d��~�lڑW����B���l�k�a�h�g����x��wcF�p�¦I�K��h"8fk�p1��h����e[��aϻ$e{��.�'�|�5a)���Cbt5f��+�Lh�%��t��7��a�6Z@�.�[0Tg����z��m�������Bv�%�2Ѝ������W?�)�ѥJ��q�g1.��;#T�z�a�m�c�$��h�� R���`���-F*`�>_���EEe)�D^7^�A��n3�v�2�/G��47�������pZ����C`�l�!&5��?��d�?sS�yF�䓮��&�W҉"ɱ[�o�0r���[��Q����l��l���lw��4Xc����h-2ap��l���+�*�;ə����݅g$k�oԋ0c�&
�	��Oi��YI�{)׻�j8�`�C/��0 1��L|'Q����,)��e��nFr# ��M�x�}��`��.H)ox@b���_��!��VBͨ��۩GkU����m���<J��_�gM0O��Nݽ�����˦�K9�jF��3��=���]��K�%��S�`z �x��}����is�R�rK�E	�(��]9H�����}����륕��<�6[���i~ɚ�y+�1��ܿ6O��iց��!U��0�'G"XGg�[.���(��re����fJc�d�6�J~(��Uc0���.������ش( ���f�,�cr%��}��?K|�S�ݴ������	����V�m�����~������J��~��d�4�pqh�<�k��СV����e�w�}�;>g�Y��jp��PH�t/@�)�gog�#����I��`�!_{��ry]���̡�:&|�T�2�A�2�1����Ǆ�2��_��+CZ/���֒�)��*�䉯
����>�5�́"��zg�+R
� �fS]��9p�
W2NZ�G:�����G��rCK{؏\W!kQI�Q�F]�
���)�n�"� ����Ђ�O�8x������G����n!��QF�f�Fu�j8ͧG�{���� gŭ�\؂#)��Z�i�g�A�Q����Âxt*L�w,�Xp��U �����B�� �#��x5��a�*$s�aP��l:i�W�~�ho�N�KtM���_�IW��@���&b��"��)�$+��'�È� �g�k��=3�'j� ��i�?��0�y�U�Q�S�BR�Q&��%��,���Y}7�1�t��pjf)`���C�  <[�k`���P|�K�=+��X��s
)��9OR�޽���	l�e2�^1[��d��|�N��,e;1��8�Y)� �H��χ8BN"]T>�cr���ӝ�EO͑ /��A�S�OՌ�O���m��4��<lmХ�����;�n�]Y��,7�J 0� ����
*%2�٠�+wp��~O\����}�t�9e�v��w!�θ( ����У���R����$��T�X��Ȝ���aṓ�����u�ǃ�qrΞ;MÞ�EҘi������Ѧ���UM8bz6M�d�L�����e$��}�:�7H���D��J�|c���S�Q������h[��\e^��W��������7�B\�'���#��=������)2AR�)0/k�K�;^d��e8m��d��@o��E,�Z�u�>�]�+,��'F���?�7�����pZ��|��d1<O�o9j��v��	����]�<�%��ۈ��}���t~z�m��M$�EԼ������^�:hdLr�5��T��`�p�56o�4+�Lo]-Ƃ�����>��Jբ^����'�� %�}R]���3���+<��
VyȨd�69��;� ��E](�e���q��/�rJY�7�R�����"�K�>r[~����4���8\@��H�P��E'fF��x���
|�56i����?���c%!4,�Ddhʭ�
L��.P*}^ �Lq��:	����)�вP����;���آ�<�+�c2D҇T�Q�>j<-�=E�Z��xP�Y�ڃ6:�6F������c��H���I���g�|6wcy��H��=M�g�FE� �RT��ĄN���-/ӂ�7�}�o��5r�1�X�y���v�1���^^U��LQ���7�xW�s�x�nĕ�q�Oz�S�.�����ؠkFam�g)�<���{��A����Ow���y��sV��=4ŖJ$I����v�>���!S�o��������-D�cc�A��$�:�،����gm�mlR��㇣A��ʷ;9tq�I�c���pN�
��́ɦ&Ͳ�ӎ��Ͳ��XY\.oL��F��(�|E��$/���N��i���-��U�����i:
�U"�;{���N0a�Y���� Z6>��f������s��Z>2*�-�`��
�pE�j͔!
��d{f����T���6�߻���MN��@O�вs%B��$9Mc3i���]��;�;Z����sH��Q�������+���wyV��z����;�����@�̞��9n��+��f����i��׾}ƴ�GA�cЂ`߹/�t~YAˉ��$�+���:��R'A_�-ua�O�S���Bʨ�����b�Yš� >�xH�5\�:���n������֎�F,�u����W����Jz|b�$�A'�X$��WA�F�9#˸KU����V��=Z��ma{��R"�|	���,��K��\N�����%q+��� �=�w��z�����%ȋ�<�!���B]d9���|>|����D�1��"x��c�B�^�"W,�qKv
Ȏ1��!�Hv��	��5�4u�n��x���_�P!l0�+�|�~5?�S��X��z�v��q>8e��g���LT_�d�x�;~���U���6������yIy/}k8�3(��`Xb9s[��0eE*ˈ9���$��2����3Gl�5�����_P��*�?�xl�\�M��vK�J�*�	�4�h�p���&�Yfin�<���]o��Q���<psU[��~G��5@�?]�6]��N.�FkBX�����������`����XNH���pJ��񔳽Y)������Gh �PZ�A�����]����k�4�AA�Fv_aI��g� >��A>(���:��[/�����/.<i�C����=�[NS.6�B� @�.�M��^�v+N�U\�[%�Q-R�#K5���`�U?&��Fv&�2I_r�Lrs>�n5���y�֏�:�kƞ��n���M+��ܟ�ip�E��]��6C� O(׀_�y8v��xV
=~8 3V��2F�Y)� �|@��"�l�w��n�&�홴������~��(~�3��e���g�����G��#�T!�Z}�#��~y3�T���b�[,hU��˺n������@�Xbw,�B�1�>f�����$9��B
��2ݹ�N���ۂ�s�X� �4�o�U_6��b�T�
���	��O�����5����=��'cN��i6J�y~b ���{�7�����ߣ�	���:9?W�|p��%$��_��0N]
�65`V��� �+>$F�Z/	�D��ҩ{��Q��bb$V$U�ʷ��)�$#F�p%ߜ"{&��T5���k�D��$_�U �%YYp�l�ೇֲ���5ĺ�\���F�1Y_eH/ԏ"��1��^>[��Hjc�_�w�eb�r�U���|[�M	_���9�H��n��ly뎀�o�| �M
�� ��{�sOu��w�!銣��AL��<�y�����k�+]���o�ƣ޺7�M�����Mi�@�a�T.cS�xѺ|_�݃�M���7]0�9����0;���I!D0���l�����r�����A�YLO2j���0��Rw4?3E�A`7tȠ%m_ƯP1,��y)gµݺ�����.�t����T�����fМ���/]d��ɝ$��F������2
b�W��#��x�D����A���0eW��ie�]cj�b��J�U?H�=Q�($��$�r��a�"���3b�d#(�u�{�{7)zǦ=�6Ļ�EV���.����h�=�w�u�9�_���?<�"p�\Ȑ����uB���������:M#ڟ+'��c�jµ�
5*��"$�w�c��^7W�j�]�j�ʻO�����cL�璒�y�@��(��6�11w�_"��ҼK������7�uo4��|�WZ��\P0Ryԗ��^���X���4��U�dFL��z���ٛ�b&x�^��4D3� ��݉
҄L�)qu�0)�K�X�P�ZSt\��^Hk�d��>B�����i�G�8PeG�����9���D���m��yX��8Ahlu#J�-��Ew��Z�=�B��\-��#sAF|��� ��3�D�Y�֋>�������7��r���=k�˞.E<������;��8����'o���&ϕO������T�P�.+]ּS��ߣ�6�pe\�j����̣��%�U�5 ч���cY!|i
tr"��B �P���mow�����Cf��)Ehp��J��������o:G�X�5%�m�+�2O�f_�����GT�J���?$j)��0+�ͩQ��)#�'���\8=��j*1�;���H#��Ӈ���I�&���:�x��A�}	�N�r�ni���RC9�����t�ǧ}��{+�.�(M����s ��&[�!�+6�k]�������/}kD�qAْ�Z�������Ʈ����g���eK�v��J�vU���H�*P����ͥ��Ao;�h�ȥ�p�{F�����!� k�_���9�h�u�\2d"A��F���r+���E|�����ow�I#�|�?�,2��	:Gb.�܃csYH�j�kU��4���Y�[Γ����l���@�SC�Y�*8�Y�v��{���b��?g
�5��U�`�];x�רo������],}c�{���}�'{bB���(�6��p�q&���O�S�䚝&��q%�z䓤��[�9�XX������D@y{!�2�ܯJ`��,���N8h���v���\y��@n���3���kx�pD���8�	s���DZ��o&ׇ��0KI��b����f(������lt�S����2�+]~I���6{��[ˠ��O��,3�h	b&jrR�*�U>n����^�.*� �,\�YG\��?�L�ί����)��<ڦ�J��\�� �)r�pR�T�vn[�g�����+N�Zᇨ}i�SBt��ei-$e&�lu�g���@W.����݌��\�eo���I&�]�˜gk�]`X�m#�d5�l�dwH/�qz�-(˴Фa�2��*����彔��/ ��;'��^��^��^�>��.][�BU�J+A=g�)W� �ֶ[`#r�W�SF��@��ʦ׻Sč�)of�9^*|D�[!��Š��o�lX���P�"H����[�#��e���,Mb��6�]���l-;�2�i6k��y �p� �f�!VM���F@�rS�Ak���-��/��0r�����.�&_xa��;�`}��*%Ȕ����^�r��"�i���R��.�C�U�}``F��[5*[�f�����΃�#5xJrB-D�q�G+`"\r���8AbV�$����$�#���֟%b�$��G"��7u&��,��D�):��껿���x�M����� 6��.��.ZŖ��?@ߋyFZ
v�6����i��� �o��o�2�ہSgN���_�����
:�Ǯ���ߕ�=b�[/��J������C~Nl^m���,���%�}�,q�z~#о5p!-��/^J8/�%�m��@�,اw�%�&�XS1S3�VW�z�X�c���@;o��O�B+����fNY�N�3bX�i���Or�B*`�w�U���Nz#�f;��݈�BD^�˦;S���p��8����k(���ɔl2>���4��8
u��|��e��펶m��:� ��҄�	�`<�Ot�o����/@��'�^�l?VM�X0���P5��j}�dK~���7]v�gQUݭ3�$�Q�uh���ɹ�OA8HA��*�B���o���_��$cX��L�����bT>s�v-�~ݿM����t�|���I2�}��,�__W?ɽYU�^Z6=�")�Z@�:�X�E1�J���Sw�B�0I"O��@
'pj��J�Z��җ�'��mY���Qc�aJ���8�(/�~�Ȟ��s���R�\�5����O��7�fEΐk�2=Y��F�?%�MI���P1i�;t|}Ⴞ�7��A�8���
��r}рn�e�P�w3�&��W���� ��,��<��|�ƈT눛�����×0��Z(�����Lƭ#"&���O ��U�4�X���eɔP�O�U*�<��퟼��r������*�qD&��ߎ�*%������W�����k�>��Qǂ���!���]�HwO6S�{�a��~}���Y�q���I��q��&��gȱߐ�r>�0��5uv��H;��$����64Yz��r��
r��}Ҫ��������wȆ�:�j�WF���!�:W����#��J"�&D&˰1���ķ_��V��W����(��)�77�!��--�5�a�?��Dv��z�Of^��]o�Kv�S�a��ZcK��sq��{��c�G	)�%�olg.q'M1k]�su����=v�~ʵ:o�`�UkU���	�r��/W�e�C���a�85-�$�J��ge=�&9I�xJ{�Z���.��On�����<^�:���O0)�q�P��}�������9��U�=��0]0��>:��k����B� Q:TS�f0U[<���ж0��� � "�ŭy3[x|�uX�2���б�C
������~��D16��ʜ����u�x�6�-Mռ�.:��D�<���_���+X\JO܁~}E�!s��]=j���8�|��T����q�"���l���A>>�{7�~8�Źvl �_U��뜹E�`M�! ౯�]
�L:(�ºB���](���\{��K�Z�P=�TV�Y/O��$%��)bg���BL��8���+���N�D��WA�HË�0��� �l
�����z�gr�O�G�%˕�=�`,@*�q�F֚]	��S�lt��؟g������M�br�C��*��W﩮��RS͂��;K<�{Q�D[��9����x���0Pp[E�'K���@���;��X2Q��1�>o��&����h��nzi>&�{s�P.	^-?G�A�e�)���6���W _�9;�� �}�ʑ���k�"Y�/��{|hg����P��9�Q��̉���Q����S��!'��W�����'Ar���t�Џ9��X����*h%����ע�������"��?�c��ڢzc'�QIe�C(��H��xQ�J˥rLb�=��'#[�U�{yn��ɇ�pN�#@\�?��yS�^lf�� �	ޝ�N��?βK��I�A�r����L,��l����$f�8�4��~����/��� �Չ��Nkp��s�/0��E�0�1��,�C1����$+����_xh��l�g5���B1~FP�ԨDu&)ɕC�M���̠��F=1H~��o9!y�)(L�x�������w�Q��W�m�s�t�&��h���2xB)�ة�v�"����XǍ�mt��<a0>�\2:K 	;?|��L����������p�T𹎖|��C�q�y#�k0�Ѱֶ��y:�:�$�;D�%�`r^K�J��m�V��
�F��,�=o^�}Ly�sЃ�>~�sט7����A�X�[d\3�"+#�ɹ�@�g8�
5�⽶`*I-�6?��C{�I�WE[��T6K|�1����[��,��WL���Ut<Q�uO�N�5��W��w���|W� ��m��/���[:`n7�Y�^�t֏�5=���(Cf�Z#�l_/�@�4�P<XR�(*[��u��̙�t+����f�LQ����=k��p��Pk��'N���B'�cO@�Zy��+� �O���F�>9�i8�G��([K�Ix�hoDq�}����w'5��Z�H���i��1��P���d�����	ܜr��T�\��x��_�E��E�+8KV3�g�\Ь���@4�b8�����*�W�֟+%��
�ޱ���s�v/��P�_tp�R6��1�#��'��r�Q.����a4���/w��.n�$],�^x��a�ؿ��67���J�25��W��_�����%�H�7�y����z���=[��}���M�&q{��Mm4�*2�&��s!�*K<��AO��a�Mll��w��-!#�%CQ>��$p�ME#ؠ,S�]� �gjG�0�@|'��y�r��D��P�!鲆w%��>���5�2�D1]Y[Ts��er��������_	�u�K"�x��n"��q�M9 �	�翖��w��&�	��z�t�����R:?���K�Y���C��F?u��YnnG�*�J�yb��D�s�����@��-�Mاa�[�!����96Pg����g��f�p��6�_!5¢�l��qb@��Ei�/sg���T�����6�L9�"0
��@ɔU�̄X��$�@o��6\w��uQ+����p�<�k�-10��	��^�U�Qg��,�:����S�
�iuC��+g`�4�����I�z*�����w]�Q�`��u��V��M�u��3������esP�C�E
���,��b0=k���-
�ig�e�_�yLO�f���4�|q�<y�(�x>{�3m���L�Q�lI�/U�s�`��F���aB�����Ʈ��a�6��If��J�lUّ�9I����C#W���]]-��>`%��=�g�v>@���������ȶ���G040t��$�ܤ7Q"�V~���s�t�ЩA�,~J8Pa�+���ؐ.���i�y��#HeaXZ�Z0X�GD���`6�)[h�����w<���u�
���F�9�ub���H�"�* ��K}os�X��bB�gꋅ�e:1������չU���LU������3F�&D�������6�Y��_w4 ���N�A��2;/jxdB��P�&��ܙ�%=�<�zt��s�^ �Z�у�q��h��1�������uJ��j3��y&�K]*��}F�� �jӳ�H%k�7���KJ�R�M�SVa:_'�l������Dp�z2Q@ZN�=ic�g�g�
���HD[��fQ=��#��z%]$�X����d�1���xd�eu7�ry��5���X6�oĕr���&hxVɻ�8�)a��S��)3�w�q��#��6�����!w�����3(��K��"��H��W�S~�~l);�%#��d��G�"n���b�Z�	�Jt�L�A%�@� [�������ۺS�$�r�̄�6�.�d��$C��D�9�*$�n��X��O�vtԤec�������6�o�����3��k� 
}zg�N�/~������n'�N����)�1;��)�+4)�$��և���U�6��)���/�&�[7ef�1��U#C
U��8䫖����ٶ|;��\��}<���Սdi�ׯn��	�X}���CcXG��4�i� ��_���&y��z�a�X�u�i��{R}Ƭ���I���7{ʀ|��"*�ouu�i�����ݢ���4$(�ղ��C�
��M�aB:f���*���v��c���2��5��U�@����9�(v��ح��I���I*:�V8oH�/�h'��0����윂���1A�sW4�W4_$尴^dr+����;zb��i�Swg�Myw8��x�a�Ӧ��6�ݑ��s\3�n(�.��LߙRl��\�ÞYt��-��@�
�j�'������ �Z���d?C4	E�A�I�������)�Oj��f(@�
�`K�(�����7p�0�o;�� ц�R8~�:z��� 3^3���G���\J1��������i�`ߧ_�n��(��<N���f��bz�%�$T\q�����N�`����� �R5���b*8C��'�RH6q�'�� �"e�]��|qUѰ.�Gg�uxZ���6�<S	C!Hi���2�'�M�Η�C�⣌��x>�Zh��Q ���o!u^a<?��}L9�?���QVh�Wl��A�,�ň�4���?�{̠��65�/}� ܐ��7qux�MG ��Ti&��R����)wէ\���Hw�M��8����2k�g�6��@��fP�;��&�TUs�ڶ�r/��i�`�P`��BOI�zh�u8�x(��ė���]7���Ve3<@�����B(�������?��<Q��$��a�vq"�I�&�3����ĠhH�op1(j��^e��mu9��9]���5���yc)<�-��/���)
��`���i��z��~��V�~57��]�u0��;���X?�Z�eW�B�ұ�P��F֝�B�jw�3H��=��+�b�M�;V��0�j��a�d�i�V��W��+p��2d
.�kb弳Z��S��*h�' �ɜόF�s�#�}�/W^n�.-=�Ūi�Mw\"bs�>�30O��V�&'�=3�#T{;y<��8����uc@ �o97��� k�\�DRa0�\}7�z8Q�,�b&�ҝ���d�^�o��x�C�0J)�0�|�Nd�7+���j�A�zQ.�Gsc�Kb�	"3f��Q�J^:�Ɖ��Q_>���$H�V��~�{���u��c�@��ХM��cЉ�}���n��2mL��cӭ���^&~��)�X@��j�]ЄL6ȹK��{��b��0s��KpC�7���%�hR��}
f�g��o0�feu4�˿R������T��YG3$�)��+����l_�Û�d�����%����h����	bg�`gr-�8N�H�^�X�,Y���k�6 t��q�}z��� l$��
Os��
�5�{��UNo�H���J.	�])h�0��I}?��֠ �1$�}*2ƥmr�!a3�A��ֻ%��~���#��.�o��I�$����U��"��l�����[?�͹P�ZAp���[���{o��%+P�3���1�.��K��_���T)�y%]T|��E[���?�6�I�Sɂԃ	Wɟ;N��&�x���\:��K�T���S�r�1�,ĝ�)*3/�o�Dvίf��(�]��±���ErJ��z��\Q�$�w�������*���{�Ln�]7�,��8^N��-,�{���X�m���|^#��H����x�ï;�yKA����oΑ��+�KD!�?�*�̇qlé/XH-_♗��o�=<�}zO�4@TЦ�u592�!�����6�D�4JZ��VNkQ(��|��x�{ P�$:�̪�\���+|�{�������Y}�a���d���e.(�d���J�j������[N��A��k�az@qq���N���/>5������x ��j�����T�y�x�.�`����&�4�{��Q`�����j�N��/`���MD3Rp:���w���� �du�����$��*:X.x1�#��t�̝�2jl%y���7��yH�,�ʼ����"�=	�9S 8�uҦ���ꚬ#yR�Pi�"����QPJ��ROu������0�C�N��x��~rd;���y+�^I%�I3��K�S���������}�rF�z �q��)��Aɐ(wg3�߅�+��!6�%�ޞ.����}ׂG<�0�W[Φ ��4ǱZb����]8h3"7����۸{�_���M��&?i@ 8���D�or��� ��2\[H;�j]Z�G&����Të�pl��2��&���K�ӆmM��4�4���F`Z�=-U����x�$%�� ^�ž�caSm��|�"7$*k��/���]���т�Yg���J���W��F��0���_]3Z_*����G���T����IM0�#��D�����t�#��I"���۝��6����%[�k����;Mk���pҶ�p.�=��^U�D�Vj6T�Qʆ�� X\�ډ����)�����z��&���H���C�Y����h��!��܃dSPW�!�Ո�NHeES��*�L�CE-p�x��RJ�)�E�dDr�0�	�{[#��t�T��5~nυ�Ho��@�S�d��w�+mu;gzq;�^D�E��".��d�ؼЋ����`n�ģ��(�v��m�4d�%�Y[�%}G�z4�ځ�$8v4'��VhUwâY���P%���1Zm-|�o�5�я�#Ծ�2�,n�Չ\nv���J]Z �`��e%R�+%�h�G-��Z<��p��P�0%�m���?3�����YQ�(�p=�ƓU}�{����],%�E�lJ�oF��,ޘ;�����#�߮S?�����ґN/���]���rSu��-�%�zX�Jx|���{x��yC�
C����PT^��ҭ�|������v�H���^ȹz����}�z4F�v��1~ u*�HQ"/l����N�iϫ�ͺyo*ת0S�Z���N8��!���Z$kpAXY���)���T���I9�8KB뙾4J���h����l_�D�Ei�%�^�!Pσ�f�Q{�|�]x�J�����_�}W�b�Q��7ʹ]��\����Li��`bQ�����(d\�y��H�0�p�&�E7�Y�����C\� sC����P4��V�]"q ,�c�N�̤@]J(g�ӢЁ�̡ �r�o��^ٚ�2��m�ޞ��&p�r��V�ћ�DN�p�#�''�I��,D�x޲4F(���$b���V�ڦ�5r ��U�z�"?�#�F�r�N�3�1:�s#N1�s
D!X�A�hHU,��O�*��C�8<�9���8��1�pՇ�x'z�Ebwo���j�e�X����s$�� m�V�%�B� m�d&"��y=q�y���7?�&���!@4�~�WFhm���Rﶲ}�+�AM��gb���6��72��ign��(��P�͵iS��kML�'�����ƌN_A������_Tu���nq����+/�ne��)׺p��v�\Ȳ	���6a�d��b֥1
��^�ج��'jU_��ym��)�3��h�����D�(���F��Gl�C���H�^9�l]͘������U��?V���R�a%>����1�cO�|�jo +�=��ro�\'%u<h�ڗ��hL%TWG���ґ"�L�w�|�J�L=\ݣ��Í��x�ק���^���U���X�Tx14��Q"��f�����h'�>yÉ�9+�Hg�������G���c��X��Q�/�2T˴Z������xt"Z�R�}�+j��A�Ws�
YX����t�;�W�1�1�HGH��Do}�_�M�Vn؏P�i�;���QΈ���,-�ͫdٜ�����#��_��a���*�ĒE�7i	�٩ƍ+�y�?	�v�ہ���:'u�B�-�pp@'��w᠏ ��Ƞ7Ԍ6S�g��7�����!{���Zs������V�����/��hv��c(���x�G��;	-�j���`�8�8]?w��=�#�Oȩ�Η��I�tA�y.��E����s^�9��	�[i߱J�S5&������'Su�?S��
+��v ��A�^��܁c7�1���9 �����d�84�Î��m6��H�&��G\Wjϯ����k�
}�;�r����9,-]��f����#��j��5���S�|�<�O��ա;W��qJ^+�?a����^�Y`�XK�r�c'�~w��Jk�\�s˝�����;mZ�YDŀf�4"?�!Kj���)��Y#u׺���|�Yo��BhO�6ۣb�F��.,MH��"I�r�|��&Hw�t�.M=CKk�����9s�ˉL�Cl�u#f�듄-�+N�O�!m��It�@2[�@��g�+['�����:�'��7^���l@<�'����qOŃ�"nDV�*�䖨Gc� ����-�h,C�M8&zt
�Oa{�T� E�7XG��]e���w2H����" wB�6(H9P`}H��R�~(�G^�����b���0�Xk����i�����ʱ���ʅe�ɩB��,/0h���)���(�x��������=%��V#?��+4��8hL!�{�0Sl��?c4d�\
��u&՘4.��ҳұU�|z�#������IN�Q�@̡>���0�@�I�?�#S��I�`����K+6�#G#\�*o=�d�Û���==��O�� ��/ǼЧ`�Mo@<�_��@qns�	��u�Z�-���x&�`�NH!�yj�U���T�;/Uf�XP�wi�8P�:�쨘�6�"�L�����4��[�6���Bϓm滊�j�g!�(me1͵�<U�at�_����z��K OS�+�WM��g�s��F�>��'*7t�5d�OVߢ�RT$�X���Z@_*K�m�`�e��It��p�p~����u؝S^-)�m��R������w~׈N�џ2���<��Ij���v���g�K
�@7<��gΣ��g�%d�*&�W�����W`��������ɇǴ���Bgo�sX����[s�)�&�d[����Z�?$H������	����j#'�����;E[警���%ʔ`�݁�ŷ�r&&�=&8��?��7z�D�żW�7D�`r��v�r�i.��DO��w��.z����V�N1��ڦ�d��\e3�8�C�"*�*���n��6�v�s��#�ði�ᣦ(�ebC�������[���S��e�b��7A�����V�Uh�m���8~��PT��f�����r�\wt郋�^�/�R/_C3��/:�
�\JA{�:5̧zK<"�����Hw��w�-X���}�bQ����hݧ���m"6�l]��O1�s
1@�UwP3�W>5�����0�+ϕ�t��5.��NC�(���Q�9�ǰy�w���{_��ܤ�0XA��	�]�ܼa�Ⱦ�1?�\�xk�WIq��'��m�#^�Q+�fk�D��4=лr��7�lv��t��d]�R�k�6�(�_i��\��E{�#��]̖[5/���af���������	A�1$G�G�P`ֈ�Z�x��X��C�(F�"��Fh�5�u	���y�C�C��_�\����ʤ��p�j��96Ȗ����X�W���oue�v^x��e�����A��8�Q�yB����}z�)���z���.I�d5%ͪ�,�PC��ܸ��xbIf�KC��Јɗ�o�6oZ�����ԕ
 b'P��8=8e8��H�۔H�����s21�� p��詀�g*�Al�&��_����.��~���1���Ǎ��B�l�po�3Z�R��q���Y�Y�Z$���{t����⟜p$l~@8�����W��,��i���S�ـ&�A��	!��P}.G`�E�y��⪾��x\z��yK�L��$UQiV� ^9*؛���{�Tl�<}4G���d\ۋR}Uc�׆g�R�(%l��D��/p���]qtk �)���v�l�35s]s���o�?2��t���� �q4`)�
�Nt�0��ݳXT;��2�ZEK��n£�e��� �|E\0yЪ��rd�w���)��U�KI����B'?�/}��aV��[�1YW<����ⱲB��\/�1."�!�g�[W��RGƲC��`pu�s�_�M� @�9_�����=nFY�$�W��H~f5��g��˖�7"� ��I1��U�v*i-%`��5JM%;��g��7I���Ô�O=R@�L���� �Eо�-σ�)e`�NQ?��h{��| ǩ��o��^й�;=�X>�WFIv�iᔃ`4�Y�N#�Bzp�����4st�l>$�!I�Zp��~�����Vz�P�;�axDl7U}��i��m]�u@���n[ ������:G��^����03�لe�汥�SY�q���dY�j�­����Q�[V����*&c@�RVðGϸ-8�-�jY�������Rd�Rv���	�t�ޭ�#Cra�~�{@}���)��[#���L�RJC���q���6Y]|��P�	���u�a(dG7�}{�	$c�@��z7�����K��1D���������	���W���Z�.Q����E� t���&_*��D����鱊�¶����qt3�є�F����������5�]2[?���<�	%��Uf�ҡQ�|���ľXo;��⍕�h��#��{�t^n��A�i��!��a����������<�<`)�~ԝ��(��b��U�t����n���N:9��w���}��3�WCd�'~���uT���'����xR�<*j|����D̻��̶F�C���N�6F�p4˥x֫��@���]��,�wv�zA7�HS�dM���T�������prg6��
�V��*G;}���yΏob#@�O�UI�C����4��?�e�X �H�,&g�4s�w`m/"���Z�x�H�2I|�.������ۢs	~���S�ŻY���������n��ۿ�Y�-R��'�T|~���Uŧְ���6W�F�16�J4�X�7���3Vg�@�v|�lppS��)4>� M)[x���*�Q��NG������>e��XuI�2���g�w���LkN8n>#��/���ʒp���3��ؘ�����CP�|(�}�L���(3���aO���)j)�35'ZCW�
��5��.P���eݮ����wUy�ؔ��֬�:�k|�{�l.����х��:(�o�J\�#�"���ESz�yA�6���',���w����~c�_;~@�"gEpv]\5���˸��"v������O�5{_F��;D:�gW��m�;���3=�~Q��o�����׵ƽ\8�������2���d$�p^'%��U[p�Q�ӏ#%�͓� �n�R����*�/�-k����#��e�֥(K���{K�^��yOǱە5�l2����ɹ/<}Dr�S\t�S�%Noj���8�z����� ��o0|v[�
��������v�!Ӝ�TAʎ~x(B-�ѵ���(fy�n¯\�� X�����@���_�L��ݶ`k���_"�<���R3��%��Z9���D��ȹ#�>r>�\��ԅ��8��&����C�~h�
a�M�UN��(<��t�Ɂx�B�'I]�g����qW�� ��j�ٙ#���y�ۨ�*KȘ�������Ɍ���H�qm�������MY��K�ʉ�k����E��2& W�>	C�j�K��(��Q`.4�\�+�C��k�"�"�Nkf��w��Q���u�x���p{���̛��KlD�Q����a��P3H�ȉ�L�}��g%[�ۤHi�N�s>�2g���g�@2�Ϡ
z��?(���E�w��͢I]Gc��~�sOQr �v����z-V�R[��C
���qy��I=��KB�U�����?�����=$��~�d�M%�=��4t�gk$U��
���-Wݴ0��P͑vJ�@���t�2�B�j��lSs��N��7b��`	��d7V�sAU��M���As��&C͙ �����������%��;<��譹U�������Ey������ߗj%B�J�Eg�I���Y$fE��JZ����1@��&v��ETsdr�����)���Z�Ԙ`�4���g3�}6�7R�_L�����7Z)d�P�z�8�2��%��b��29Jg�����ty���V(�L�>z_��ֿ���=)p��wg�Y� �l�*?�Y����<Zg@��d.�r X�|�V
��Sδ�u�_��r��CMڕ"`� 8_�u$�gw���um4y�
����c�C3�3�[NW�b��=]����4L[,s��~��k�5,��~�}��p�'S5v҆b[��v�K����������KYq�d:��^�#�9��5�*��ǹ/;��*]��l�B:)p��D<���k�'^7�7PG�ߗ�"����:�@'^�( ���)L��1��$��`�\N|�	�%� jE�`lD?�N�F`�}��B�L�g�$As��P�2��^�i<+��Ҧa��#�P���Fй��/��H-=��lr4����*`k��O����B�I��3;�E^9�`�9����X.sQE���G��V��L���b>)��"Ք�Bb��]��Ad�&���m�l�0!�t�l����Ă�)�����2��MZGx��B~-A��-{�0;�3����G� ��C���"C�F�\�i�v~��4va�G��6q囓L���u�L�L�tR�ꛘzqՆ(F�=���?��ɑ��O����F����8 �-�7��]�����+?�\�.@�N�7���j�3SA��F�K����4�=����g)V�F+��L/aW�=;��h[(_d�d,�D��g�ŅTmq���`��L��B��G�a4���6�|ږ�JЂ�R��)ng]�_��`�D���ߝ�S��ReШ`$4�ļ��Q�iu�����X��6"�^�ZWVj$v�+�)!(�rK��Q8~i}�������d~��V;P��[�����iW�#�N�tv
���~�e�{�H�_�eM��P3e?]	��ɱ (��H���D*�����߇9�����A�$߅=��=�����C9 �I�E= �δ��vqg�`r�O�ޣR��}؍;w���;06��O����[g�6SE�rE�}-g��=�P���4�qt�9��)8���1���L�{6�G�)"σ͞` A��b9p�3g����\�\-�����Ӿ���)ex�������޺��wt%r��5D;����h��M ��d��
�����ax������-ŵt����B�C4�W�n��*� �R��D!���k1� �U6��}�r�yQ�xK�L`�U��_M����a�y2i�0�b���`��K���Ӻ�PVC�\e@pk'&�Z��5��(@�^� ��g��-C�&~�*�����1����R��:LMۢ�������3v�����`�E`Y��qV�����l�Wz.b$t�~�M�����Z��~1_4Xk���+I5�b���eR�8����-4W�7�����?�1�;(�
_"����#*�~���_�/��;P ����Q������o���[%�������b�w�$S�͌�_����m~	a����p�j�@ꦪlv��8���=�݂�6�cCU��B�A�������@FA����HT�{E���R7)�=��Ւ@���k�����В��g� Dg=�*�Od��vG9
/�3�7�ɵEn= T}����K�n	ea�Q�,~�_ �W�#�"2y�V�%���*� %U�9��$��j60����>��D�8n�E_`��)�Ґ�t@"�#o��	QD�p�Wsp�'�ޑ�q���Sߪ�xD�Mg��&'��<��~�iN{�� ���9,��g��(c9u:�ʧm-�(��:����
�CI1��j���?z�W8K��+�9/F]��a �'��
ކRZw4����IIؕ�xȑ!�����4rj[?�k�s�?�ηbp[�1�
��_=�^Z]s.P,�<m1�hZ2炞.�%���T� �&Q�_v8Y�ސ��-�� ����-��Ku�πd����!1'c������o���D(��'��L6-�;�����fX��L������" p��(�"{�ݏ`\�/5�
�j��V�p���m�=�h#�R�ssX�V'T�?�~K��d$1�����:C^ 5Be7H�k��L��w����-��)�7OL��5_����0�W%�=��e��K�i�������(a�u��.={��d�VS������#��?�LX0�}bcnſq%��3pX)m�����#bP6�pP���8��Ȑ���X? M\�?�?��	�6�7�xF?��+�;5����3����
�%�4�
��D�uZ,h�۬CT�D��g�h���t�3��n<�Aؔ=~�a, �9�7���|�P]���ax��=��oa�a԰��Q��L��:[eW� �+�VR��%+Oր����?��`N��_��ݸu7*AD��΂�:���N b{��ME��n~�T�ƫ�W����|�B��Y�����29Iy #��^VKW�T9rH�@,��֩�����
�sG��=
=<ܔ_�Q�
�5*6�@Ԋ�K�%�җ��>"�_��G���s�1��4�n���n	�Х�|�37����:
�;�ۙT����H�s���Ů�,�7�5%�i���.v)����U��iE�,�Ŷ'�8�m=5�Kc�j�C���ʗc�X5׻t������4���\J ���ڈ��0w�b�gk�x�_�b������DB�%[�Zs�꺚0{f��Y@�h:3�]�$�W�����p�P��W������w��2	�q�Rr	��)�:�F%�T%�J���U��`A%���C
�P�rX�e�з=��<�U����{,(~f�I�F�Vs�᧌��H��=��F=��Rv
�6���ڸ��<k8��>�ݸ�D��?mY:*�f�I���9lw�&����y�\��w�y4@r����(�� �-a[�,�k����&��˷��:�u�i8�8�jZ�Y=:�Ť/�m,o��}�7��P��mMn������w��$4&��p�ĸ�b\��KF�Y�7��Ǡ36�^{}|����ύi�y�\O������r����r[��o§ɊOh�P$���!���G����^�lɩeaZ�*;��
��t��&vBb�׻"�_8^�UV���Q�IY�c��Bb����g�1"��4��{ެ��Ǌ�jT��������7DL�JuÍ��'AB\�'�o3�q� ����boz	XÜ.}�¨���ig@�<FS ����nM�T�)̖.o��=t�mDI����JK��,f���9�r7<�u J�Ʃ�8�������j���_�+$X~N��P�3>�� s+T~�h1�����R�w#��#����iP�*�Y��q"x\y�*��
1>�?����=|���PA�Hz_`������X��P���>�:I������cQ��Y���u5�D���5Q�`o�6�'���n"��~�����!���al��6����~�B���~��L�P��s˾#)R'�ξʟ �*��k�7=���;{��fQ�[��BO0N4��>�5�UAI�- il��,��V�T�h��f�Bي2
M�[E3���u��"�(��݉�5��k=�f�	V+���g���"��G�����n���1D}��s֖��l5��|��蛈�9�����[o~ k���d�@}�\:H�AwǪ>5��]^5�o�0�Kf�n�c>��bE�Vf�a8�l�:A1l��/�j������*��G�/$��-��N�������GW�w�^{�B��E��Jiar�;�{�vt���8����q~X/���V@� �x��1D�;x�3~���ư
�ث���O4Ÿ;�ɴ���8��Qsou�x�Z��kx7�v�(_%�_�*���`����Ea@���P��cV�z����#ޞM�M��w�"q��=��%'����A<���-��߯=���f#5CV�,J8��^	������肕(�|@zrK��g�D��D��=��2T�M��?�������<��Ƥ�9���}�q �k��	�-,>$�i�/��� �
�$���?q\,K��׏}�ik��!�,#�#�p���Rl2��k��c�{`]|�L���\��"E9�)��أ<u`!Y�8�4�s5l��$W��������x��Qu�ò	G��}v�*IZ�O6O�P6��O0���ܰb�d6��׹C�(���;O�A�Aܶ�q�n���_�6���k�Rd�D��V)�p
��7�����ًM��v��dI��,̺�(,���SP�&_�R�:��#;�{�Y�%9Y��
%c�cXlVM@�,�e�`�/J�$s<{�*;��7�5�rs;9�R�˻������ �M�Y��mV���QN���JG�ܝ��vG��$T�P��,L��!�N�I���>%Y
h܀Q*��rc0/u���@�wd��'7��qc 󉘉���l���H1���n�r�e(7`��dz�G*��v�7��_��^E�L�hR���c�"l�(w3Q�k];b��Jrڃ[�Q�L-������rh�gyW�g�,ʤ�$��&��\����7�寸^�DA���ۻsՋ5'P��b�!�,HI��a�PS�> $�6��!b�ף�7 %�/�	4��-/�}f~�&���w�CՎ,��A �0� �|䶩��bN�	�쓴�w��k5�N?���8�z�5n��g����{2��t�[P�Hp^�<��j�� Jh/M�/�U[�eo�PQs��b�E93hq��~CPe���$�����d|H��rl�xL"��o^�4�Y2:�\9����������W���t	{�[G|�S��)K��bf���e�͆b�	�f��������h̵�HcF�sr9��o�w���x�L��6�W8F���mh�V�!ؓ#4�Z~���j���Ya���ۭ)�F��?�7�Bh���"��_$>��N��A��r�ġu�\��,��Gb���n�X�US���)�W�֋���	��ؠ8*��3�?�]�<�s��1�5+1iv(5�:rO��=փwM �{H��1}	��7��az�o�e�M�����V���J ��Ɋ@Y�ª�dF��6����DR��*Es_Õ�X�@u7���K>���85��i�ůC�Ү�ߍ�$�Z��~����
q�s>����틨�9�:�dU���+tA�����}I��ׂl�b�{[���=��k/D��u��I��m�����%�%ؒ�]K|���g4e��Ƃڃ�ԝu���|���3ib���SCۮ�΀��i}������_�ؐ��qFz��3gZ7y8�X���y(�z�����<�|2cQ�9�u�|E��S���V� �:���@։Ν4���ԥA���̕�<ŏ���G�֝�gu��2�Z���jv�	�!�Y#���_�#�k7��|G:< 9��]�����'*y��nAiV5���7����-���f���zO�,�2g@v+����2I�[h	�z�@%dt�Oڈ�U}����
��n��4��Y:[h���{�G ����mD�*���J�/��� yL�U$Eh�%k�N��|��>����ƾfa���#E�k��%�J[��N�-G^�]c�Ȱ(��M�*�U��rdG�\?Ի�}��9L5��p�j�a�}#PӚ����FI ²'vɕV"�D__�K�F+��0:rDWA~
��g8�@5����a�3�G.��1,p��1�FUh�.��޾]JB�ӣ>�K%u���� X�W2�lP�s�w����W9En�~}��4��sT�X�F֟���Ř��� +�Su�ӛ��;�F�˒�z�86� _�v��Մ AWv
��"�,;����K�x�'��EX�M����Qp!�{�s���mN Oܸ���e$W�C�|g_7���pR%�;C�A=�r��bu�V�}�t�P#f��Z��:;J�ϵ�D����(��ډR��AO�ۃr_K���̼�8^DXɹF!2c	��A$��Z��Aκe��8��74>i�6�@Y�'���tB�}.BH�k~��	�V4���eH�1P���a~�qd��_��wJ]"����6ƅ2}@�%X^�0c��߯�EY�ڼ���~��K�z<@����B�t�ۂ���y�<z�Ā8����Ar���g��)�~���@ֿv":�#(C
�F�/n6�:����~w�u�~~�ӳ�~�U�r�#j�o��6!4ChJ~�8.�z�Cp��$�eiل�7�ɑZ��� j���0F\�������a��\`�7#0ښX�&��A�V��7��I�N�	��ckp��MR��h'�7,�]d�����R�G�Xw_���y1�Hv�N�ʉ���Jy���_&M��N�+���4��oP4%��;�#�Y��&���޹�'��xIWV��;�r�٢�R��{�	�g�O�[p�n���9��z�*�ȯ�����&ZV�:>prr����g�6�M`XW��H+='Nt����l�48u#����@�Ne`��ų�#q���E�~�������M*s�4�>ʤ��*r�P�(BKO�Z��)���PEз��Z���)�#5b�2"����8����f(�۠��d��d�I<`�<���bt�66�ꟛU����d�˥l?�+�������2��-J��,���"7v�����9b�V��ٹ#"te��'��r�=� ��\���J���:�-�:����?a*vT���ek"�-��	Uش4k�@�uL�K���ie�z3br�dN_��eK��=�\��3κ�m��_-�^��h�%�3tte�|0�%8����7�^��[��8<{7����7�M��mZ��/�4���m��&�{)�@	ʤ�ѡ��K0#X�Q��"s{��Y�7U�L��S�9�B�v�?�*�G ��07�Z5�n�rF~�d�Y�N�(	���]�kͨ#ԏ��F��ȅ�5b"/w1ȿ'��-譠U���������O(�Z~�Jϰ�\R��
��O���q2�#�!?"��^o[Z ��9�sM�R?J6���v�X�
QP�˓aR���^t���B� �U�p�qPbwz�+��;V�T��?�:(FX�b3�t��Y��>��RWᭁ%���?������.� ��N���J��W�:�������%�ش"��˖!Tք�YPڛ�ԟeVHAsd!�wHfh &�K��z&�I���h�։I�,*mO]\�eY�"���E�xHnLX��sg26*���ܭ��'wȤ0���:p	�b�.����z	{�pd����)w��ڳT_�Ĝ���b���ם�t�]�e�̅�����;� T�=<�����Γ��%�"^��֎)h3Mf�:%]��Qh3[�VC���Q�\�%�����
f��x���YyPD&����l~�3^�J����6&SOC� ����O�P2��� �%;�����J���ě;�]�,~�\q��	�)���
x+��x%,���w�M���Yݟ�l�T��ѩ��$��JT�,AJ��*�ib(�L:�O�@���W����}�T��̮�h�pT�D�6?��� ҪxCU��RXP��}������c��eW��	W�7p�d]�cZ�8����W`N���3O͓�򙢭��)��>�����	��䑹���i�B�ڹn��T�Wt���J�m�9�$���������˺{{*6ۺ�ߵ��o��ԗu.mj�8��Ɯ5+Ub��Ϥ�|U�#�1�����%Ȉ^��9-4��>�1�S:�p�I���:��o�� |�gO�T}Fy�=�O���d^�@�����J]-P��cw�� ����M�:.��ZH�x���d#��
��K�� �� H2Yg��H�T�Ԏ+�F"�X/j!��;��N��`��d"����I*���<�3y���D�«��pԽ��&T���'�t�tT�}A9��D8��e#-��0���v�S_�9�'�� el�L�"��/ǎ��I7�� Lp���8Z�.ʓ�c����Xăyw�|�0�w��TEY9)�"*��{��0z��1<h�� �v�	�X���ʗ3��jJ1�,)�I�$�8�=G��o���H��b�@�������NZ\=˂c��6�H�8�?1#�	��M�-����lv�lnɸ�=��v��B���D��~C���Fa~7�3dW���~w�c�j�XT3qP`�-w{��` �S� �ש\Q�����Oq�d��䶽�˰�uL�`ON���\�n��&��E��Լ����8�r2��������6�!��4�f�$L�M�����a���u�?c_bk�w�ȁ`2dةjqҷ$���ު�#��Y>�I���ˠ`�W�m��~16�+�s��4�ĀF�%��r<x� �ƋƼ!Dֳ8����k;����9�������e�S��^�s����=V���݃wɦ�K��t�G�}���<{�F�e#���1��Lh1	�!-KE���o�)�b�6?H�ؒ&8��GǞ��j˧��p��V�K_Ć�6�1jeL.�S4!�v��^۹�l�� A8���R�\μ.秩h��@�.����� A�!3�v�U�8@G�	2�_f��aX�����P�G%yS�SR*��byN��֥���$)�`7��謚��S>b/���,�Uh�8�L��هMJ�����lOiY`D/^���G�}��(���6��v�^�,ׂ	����D)�~D�X�ĵ�ؗDЏ<��[S�ù1���c��Z�����.���GR�8	�H�.�ʳ�B=������0�<�1����v}��0|QC��O�L�1ā5M&Hɑc�b>S�M�@I.3>����C�����`u��Y��PmLD�t<�t9Ed�,E ���{0�Y����3`k�J�SN�2�=Fb^\��7���"2���Q��An�\�$;��� 2I 6s�Y�iXg�Usi���+�/�Q�?��0��y�=��?1�ia1�{�7P�����t��n6���� �V����Us]��B�^z{kg|X�q�s�;P���t�3�C;�C�ڶ����EU�����:'Z�Q����|�+=9��6G�Y��C�]� ��dXݮ�CB�*S}�J5�}��0՛dK��-�3��ȫXC��N��1e8b����	�l5���+����a�z����~�ځr8�'l'�{M�'^'g.LM��,��"sD���R�$&V����#V�gg��5h�V9�3�ǐ�w�D%+��Xa������P|
������^Σ��K#=���^"�=���^D�V���._��`�"g�#�C�T@E�h�Y�rf��H+!����닾2y�6��.e1��g��
#�=Q��1�"H��wN�F��.@� �;vVo�w�J��nv�b�JƱ��-�)�(l�R���3R�1A:L��a{�&�b\��ڗۭ.PtJ�I:��8 z~)�����P7�ʉ���ҺV�����?��F�1�+�.���1�	X'��	#�wq�g�c���/p�\B<��m��.��`p籰֧!�V,(�W�S�bAx�D����&���S�c	s�c����J�|� ����R���+��1��h��nK��ʑ�
��9��ْ�� ;c*����E쥄��0B��$Z�lX#��qզ�+�v�'@5���
ю�4����J��I,��D?���e�i�gF���Г�ּ�H0�@�r��1���LN���R �$��Q=�>�	� ����X�H��u�UT�C��4ywbd�ۦ�����w�\0�(K�.rm�I.c���]������2�kB�]>�m��$�9���{j9�S޾S���i��'Q�Ҫ��G���\f� SKe##�ni����m]�_9�H���ڇY�Pu��-��G��=��%�����60���c��?����#\���ԧm}1�����q�̄����W��7���G���Ȅ�64H�Ԅ�;I���{~
���E'��񒷄��Xؤ�C;�w��]��)�gVڛ[�5<�[aS���w_�O�8�0�&�Kӕڥ���m��(tr�����N�4��}��I�a�?�kO�a��h������՞kė?'�=��x �%&�3�9��A�c��?A�D��Jl�4�r8���`�	-5zvǃp��T<��{!���E��C�\�%L�B�>�&�ؿ0i�ݙ>�agĺ`��;O�����AD�@qry�>-�7��f13�B�b�L"��s`	���Lv�놻+��h�$��3O(��	$�dn�6� �P����{0g:���0� ��v�&l�*�;LW�_���������Ɠ���:^��8>Rb�]��!k�X&H����ܘ&�c,�q��}���C�S�;�����B`Z+K�@�1AZ=����/�M��h2��]��3Z�G�r���)g*V����
B?{
:n�qq�Z�nԝH��%W�H��
Ljd]�n�~�圸�g�P��;���Z�7,�T;0�!wJ�.mA��9�I<Cm����l�PH�$�dn����4+�q��������oۦU�� A��+�$�۝^l;x�h�J�g`��w�0��@�jIW�}>�ݾw�����-6�>�q��Ƞ��(�`�ۣ��b�.��GFQs�V���4t6��O��{�w{2oяW�7p����#褪U_L��7q��i6�f.{V���y���:��K9ǿV���bq�T:;�`��"�s9��(y�%ޢf�!�"S�t:�{��>7����RVY�`�x�s��|RҎ��Hk�D���w�,�.}>B2��Wq�rb�>��c���-&'��O��]�����RA4m�\P��k�^�k,9Q>R��Q��Rm��o��x��{7�Dޒ0���RwV-8[�Xs-��8:nUa��`�'�v�>��Bԑ\D�c&ʢJ���~�;Zy7(NaVц�8��:藙��xr0�q�M�o�\�*�z�J"�K�W�>�#S������L9K�ʊ���i�sO�~\���<��[S�������2bw+�]P)r-v�\����0?`�(�c������B:������Hhf��x ���-���ޕ��F��ݺypW��EZ;�B�.������q�3�0L�@(o��b: (�	sy�7H��N&������W�;Ж�@�Q�9��m%�� �ˌo�
av %����Q���}��B�1�-7�zn�-���۝�b�V��&�������L��F�y�� ����dh��x���|�f[b�˘sF\G�=����n�AdZf�=�!?z�b�ca�}*�I!�Q`�!RZi�rٕ���b�6�I4����������fGe���Ul��?��v.�nX�`,�D5�[t�/�N2�
f(q,���e{H�W��=���Έ�)m������u�ܪ�9!ΰ���I& ��,� ��QmW#���*����l�8}|֮J���Ql�C|��k�`�T�|j��,����7�K��9�b�Z�����/_H��#���=f��{P<���
}�T#'�v=`��>�b��
�&$Wx��ZǤ�W�@�t��~qW�e��<�>0ً�{@%��s���e��J�r��w���x!�f�؇+F�^'Li�S�?����-�+�{ $gM6����̓!PW�p��`>�x��F�ίZ/N���a��_��x��[Щ$Hλ`z�FC�)D�_��Y���9�9����5��j�k68�ŕW`Ω}<�Ex����)�L���� ����
N���MA���Zr�[8C*0��9��RҦ�/ww]<���D���.>kI�P�w�]H��^*���&PW�wi� �M:��-#�����*.�|�St ����a���;���'X�vIۻ(��gJ �^.�ܣo�U0iw�{�j�Ax����ĿDk�:��+�����lE�����6�H�%�6C����֊a`~�\�Ƭ]�#BtM-�7�7�cJ�p�С�8*�1#�(8�on�`��f}�p�kT����[�S�cH�e�&h�',ײ^�j�ъaݴ!۴c��SO���+�
�G�y̭�C��z� &o���IJQDaSC���>������?;ʺ���D�	_%vw�?4s���׺�{<9|oF���,��!�-�<�oTg��/À_X]�+s�Qp��q�����q}~(�u�Q�+����v��2"��'�h�Y�ؓ��3����J�Di!*qC�8��!��M�`�h�����S�UV�~�+����#�]���Iu��1U�\���_9����:�H��c���gk�j5P],��8s���]����e���W�J>>��ڧs.�)���6���x�3�4\�"�eB��~bײ/n���`p��_��ತ"U��&�ߙ� t��Q�x��Z��$�����
ޯ66<��+5���O��S�bB��Ec��7�l�Wj�a����e+�^��$�U��6a͖��N�V$f�7�:�$��g1�E�=��V�g�T��D\�8�.Y��=ɯ]�UMϓT&��Y�A� �S�Y�G�9T�leYK�m�n��M����t���d	�M�;3�_�>�i����t��Xm�������[���ߚ'~�:��G�`�**��U�E��/8�^7��E�$�`�/^��=��_����D���s��D�����z��>�sw^�����j�����$a�3`z���C��]�m�!:���+��h�h�;�a�~N����a8|r���[�����s��e��;E �a�I{����o�Ęd#M_���.�bڛ �ȁ��U��8��T��:h�=�)g�)�эch؜
����q'�n�}��LD>8��D��ӄr΋.�-b�tdGiW,����kP��N�"/��,�r.�axm��L�냹�#�fpY1-t���Vg�}̽���_)�;$!�1�����+}o��x�/��y������r�O{�ъ�#=���D�43��o�[���DE��1����H�<�'*�OXN��HA��m9c��&ߐ-/w�Z5�Rr+��KU>s%���۟�Q���~�c;�:�9��09���،E��-5��T��l��<�ju�h�F��8�u���/5���BM������1�9)'�!1��T�%3u���|�"沖HW9������2M�S��i�o���uu�H��*"W,~|�=���9C�D'�y�6#��|�¸��'
F
���>ƹ�����J�,0��7{�H;��韒 ;�,�Tۺ�m����sP�����* ���(.2�1������4?}K�f�ICu���e�q�G�7Xcn�D7sy�f�����oIb���80Vf�	�]��������(^C�R~*_+p����'�Rd�Y�/.3;��3���4IW���}����˦�U��8v�����/���a�0�����w1�n0HK�Q�eɽ�	��YN��jK]Fȯ�Lb�sN���: Y� ����g�]�y@���q$�b�@a���Ue�ݕl�\[D�Ss�L��X>NO����A���n7]�y\ �y7���{��#zb�v�%��ٺZ�L~D!��9��UO:�4VWt
��{�)�\���}��B,�V_���4���C����ˊ�8��!0�W%nx`İo�\�(ND�ȟC2�Έ8�U��I����Ng���o�aX!؝�?I�J�����9����f�uYVޥ�7��^� �������W������;��e�,�s�m���;�٬��D����)$�erg�+m*jB`�*U�e�C�ͦN룷���I��[x8��VWz1�Y�c��I|.�\�(���9c��d�qlܪ��p�7�������?0J�76�y�dd�r�(��/�|���U����j�C(M���/O
`������3.o�Q���X�Sg���ѸMf�Ϟ޹N�B}����$����&�-dh3��y� ��`D�-�4���Mc��k��1~��>�R_S��{;�"]�d�����\���O@I�=dEx�.W�<���b�k��l|ھO�;�}���rXJ�������9�T�]2�V��9�DY�"�e��5���ĽLI�*[���|,m�J�xZ��(����5��a��i�}�.=iaKN|�	xJH\�
�p�GWz['�f�
���H_����Bo���:h���h�t�|����c%�������4�/��`ç��7� �4:��;ڦ�OeK�.X6��wv�qt� ��c�]�������$y�K�g�s+�Lv#�t��A_�y񍿧uy;�&��<]��&@dp����*h&��$�����<���^q��H��x3�|�V�L)���;����w�;�G���/�`h�� \m�\_��N��A\��Y�Cn�N��%\��AM�j=�T||���j�P�k2�Q��$�kv�|��}HK�5���O����̌�FP>�y���f���!��j$�������bav�J;��Zk�Kp�m��v��M2�Bt�Dcs�~g��FTL�<k�v-�Mּ2�U�bx�cBd��A7l������ �'�D+�6�+ �ȷ]��U�Q�4#e��d���9���\J$1s���'�p���
�~'��q{kҢ�0:S��A ɔx@=�$�c4���5�p|d����t<Ñ��"^F6Ӱ��U�mv�� ��khw��]Ng��*F�B
|���Oc#�ztR�� �O8@�o��9ᕏt����� ��uo������Xߩ��{{_���@�֛9R�h��_�h����D]�G.J����.5�Y�A�GP!�����(E%\�nFft����j�ڻxr��F��Ύv�QgN�����ƒtEkRU���:��d�q�|�����""3o�*�u��b�C\u��7<����+
p��8�,���Hx���H��D�F�P�G 聴/}��?��G��Pv��2T�.ȅu	d�b���
o�bAG�D?
�Pf�,#v^�a�F�J}�3�nQ��ޢe�g;qI>�!*��>��,���f~�M2�FLC%�a�6ڿ:/�������wbG����"
�k� -����"*���ج���m�pE<lG�s��=�U���Cqz�����F.���;V �|Oi��ɤP���ϗk���c�
��Lo(cD>Y�5cV��hg�s�4�!4�/W�:��Q����<�M���چc�6�Ɨ��z�f����1�\�>Q�X���(?���Bi�`#҄��)Ze��n�ċj	���?���::�Յ�d4����3��� �6o
��2�����3V�y8��E���[�wo�GG����ܥP}�Q���^\�2!:��[�9��>����x23!���m�P���L��<o	+�-��h��53WN!�ԯ�7e��js�"�@�[:Fۇ�e��l�����A ��HN�k_��[^��`��X�40�ȭ���o��(�P��x'���ȴV}��+DFߒ�Q���iP�4~E���hNk����v-y�|4(M��´m��v�y�	r��ڛT��s=WR�UL'�An���8����7�@ԛ����pJeT���)�:�e/2QQ�����3���$/�i�!o�f����VA�r���=�&����~��� ����PH���Չ6�� ��������p�Z��e�"C���z[�����Z�en�����y�!ҟ��kK|�EO��-b�N�4��V`�b��3�Gp�Μ0R_�&~�T%ňAV�%��On����]����fC.G`> W3`�E���v�h�.����
b�y]א�
U�;��]?`GAi��y�a~/*0� n���/��mh��*E���6~�4����jq��Ù>�#v���,��EO�����C%r S�j�b�A-���PI5?�����^��4��X��ͩ	��W��Au�͵nQo���j�8,ˋ��@1L$a��A���h35��mxw4�_�-2)�ߖ�&�)N�����  :��#��5�W�?d�л?�7p2��F�֠>r}�&DÊ���<5j��X�m�98\C1oHXQ�R�QQ�b�:�(f5pi#Op�sr��s�<�/AC9�=!����##`�(_,x�.?Ye�SU:���$�/���p�i�3y�}��߲��A��7@ٯ�$�'��,2Re��MES���GMe��z*����Q+��6J��X��r�\�:�g�X�Y7�k<��H�l&M��8����>���sf�U��?J!}&_/�R��f��8~Ȁ �R��_���_ؖ�╅ƙg���,*9)��C8޽����{D�W�Q���I%��!���u��5ѝ�J5Z�j�!��C�B�š�U�\0�9&��̚U�=f��h���yd�1f�������*�^?�?����Q' a��^�g�*ك<�T���s'����n䴡=�� :<�6Ώo�@�'O��tRn�����c�BK��v���<?C�5�b��TuI�U��^r��g�Uh�j!y5E)MM�g�+号[D@��jջ�:BS�. 1�=n>?˓��e5��"07�So��푕��0�81(���d�=��:�fc9�1�m�ܪ�(n��v2����ujX^��p���w���&��(0�BM�<Tț�$`R)�X��6r����BF�u�CNK��cġ�a2�Z��b�5>L��x.y�H-� }-s��@�J܋3����P��C�)��<���,P��3K`����Y������Q���e�z������!�h�0�=-B>�"dK=��f��Ŏ�ɖ4�����FJ���s������ɺ���Nbe��c��38/�F�^�b�� t[�k& ]l$~,`��;EḞ�N�/@���mC	��FFX�0C��<E}�o���rĸ�dvwXFI�S�����ǁR��ini�[6v�ma'aL{��y����!��� �i>%vT�3�Kyc
ax����o��Ɂ�/Z���	<9�R�g�i���밍�%Y[<xI%G?�v�ua��.�<$��A�}���J�#|BEB�&!	����2k9Р���3��g�Cq�c6��kl9J{�~^�Ǵz͎W.}:����Qz|؞���䝦���v�$�ڠ�y��#����V��.��ի�Qe`�a}��0kk&����������1�N���'5h������X'9GZ���5�`\�6�T'��+a����U�8�h����Lm"���G�������\���2ɚ��|8b|_��h��2�5>�/��O:��:�l��cﭟ�S��ܥ�(ʦ�0h�Xf�ki�G�!�w"H�{D�a���5������V�F=!��W�xN���	�iM��GL{�l1T~Ȥ R|�}�r)��2�c(}�$��F��v���#��P�@���w���s�VI���K����R�n���Exc=�(��hgɇe+��B��RL$�ôd6RT	Q#aVOX_���j���E�����%���9�IG�V�ث���aw�39	�=�n�<�*MX��V��ȧ�TD�#�{��9���~�31���7K�D=��9���fxp�_�b�% 7�P�2h��v�c�v�6T]X��{���ז�k��Ba�R�w�=~�;F����u|:�q	��a� �dlB�B/��y��s��)�'�W�	����֘��Q.|��{��Hٍơ-	=b�p�g�y�m���|o!ʹ��"� �3TE�?�n��R�l��5�Hc������ ��~_L�l�v��,w� X*ᶜ�[�%v�r�c�/�\z��b�r�!�wI�?�z��c�R�˧k<S�={j�q=T�z^�r$@��=����itX(�>����|!=
pT����I��jCj9ձ�}	����K��K�Y��E�玀tL�˕܅�7�^Q�C
����W��l��W͍��Ŷx��d���1�>�w@P��8?wl�9�v?���@;�-ꈧH&'��<;Mڣ�z��:>zn�R��L?��U�pv�یkOΘV��r�9�W���mdBBz��� �-�(�X�5k�ubxq�:���%\L�yAO�����&0���Z��z��xvw��A���.�2��٣+���fvй���B,��9����p�̳�0�P4�7�7/��x���tF�����<�g��N�d�yɂ��![ݕ-�^��И��}L�AU�V E&���,�h�jJ��+�/��:���JS�T���7m��*!��9pk~L7���j�H��C֘��0""4��y����ȕ)��U]Tn��\C�t�f#��Le���c�����Q�ۙ�6Xi�luTbF��:����B���A��봦���*�D�X#�[B��S���Y4<H	w��;B���݋���_I�i�יI�E���NR�R����2m[�l����
Ḻ9"��I�V���D�R�Y
LV��Q�n���H��~[�11�c��X�����ߧ�y�|-���ek7�g˷tF>�$�n�ưj���"Y����ʡ�/�B��#Bt�g9�g"IJ�'��C�6�N�[�����[�>��2���m�����Q3�l�^1�;(�ё��^���e��g!R��/�sn�յY��Wɦ��o޼�Z��(B1vZ~=�V��!4R���V!"�Z`괽�"� ^^�D"|��O;�-.A�C�@O�e�����tv�;�zμ�R�h��0���_ejѽ[=�Bp��!�N�T��=�S�?�6g���5��i8v���Д�>���� }8{���q�������c��:v� 2���=o�HmIa)�PJ]Ǆ�������0��)im�|nX*xh"8
1�-��()c+!���kx?��*Ӣ�x��V�> I9H�� �����ǟ��jP����lu��jݖ�\r/�I��?2XG��<��R*��b����0��>�/H���(p�U�ء��2g��w��H�B�%O9_l}�S� �OV�������w^C��%}${�G�~�3Ă��]wn�\�x��Ak��6&�qw�ĤiSPRWuќ��vk�� ������pc
��Lm��	�������ڽ�3��X��OMO,et���- |<c���l�9Cq��4]6H�	�XȐr!�F��Q�pJ�{���M*=EnZ ���o�5�iEIp�mo5���R��H���¢�>�Ũ�fQ�T�f�>���+_+z��������˴sP������������GTx��d(}wjݾ���f4�dfNq^�6}��l�wa��cpV�V��N�.݊���� ��!�̹��������}����C�+󩠛 �
�U�%��@��g�)�IV�7�'�Ak���]O�"S��l�,'vbw7�4�3I�n^�#ۚ���{���T3[B���5����]�}%,WF7�3�?�T�ɀ���!��^��~kB΋���wp����y2Y�r,^q�2� C���r�g�..U��{�:iB��{h�p`%�_
t�����h�s��L���BZ͟+�F��&6�"+,U�3u3Uϔu�ՅL[fJO� L��b����ю�\t�,�S�lLu�M�X�7p�~bĒ_F\֪�"-�솷L7����=�d����g����惲J�B�����}i��굉�����Jd~����I�o2���d���Hl,�R$����	�V䜹T�<�W��ؓ$���i��^�kO��< %��/I߳����ؙ�x��>���J�|C9Uk�>m��~���
m���kb�]�)U���Ǟ	:�Qi�"\���$s��t�Z)h,�4���b��X~�� 6�:*H�M�zbRvk&�(��M*����G��F/�Ϊ 8G��l��`��I'�Q	��W�r
�00�����������&�_1�	��r���W�ԫ�jP�A�M��rr�&\lC�;�gerC���*A1�cG��TL4LDJ�F�>sA�L�*�L���H5�LVx��d����C�&���L����&+&��*�F��
���b�	����n=⪚�X���*���D���_��g+tS��ha�aU��}*�E��Ӝ�R���i#[R�P-N�ĉ�`����;��� EG��=��V~ˣzw�F�%mȤǟ�&a��f9K
"Oh����y��Pa	~J���v&:���&>���{��$M��e�2��u�Ib�7b�C���B��N٣n�L#"���R%�C#�dl�*�+��ٓyd��Q�iH���1���U��^
]e�z<l\�J�(_�np�������tyN����C������4��ꮢǏ\�)ނ�B�ө�4Tf���͜ t�}�Ĭ���x��
<�۶È�A���.>E��m�K�2$��V���(��\�AP����}��X�qRרڬ/��,�X�_�]s��`r��7�#�z�F�����Oŋ�}�����T����L��%�B[_���<F8mr�v��Qp[35`���(Ŋ�:H���A����bI�Z`ӘC��h���a��쯌6U�x1S�x���O�.���r��>�m�)����F	�DDz��#�~�������q�Ak�g��!5�W�"��XU�(e��?�Q��Ԯ�G�P�;]�lȥ�+���+�� �K:M�YZ���W�LO�;p��B�J� j��N�ݩ��t���t�%u�.Ԁ���΃�;�E�suRH��'M>)#��� �*g�i=?�$��m"n>�;��aԞ��ޒ�D|��ݙw5�u;�݀�:�ꮐ)f�H�B����Q�Ӡ�0��3�%?�.�:]��TƲ7Bt���ptᮗp{�VV������j̃�̴L��^�B&�aq�߈p�i�	%�>0�]��QY����pk{���Ձ����ʦ5�+Kix�p�yP'�Ԥ�sT�'��������Q�qȱ�����@s�gerb�0[g�0U;̴�Y�^�G��s��7��[;�_% -���@��f}r�����Cu�L�ˮ64FC��cjE�~�w��v�T}ᑡ�T�#��r��M��Ӓ������Ge,:�����t�ށ]�W�x�]i�Ťk���s��*��o�U���uxNm�mJ-�$a��~َ?:�|N�$$���`)i|6+�����y܎!�eJ4Rۿ�<ԝ���Rl����0���M2��;�����nP�{�xB�!5��(��et����S���9��ڍ��\ c��,��Y�ʝKA�5·L����t֥�H�r؆>D�9���Q&�aY���T�B&k� 
��$1�|my���p�����!�R�s�i++U6�A������JE��纨�b�V(���{�*3���Ip^_�W����ZhuX��Z]�o{����X
��ڱ���Tw_����h'�#OzՔw,��W�9�SQ3ϵo.�b������g�0g�j_����mRة�g�7zz��fjG�+�M�I̸;9�&j}PZ��=�jC��!3��	�ͪ�H����cJ)�Q�����^�b��Y��ȋ1�z��W55�Q�g��C�7��?���Č�'�l;�y� ��
����>����Ce�_A���i��R$'X\�� 6^ګ�(���A��wT���Җ�b'�O��<;~�����.�3/�n���c�ǧ��kY���#bG��^�C��'-�TH�� S���\7�T�?�g��؝g#H��z�����6��i(�!󚟁y�����밾n�_�l\����� dG0V��	B^�Ba�\Ǡ���q7ҮbC�%��_�����D�A}�Jq6_A/^�s�}N.Y"���+��y�M3(��}��t�On�=�<YT&�}���?�ZX����<R��?U� ��jXu.n���ɪI�~i��u�7j(í�_T��1t�:�{�<�į��q����7Ҕ��v0u����U�5)�j��ϖS����K�]Y;���:e�l�s~�=�)���g���_1������oYYD����4B��-�(k�>��^"rU�u���d����{ Q���G��S<M�� ��XE�_�ۚb�w1SB�8Lث1���i��N�s��tGv�Q�3hV���%�ݔ���>�]e��F!�[�v�8���1��]�����������Xh�VE×Y��פ��������<���.��&' �1xy�ࠧ��qH���e��	�	�lV��g�m/Wo��X�a���X�M�M�߽mn��FJ(�l\�W�?4��|��d�3�Y���9�]�4�j�a	B�֦/$%���h���z��,	�R��G�*��<�$��z��+ǖ+��l�៻0���|���οSorA�^��#L��; Œׁ�/��Z�A�	n�O�-_��x�q]g�T�a.�� ��ϸ�[�ep�xd��Um��{�V�b��c�t�9ܙ�����H�Qp\��Ԅ&�)uR�;�@u��00����5x�1'���M}e�0�7�%VƖa�ك7����ʦ���P(��I�0Y��q�����D��y�9�b��s隰���BR:��1� ~�cЊ�V��#���*�t�+���S��&gw�̯o�ҩ�珟è�m�a�����}]�CCg�C��/3EOR���)6��)d��N����o|���3_��sX(<��'-����J�*���Iz�����Ar����a�����E�Py���/j/+�m���'����j��|)� QOCݿ�t;��Ͳ���R�?�F�vO�'rҟ�&&�(#����{q�zU��A�Z��_k�L���T��A�9�b%Z���G�� �1����CH=p�\(�6Y�3���g��$ȫ�d�7蠤�`nM>���Tc�D�d6Q-��T<��$ٯ��������XH����]��1��� Hi�������+T��?���%�>���zW5� _X���x��*�ʩ_ó~�V	���n��O�c��l��j�����"��C��ggg�O�^�9?���v�VᾺS@������*��x�'d��z�M$�16i�Bbs���z��L+�.�R�3,zO��M8�)>K]";u���/���o�zu<����r�B��G �r��ŚJ3��%���qg�4�� 67O^gb0 ��2�~=(~�o0�T47��	�&��~,���U�p�N[��S�s'�GQ|����;	���5�`8�v{U���ɿ2��M�3��Q�:��(�}
b&�=Z�nT���uNh{�K�16�v�T��E"	��8�2�~Dq4���D�����Q1̲ʂl����f��Ð%>"g�(".� .�¼���$�,i��>�a�vX;�ſ�*hdS<��r�gn|�]�͐"���1��L�B~��z	Ʊ���+K�wEPI�/lCD*ok��,�ym��^E���
�n-�H���O �t�]���7�㍌�7҇�%o�}� p�*���E�VI�I����f#�6 N<���4��U��Q�%�B��|y���X��0�Ug��!�A��X1�Y	X���N���(Ƣ��AkZG���}��i zYZi��䍽A�U��'b�X���7�d��� \Oַ�4cޟ����]�0յ�۝4c?�>U�K��@G,/��K��Y~�/cp�{^�y�a�0ѿ[J��6p]�ൢ�٦'������a_��0z��97�A?�[�E�Q���k�x����G؆�u�Y?��JK�7��=�$��ό^��m5�5��xzC��[13ߚ�yߴD�q���T	�/i�Q}�|�K�����k���L��*W�A��,,I�5ӻyJ�-��C�O���q��+�� �6_����p�k�X���og"�~���_L�G#�! �����/�_Yo�0�F�Xp�ԋx� >d��~�L5e��r��ЄE���f�ڤ݀��W"&��C��*:��qG3u�0"�5��9��v�G�㙒=���u<zMz�7�[��,���H���&��3�:6����_X��0M(��e�0��1�iG�[0�ӠB��Z���S�6э�.�	�<eݖݙ��F�g� ���vf�C���/�Ð}c�Z�!�k�%�h�
���(��]�Gڒ6}Vۢi��k�2��)7D2%86<��/Dej^�<+�����Eua�YRe39OPT��g�x��O��Ο�3��	Kh�b@yǝQ� ~)�y@������o���P��Eqtȯ�+h)R��������f����b9ös���~Z�̙��=�PλL� �#��iue\ "?C���Ҙ7��cf�r�	�Y� ����0����G_�[z޹�g�A��_Xє��="���6�z�,6���`I�E�CFc��xs��xG��n�e�
<)%ň��M�E������:@�O� �)��f����5���}�x�3~-lx���6��i�?N���92�N,�rh�h����d�-�:���8�?dh�K<}[�� �Nw/��$�dZ�76mX���00#��5
3�	��j�pnO��߬�W��)�W��b4-DR����>�h�Gy�X�O��=��-�4�pCx��)�7�&��%h_ѫ'�Uˤ̰�_!�ybm@�!�ض�,����2(�T%��gzj�����&�v7H`$�RZ�0:I���P
tZJ|�ѩP�6əV��ٔ�<�-e���+ն�I�a�@��(����T��Ǐ���ˎ_��ؗ����{��c����&�Z�*���L:� f��G7��Q�K���>��V��?6fN��/`�q�����Jh�,#rq�t�4��7, ���(@=��n�.�4i�I�P�l��MZ��D�,�b��_�*tS���v��<�����&� ����)����dt��6bMY�Rɳ�h�[���˒�yf��Ho�g7Z'eR��]�7��Gf0I�<�Ě
*Y�,w���bwh00�����dЗ�<;�	�n��7�5 ��n�%��&�O�i>��rE��F��T����}IR����dH��O�Ӡ�1�B�ό�ԥq�s4F�<��C�M%a�=Ҹ��M���[ץ(��B��G��Y�ܩ�N��ݸ�<�b&�f�q�.}2���2�"�}��߭��3�u`��k${J(K��iV���V	�#����
���A���).�§e"��nCl��<
��[G�VI>)�>��v~uZ���|^�"iξ|���cy�4�{.]�ҭ^1�Nc�� Z�Z���G�[������A<��V˓�[�I��{ð�Q�X����u�S7�CˆT�R�� {��eqb��C�����OH5���EN����/�ګ�8�i������s����
�l�f|H�]���~�/NOQ��n��~|�ǉ��r[>0��`fl�GW�+����[��N�|G�}_`�s|�E��"T���	6Hpf��Bt��_��\/�;~��*�E�W�S�F!R��z����jy���a[��}�@q�����$���(\�N�'66�m�C���F���|�t��� ��o�J���4�TXS�@6`�ahX�}��d&��埞�� �E��M���yƢ�� ~���}�	(��5vG��V����v���&6	�)'��d6_�cqAD��֛�j��g�}b{P��L�o5;?(�우�C�=��g~�Y��r,~�koB�s�8ԷR&*�Y#	�qV�޼�Xv��J`���}#Q���AFxj>�AC5{:Kc��7�|��%��!��)z�\�喨3*2�b����(4�+�䞦#f.�E���� Z�`}��� ��^�`Gϯ��fr�R�H�߭V�O;��訥GH�K4V��2����-�:@j��>,?�<���{���jz������*�ޢL{r�6wF+�z,koI���g�h���-�ir!���6�d���,�6T1ݺ��y��4�|dv��m�ɥ�+�G1k�0�������k������1�#���"��:b�Q��9�1���sԾ\���s���� j�}w�������Ԗ��w��]J�L�<}ݙL�l�`ɪ�o.��´��A�`� A��^�^\��M�<��ƭ����"XL�)Q��2���+`3y��Ce��T�F \�G�"��\z+Lu�V�u�%9�Nߡ9��+NH�����ҟG����\��&u��&���ok"'���Q��s@:I��m���U��Pc'v��A1�K�5�/F~�ؾ��r����:�.��	�p{+��dT�_CL���9y^u]Fݾ|o�Ȱ'M����vW̡y:���_�2��*=�M�V��d�{'�yYʋ���J��ZΡ	%�3�#�NCg�XwR0��6��g`Z��p
�,�sI�ԃ1T��xd����h]5ѷqJaG���&u`A������ly�@�A��3��Q��S��҅^L��\��nw���W�������Ux�����%fG<�YL�� P	�_c�
{h�\N~���R��F�48��J�|�����It}�L�+8E�r3�Q[�؜�F�l��hw�<�����"� ��I:S3���3���;s��'1��wU��x��&L�p �L�]� ]U�����wt��I �S�RH8����ڧ�3�~���䝅/��ǘ�յ����n�W�n�JY�2]�����v������۴� L����X�OX<��~�n?[������3�{�ff.�Y�zxY���7��Z���exa�R�	�|gI+A~$H��+T=t�|��Wr�r���dή�r�Zn����1�L�,��M�3�P*,̆��SX�����$L�\l��d�LI6�㿅9v�v ��=2r�%�j�����m	DF�����RTȏ��'��W�+
r����܉3p'����̿}��-��}���Xy�P"-X�+���þ%��yI
:2Wn+���-%�������5R�L��l���e邾�Ah �A/a����V�;�P͎\�:��UӤ��:���R��#��fP�ũAڳ��t'F�><m����ٶ.�;�36��GsJ5��Nsr�$g��F�U��	�~��[�h�j!�P�ƣ�o����ܫi �&��S���|�K�甤G�Q$�%�i�u����_���3`�_�x�3I�ER�"��Vb��}m��^�sƹa"��@Ƥ!�z6r�~T�n� �9�g?���)z*����	u%yl�>g���p�ɜ��ٔRv�����hm.��o��_�Z��ᷩ���Ћ���b��I*�{�q�I���SH?|~�9�-�0����������.��Kfm��R
$X����5��$^��u��,+T#YF�ԝ̿�K�S�:3q��[�{z��8�$%���R����k�&\���镥�_L]�����v*�Sk�<�F?��E�:����6�3�E�#��Qh�r.8B�G�m�K�ynN�y����uw�����[��{�����(X�+(����x�J��ZIU��j��[����.���r}^ۺYA�dP��� >�����Mmm�*�/Lg+�85�|��������4�Yk�eJB��7�R�=~�ڛ�q�R�7�n㹗�§������sYm
}){��8g����B����y~�r�pi$_�=�h����V��|j��-�J��4��*�K��	� ��w6��d���q���:�pF��5��|9��˃Zː��k�e5�f%�"V7���������H.2�$�2e�_��b���^����A
.�s`4p��7��� 3'��]�7d ��7\��p4s ���k/�Q��&pH�D�y�x��<b�s墪9˜�Z�� jԈ
��>��~���y�=請�}g�n���AnO���D3�ډ�i=0�J���Y3HrR���*����G#�������3���i��G	z��Fo��d7�y���F@Tw�v���(�٨��1������
i�8e\�Z���R"so�so�ci�$�1=���,�
�G~r#�S�!a�M�ξ�,�pDi���f�R�/)P�:.���O�w��/�[�T^�t5t�N`+��ۤ�ci�-9�`9�5E���4��Mf�ӈٮ���'\��R�=�\�Z̷l�-�>4��:)h�b�;�.J�Xk���l��{��dx��`�w��rr�kZ/�3 >떑�a�������@jI�u��c϶�q�����v�R|�\�L�b�0��	{u��m�b���h�˲����[�o$���X�U�ԙE~1[��ٖ)�n�HspĹ�?�f,�C�&��{`�V)��u{P��l'�^�^|S�0�2���yQ��=�6z�8%V[IF���\�/���v��糝��H,G2�{��s�w=�q6��\��KҲL�!/F�}!h��C��p�����[�Ӧ,�R2�F۳����a{=)E2�NKq>j����b�ǟ�L"E4h�V]�-A��9s�%^fe�jO���:Ӷ����0ռٰ�e:	'��e���z����DZm��.=W���6aR��95���F'���#KH��;e��K#_���|���HM�Y�м��EN9Y팟��E&I���ٲ�g�(�V4����A�"YW7
+9�P����f�[)[�T��1{�
"������/\��A�>٨�i������~���S���x%x�f�^D��0x>����ܨ6rˢ ;==0��W%��<�Z{<G]"�~@nC;���b%w� ��$�F����Ld�8�+��_P��,0I���*��Ҵz��'��M�3a��H�il����m0��ײ�Y���&Δ<�
%k���s�
N�<i�.��Gr5�ȫY$G��4�4AT�������Zy�v���k�>qR����E!�b���^�����O�o��]�\���_W�,�C'Y�rڋ�f/�=F_�YR��)h2�����r	3mZ���wx�s&P��V��-�i]�#wR�h�\�k����*I��e���o��,���$�ЯF#QR]~�׭�c�5f@&�kZZ��+���H
�tY�/�C�V����[�v��}�^�x�#s�%����]�Y���4~��{��?@�����[Hf�X���	�^z�S��cg@u>`�?�eGYSƬԶ��1ޟ;XYX;0�N�-z!��^����t�\$/����l��[���t��Ӝ�V�k;n��7G�8�"h��$�1dP��0��z��z7��r��Z42�[�O?�	D<�ܿ�:�gw���c�����N�o�̤�p��߁"$ᘡ\bW��qi��cj^�Y��<x��1�����*�U9�u�����PXvSRd\����iD�
�M�g�h���fh$�H{zl4 C��V:IȬ��kC���vf��~I�/�)�Mi�jB�b�͊��L��o*;����o;�u"�f�ꚩR�\0��:����zPp�D��Hv*���۰g�[�B n$�FeY
�:��J��.�a������E���0��P��Y��W�>��Q$w})�Y�r�f�����Ƈȡm*��o_V�K�O���B��[M�G�w������/#S���z,Y�h����%n�~ʓ��Vd������'��}��E���p��q؞3]��v?�������5 �t�^CXFjxk�>�E����1[㖱D}X�H���I�kp4|��M�����w�GY��P���3���E�gI�-���1��5���o�o+h��<1�/H��[�'�pm��SE�%�U3���>;<L%2�{�����!c�}z�0r��#�˛��޵��M�!�C<��㿻7K a���i���m���h^�(�|���b��'��K~Ѭ���OzE���<�D�G������C�׽,�~/����Y2�b�kPFTA�\\1TMg�K�8�iVȩV�;�s���e�M3��;_]Ǿe�{�W�v�0ԭ�w
vO�����\X!l� uy�"�ˀe�*�+:���ч�^�Ϧ:L䤞�dT�7z�Z���z$��,>A��lȖ\�U��O�e��k��Y'��W�b�~=�O���_Y���R�n	��E��@R�<ʹ1��-�P����C��q
�:97��ѯ��i���*���sdV�w�F�e� l�%f�_�o��K�ҡ�b9c3D���Uc��Kǲq�y���
�k����-ȞȻr~���n[$~4������Ĉ�{nifvOܡ�*��^	�����ɝ�$ҋgF�z��6y'��[����)	n|2tJgK���4<��?T�;#)8��(dΔ��T��I��Z�1)w�0u8�nB;糧	��#��J����Pؚ�~�b�A�����u�`���q�<��	�N�)����[좋$��2��9�5ꑟ���|�eh�m�2�˫��I&��RH�"���2w�*�b�ܙ)H �F���RecUy� ͚�qLP�Y$TP��P��T={������8.q1��L�cg��jTJ�������n�?�qן��ZS�T��씭͇royA�\�ЫB9��>�|s����)��s�����a�M������`��i?���9�a�u<�gt�[�7�PI�ȍ]�=�g��1�%��ϫ?����Zu������.	�#���*FE'd�D�����M�^)u�q�{قՉ�l��hȕ�.�oĩѻ�:����1yَ�c�)�������4�t��W��ӿ�L�ŝ��c�w�x.UM�=����$ќ�(��bm� ���̈����j�
���K�����&�4�׆���'ae����}�����B��GK��@O�[���V,�Э���W��m�L�7c.����}0]�L#�H�.� �d��������	{��M0+Ԛ&��5�n�D�7gQ��.FЁW˝ʓN&k��������ܲ��q�gHp7y��g�l��f��bɼ��ZI�R���Q���5�[3��w��� G������sS�j��in���ӭ���c¶s��iL�&�#�P֡I	����ն��\ݞ!�쳈L���_6��52�7��ǅ$�F�@��		`��
�E�+V��k����۬YЁJ"*����7����L�+s��U���92�9�;&NQC��qs�Ͼ=Mu�ڽ�W]<�D����=�W]j��J�w�\h�[���s��s���Yr��0��X�ɰRl��x-!��ɵ|�m�؝mA�k�Z!�s���DQf4@5�=T�r����o5Q �˰��ċ 뿙�[���'�|=���q#�G�@\}w�+Z�&HTz�2:l|2I�oo`��� A��%�.�&�M��&g��y�)K�t<v����Q�UW-��<-�#A�;Bs
�/�"F�m� �g ֚���E��a��҈���C%�uyM�M��LOʥ"a�s�[��������̤b�j���9��'�Ъ!��g�v׶�ؐ�m�[�Hܦ�͹��ڏ��ݹ|(��2-Wk.>��g�e�e�VO�| �*#�`x��n`K�������4]�|Uҝ'Ј�M�(Y�:#ъ"l�~+d�E[0GWs�v�����}���մv�Qa����WX%��HK�w����eh�3Ǫm��4<wX[#D:W�A�{�*��`f�G�`b��5y6��i�щ��AK��� &�֥����+�wV��;Y\G{���$G��WV�P��D����WT<���B����*�-�g��U1���ۘ�h�M#���g�q��
mxo���m��yx���U�*c�gd�D�y�<Uc�	�9U�q��BoOՑ]�ـP�,EJQ/�'���s��k=3���&�E���!+�Q�E�o4�Rz�W0��$ye�I��P��ئ@,Q�($��R�ܑ[)��/W��"蚧����(1$A툥J��q��o�#vFNy�����������T���45b)V���Q�w�q��u���6����B�}B���Ǯ���|�ݻb;�ĸ��YQM9ǻ|e��Ãe��H՝�f|�!A����ayq�����	҆$��(S��e���b�e<&戞����1�=��[zZ�P�>�S�l8�mFb�%��B������R�h%�l�t��Ex���xv�N5�1����O2s����j��Ю�xx���j�&�N�nD�t��|�3��Ci�:�"P�`0����0������S�<�ѩ���	�5N�4F��̥�n,�t�5�3d����~Fxt]�f�+�Tr�Ij^By�@T�!"+7�|U9?:��O�"x�vjꙬ�_Ͻy���z�����?����(;/������rfZ�H��Y�l;�N�����:wbM��4�q9EwP�Q�HU����9.�"V����깑��[�)
`q`��D:��>��o����S;v�t�T��D�2?|��~���I0Ԕ��w �t�-v⁓���U&O_f�RQW�ٳ|���[��E�ag9[��u~��s`VR�--0��޴��\Ɋ�����>Q4%�'�ga�)K��-�S_�uDU�e�	�-���D�]y������ �+��طpw��E�6���f�N���oO�Kz�Zd���`DT��"��q�L�)�X\�dw^
|�K꣔5;���|����":d{��9�b�G�ك���p�48c)�������H�yMW��H�}�ű=bǃ�,8wc��dT�7�_�dă�5f<�Bf�z�|o�!���7�1mƦ�U��1jM]bFI�8�%1U����N��PZ:��e4PsE��<�T)͉�(���jU�t�Or��~}s|ɤ�.����� �.Ր�l�>u��VB��|?�{�6!E�,
��"��g �ѭ�a��D���A����Ƞ�o���f'��b?{�B��vh�D�DI�&�=rZ��E1-�ۤW��) �N]#�ٟf��Guy8�TS�v*��DEYz2���\����ݰ8 S���͘�bc��y<�YN�E@����~4�"�[��G0�qH����P���}��fޜ���/����I��,��/@ro-��Ե���mB�a;WF��Lx/���E<�(���&�yW����L{��b�����rg�9Z��Q)&�Kv�����V�k8�&6[�K�/�O��4*
�6�Ɛ��[b��ӯǐ���p�u?��3��p��I4�ZO��E� ��J�7$!��X�Ý��@����"��~���䒜q:�6�f�2Mm�y%���?�`�8p�ѻ���~f�ߵ�����6S}2����fM��Wݵ&�\\�����
�YJh��&gDA.`%��P	]�+ԣ�|���K6�����UP�h�����ޑ�mEU9�C�<�M�#����êR'쌨�Kj@Ȣ1��L�(.2���[ǣ��,X�GN��鷁�������"W�I<����N�����}���\��ؔ�،�%���<����ʦ_6���{�F9k�j��b���� �D��ݝ�"�=���ړ!��F�[}I^�w��KRR[(�4�I-���6 8��'��-����䱤L޲��P��\Q��&��%)��iF<r�K��H,�ݴi	�BF�P��2�����jq$v i���S�n���1bp�"	g����eiC�Z1�e�1�Yr����Č}gqn����"m^Q��|���}ܕ�n�0	�@6!ᄅ�b��`wMk^�|�[�
WY�._C�j�Ȧ<��H�=�ER`������<�u��v��S�����h�*�z0ܛ�Ol�}��F�3	v��#�o��!�:\���ޮiLm{��i�pU{�{%�f_�W\@��*.DÈ�2u,�WM��~���}�@�r)���4T��E�7U��QT�_��I���n�k���#b�ˉOH��6ܲa�����N� ���Ģ�=;l�6ĉH��Á��t/$�m�XP�Z��]��ê >;5�S����SA��[���6���ł[N�!c���$*���/���kl+o|Zw&i���x)�*�4ę�n����]4i�B{�J��Y��{�}��a��Ei���=�w�վ W��>�7}y�`��:#EΪ��C�\ܚ.)YS��iV#��ѸӐZI���h<�CV�F�̀�c=R�d\���hd��l0b�4Q���g���'���Y"-z+��;�]s��G��=����(x��V��Iº]��G|�4;��V�MT�9��J��u����nO*����s����j�65.F����hY"���#^��3)���-h��7qt��\�������B�:>����O�U��=�}\g�%.�\��Tɕ�o$��e��r�>9����.(1
[��`��a�4�+�N��$��ұ6�9Bʖ�^��^�^��'cp��r���h=��j2g4o��׀��<F�2�*�Φ?d��G�}�[��p��!���$�2�>9�k��9FJ�j�o�f��UfC>ԕ�I4?P�ZA`�*�Z�r6�����;i�.�b�RV��5&e�
�N�V5��j�#���ߖ�Xח�/~{
}�RHE{��:�7�B�,��NGj�������S�9L.��@�;yM�E���|6��U3u�UZ��{r�݈7b��0�}��B@�}%C�ȝm��zנU��� ܗ_.�6���A�� 0禡|"hmw}��ƱE:��+�����(���*��2pE(��c�H��v�j�X-?d�<o���"�YO�HfRL|�s���
�<y;`<��&50�_�i�7{
%�E�l��~Z�T}��
mC-Q�k�j,��(��PR:e�;�pS)��_��P���ȩ����a�;M���5��T0`��NG���������w�n�`m��πς�R�K�y��Ӟ�+k��@�?�IT, -�k3�3�����!q�P��wWILeU��t�_�2�z\�{��	���$}��%���r��қb�i/x��L��_#�ŕ�oB́EZ�Ƽ���k�`z�Z�A�P� 6 �O�����:%�(�IA�Յ���p���o���z�5x�f���t��ߘ�����?���;�d�%���#&JX��@������h���dR�Z;R쭇^�z�T'�6H��@��h 4t�-�T��w�=]N9s�l^?��wy5�B�@_ܡ�䟅�u)HS<�ҥiS�]�mf�V�;�1|@�����Qd��H0@?⚵U���
	o�Io�;�L?n��{e9c�CEG�	���禡q�X��~$�����s��Qc��"ށK2�u��.�����QM��� �� h-4����9q�Q������DG�%�*��#\��	gC��4/��f>��+�����/��(�� }᫤���n��{�������~���%4���{��3��HPP-��q�1P�,W��5��%�T"0*�G]�:D⁢�"���6�qǄ�D�<��0�IJ-��e�qS����^K�#���'&K���o	�|F�>��IjN��9bk�o�nbt�C"�=4��u����mW�.���geeW�눙��w\�jG�<���޹�@�Mnn^�4�
sT8D�T����8uUv�E*+�/o=
�+>����(:��t"���u�x�Y��ɧ>�vs)g|U�Qo�k��縴sh�_�����kYr��sv=�wtl�0�C�Z��Ka��ԉl�Z�X�Dc�1�y��RTHg��u��x)%�$-Q�������}Ð\�$�H�D�8�Hn� �:f&�1�v��/�]P�y�=��)�=$G���"}���j�x����;�_�)7�rj�lͫ�Ǹ��r"�	�>S��˹��jWW�U��. }���SU���~�ObL:��v�'P�)���`V��YFω�d_8����3������&V��"��)%�̗����'^Nb������tO��NC+��점��n3��#z���=��e�(z�[� ƻ=ג��z���V�7��������_�����T�5t!:�A�4�L�xMB�M�Mɱ0�!�{�LZ�"�"�
�X��+�t�yR��0G-��AD�!�۸�ݛv�>���>ڞ�Eҧm\�n���4܅��jѭ�->�)¸I�����	���u;���A���0��c:�û�G3m�u�ĳT�)l3d�4��>,�
:�!7���ft�������`�ou)����ɣ�Zk� nf������b*m����gL׫�V�`Z�ݢ��v�P�w� �±���La�6���7��H��EFn����g���a�[�sf����w$ܩ*�5zdV��Hm
���许�����ROx2�{1���\J��~�R������ʜD�źZ�h�5�!S�Ƣ�Q�~���M[�ni�Ot|Ml�ni5���(h��zӄ����^2cw���ƖP$|q�n�����#j����x(�[�_X��^�����ڦ���^��5�����4n)�2è��r5��'�I����6x7���!��\e���g�E OB_�~��+gb@���X���T��H���Ѧ��V�l�;?��~��0��I�8`_?���[~��Yzn���y#q�s�,^<�|�$���8l#�F�7*f�����u
/X���Z�9J�/����|~r,��u��!~�:�A 0��z=#,��)Oeͬ�����Q`���Q�EZ����]�Y?���4�@� ���"/�/�˹��$,��6�"�V��#Z��-kE��ft=��wx�/�fBO�����K�-��Y�ͭ˒�^��ĩ���� �.��:��y�͎+���Ԁ�`n
J�,��X9,�K@j���8��K���k�5T�ʾ�����GI� �A�uO���^��:�*ߤbڿ�u��;᜴�}��D��)��u�,�`�k���a�o�C��ab!�b����7���yڼ�cg�p��bn_rP�gOJo+��声q�-ϸw�A˸��ʸ�e���eV��1`!���ޜ!�0���P�5W�<6�V/;�|^�~`@�ep�*!,I�Q�(��5��&�7�.��K�zk����_�n1��*�e7��r�7��,�bJ`e�GQ�N���_9�}�������B�^��G&Vy�V���22ap��5(�?���8�e��יѫ�=�23P�3,�Jp���|/�)��0�bl�+lcX�[����77&�@��'_�ۋ��5�;���>�v��[�)#�C�섾q�����Zu��)Ay%z���7��*2c\_�����0�>�� I�T����E�t�g�|����U���P#�Ik�M�97����	HsB��*�b�NJS���8ٶ ׭�d��il���[0,��b�D%���͖5�w�NV�хRޙnA!%��8� _�$�!4�'[�� Kd�-�� � ��[��C��E�� ��0�#/b]�_�4:te�?팍t����o��9Z�����s���fy�Q^�]��fX���\@&&yc����,[O	{�N=a	�^a��]Q���F��Lz:����W���QZ��£�v�gȞ4mg��϶o�T���/�Cz��M���-|Q�P6Ry͡b�:v��R��n8I;F�0^�@W�����`�;[M�+�mr�6Ue�k��.?��i�F�B�TAx�P-�5On�U�@����,�=�-&��|%Yo�2T8����Q|4�Ѡv�ﴙ̔��'G�q��Y�Gl��#�!���]���\�L=A��siv�_��w��+�>㨋W+ ��P�v�G�N��yz<���뽱o�K:�y�(?)­��?���>��h+�!!���,g����e����4���/��
*,bc�H_7<�b����T�����3T���M�Ӝ�^��lK�+�P�3k
*��J{��2M h�w��17��|j�D͏�W.�[��Ȝ+c�.z�t����7�xX��?Z��}�҆.�Z���<�/�̭��Z���G�J,Ώ����D ���h.B���o��4vp@WW�W��أ�����������h�}Һ�桼Z*�\o��l]�(I�>!����FSuz����Ͽ�Բ}�D��L����DjG|�UV���
���xv[��9�B?��t� �]��u�`�v���<N3������=�yh;c��H����ow?�H3k7�~�Ks���8G����s��خfk�ğS_G,3��%p`�ε��f[��o�v������qY�B�y������[P�}7xӞ������'�5o���G�7ˮB�u�jg�1F~�u`�W��ώa���5(�p:���Va$�C�o�V����q��Z���� �g~��҂�&0���l׌l��%37E�Db��T4�@�B�#d	��	��Y~3S&R��"A���h��tltDD�:�^2�$���v�V0�X��\Ч�f=��&�ó��SN#����E~FC����<��0ͭ�\� ��}(!돵�:D��i,��~�m�7��i�)ӗ]����.z���w�QU������s��=(�YfW�vB%�0�(��4#��3�`�lM�1�b�e�w{n@ �EG����"��2�m��{u�B&��<[c�i�5��@�B�[66z>�m��x���Vh',�\(m� fZ�h�@�!���[<�zQiŭ.J��3��d$RgXK�i��#�ٷt�l�8�|��2��#�]c��]�4^���<I8A�	-y箛}*���q7�������κ{��*8�<��34���H.(Dg�˓�'B{R]�L &>/4�c���,.<kf�3���}lhD5,�˙�G���'f��'̶o��kI� �{ZKTg-х�I�.���M����^W��@�˔D�>�D��(l�I�J\��z�9m2����ͥ��^���^>;O���M��Ov���$��|���� ����������$u�E_4�ՃJ��Є{G�r4X������&���Jk��X���j�Z�`��8���X2{Q^j�	�oe�<h�)�:&�P6���{+�N�o�Dqʙy�����R(q��B�p�}T�tӐېt�!+�%�bL� �)<���S&.�ay{0fv�M�+K�@��Ȝ���9 M��An�`�e%O��4΍��n1\����Y��"<�Sx`���2�ؖ�FF#�`x���e܆�����-�r�]��t u(r�"Of�f��31�G0�0��@E
g��	5�NB����N�=�����CVr�3���D�O�ߛ�%^���N�Bw0I�S#1έ����ϔA'{b���eKw�]��f�F��OQba��AS�_�E��v��0]ڃ�t���!�îƤ�|j���>����F[�;,i#���F���QTE������`%������g��b�8'3q��e��l��Ա�̑r�8�yqX[���D��.�h��˅��өq� ����x�%���.�;�Խo:��9tJ�������PX�6JCd�4�;�~,������A�eo���{/X��ZvjFqj=��{-Dӯw�i{L�'�h�My��jPk5�4��Z�0���H܌`?�U��>x�kV��q�^�dmg�q0���T�p,��S�m�z�Bm�%X?�$��E,�f���vC=p����U���1%[N�g�S�������*����g`ˬ�*�	�b�M'οu���6��g�;���������� � �ݜܳ��&��t�ʼ����I8�(l|�yL��aQ����c��Z�U�5U��*�y%�b�=�$��N��{��$�XX�g���T��HB;'x��_)�rV�x�;8"����[��|��:�ߏ�np��bL��|�;u����3�F���R�?������ו�b;.���S�Xk-Ri��@)G�;�f,�+������bP<�
ׂ�@�������A�
��3�k���6�����_�_��r�5�9��)�is��e�ݫ��eڭ_l�-��ZV����L �s^ {��RT�jD�u���ï�#Vd�e�E�i�)xq8�������v���
��mC%�h��)Ǡ}�ZK͘��C^=9��IB��^��W����$�t�_QU3	����D���A�ٵmW7�"ǹIi%^��b��(Ҿ��VO,��c��i�-�Ѹi�7����p��E�џ?�|h��x�O�W�e�O�;��~ O0F�4�� W�{�1#��,9p�>��L�4��@����FR�a8$ �u>`\�־&u� Z����.��'�����1->C�v�,J�fygp'���N�m%��w�]�0/B�<���v©��6&��'ߖ��Qm(N|3��o����7|c@}K���AĄL�/0G�M�&��e����V�az4:5�?׭:�Y#o�����)j��]���4|m-�C'�:WsEU�v���%!�?�v^�-b3+�A4���:6{�S[��x^4e�4�^�2E�6���6(OfI'��c��/�����I�;��3Ԝ�!S������۬����z�p�:�U�4M��Ƅb�Ň�V���<h���6��Rx���o���h��[������,s*�6����ir�\Q�G��;u���"\$n����3����=e�)M�Qx:[v�>;a|I�|:�s��~_?ʥ�����x��Hs<�;4����؂];���.3M+h#�}�V�ֽbX������ͥ7�c�\d��;����@p�+y��fpn�[�'t�.ݩ	3�ReoG��D��(xش��=�&��cj���5�ݘG1y�[��<X��4ho�*��|,�Ȁ�p���C}�'���Bs[��1=|.A�W|+h'/{�뿉ת�9�6fy��ţȍM�>��O2Ktc�ҥ�@ ()#�ẖ���5���; }nX��Z�a��T*{�}Ή�- �ԎOS�����դYϠ*�\�+�4'�?����Q.c�RY��V����b֪z�P�C�,9�u�Q�	�AM��� ���*60@���qL��^��������TUk�t?��j�Q�tK@p�����%�.!��T(��TL0ŧ���kN��j��E�׎�|\\_kHK50���Oii6m���!Ĕϒc�7j���m];�o��z��Lg+#`;�dN��J��|���6d��؍n�x�2G�%G�w��3�4ZR~d�y4RAe'�}��vj35\�n�CЏ��J��X�mqU)"-h?f��TZ�	�j���FQ��pMU5(� N~VZ]Ljd	�GQy"�P#0egc�𣸽��?�cC�v(�C���:��-��Z��C<;>�^��gv���������G`?>;�.�D)rxE��-�d�Ps��4F�:�,���"�ߣ��هv�����&�^�c&+E�nC��#�3#s�E��?�rCS��5m>��#���M���63��W6�FgH8�/`RB. ��ğ+��=zqX��aO���I�]L�M���s��}�$ub�v�l���;�Ǜkԝ$ˏ�t�)K��܁j���s���E��&��w����7�\)��~e^aJ�Ob&j����J˛�Me�q+\"J���깶v���I�Sr��Er*l�&�X�OY�w�Q�` i%&a��;���[Ț��,:��gx,���w�u�\��K�o�;3ڌ*�	��q�� �˃�a��z3VKK|���"��=i�ʫZ���Z��l�������$D��9�*�Ӄ	�oN�Z5���R,�����і-���J���0���i�e�_���E�C v��'��ė}��S�C�Ϡn~7gbcS���c�b��	��} ^tk�n�7m
xT�H�Mҏ�S٦t�Gr�~��ME<�KSJ�$G60yW-���:���B��}��sh�&P_�E�[�l�{�_M�(�l�r�e}��K?ʤUJ��v��t~�#��1��KI䊜���<1+�qҺ��9o~U�G������K�%�h�7���Ԩ'"�O
�)��]��d8=!��� *~54�4�wu���8!K�W��0�����4�Z�s�����/��n+�W���yL����*�/Y�B�S@ī��J�c?���۟���O�j �D��!���'��Gdh+�4:7?|̖�=���r-s!W�� ����>\ɓ����ٴ�������kb�K(gk�F,���Y6���qc{����bƬ��Ts�"�q����TaN�ॉ�=މ�p�?Y��ep`dx�
��5�f*m��}�M?�����&s����q㥶X��?�O�N��̯]�6�[���Jn��5��l��`=G��j>��*���{q��_�a�������(�B_R���F*�o�K�h"�5X�*uz���>��(<��K�G�E��b�~��*X]�wv�Im���l;H�����6�W���A�3Ӗ)�k�Gy�k/�]"�NlQ���y������]y�5�uXh;!瀀>v���;�79�Q;f ���������X�7-�9��p��ɚy������-�U0w��������,�H��kB=t���18R�Wb"@�^�p� ������`�<"�)��ٞ��5&��}H�vPu���e����6����~]�EYj�>h�y��W�wL�%R�ߗ7U��; i͜s����ȱ3O"��%)g&re�wG
�A���m�4b�ɗ�A�����R��'T�����E��ǐ#��߾'�{tS�%4;jw{e�Е��<{�Wzk�}���+��lz�e����Xi��i^M:�j�|1�7T'!ߕc��zA�I3h)�g���Ij,-�X�B|{��'�G*��˶,_�}жZI�{	>��;�e�u;����[}m���e&;�'����fy�����+k����M`��6��IR���"L���]m�/2��s���(��y�'�6s$��Q3���Ћä$j
�::\�b�udʄʐ'l��p�&a�Ҽ�ť�|�&� ��B	���cҽ[UɅ���9>��aZ�̰�4����'eK^�!L'kC1b:;�3�'����ڳn�� ��_��b��h�S{F�(�T��s��ޛ*Xt����W�],��	���h�o-�,�Yg�c����i����-���N����0�!���V,�-hّTڨ���K��O��8�:��e�J	�*�zFe�=ȵb�aX<�Ǭ��4��{���CG��-왋c�T��k?��8�[�$��2�@&��3��NXvd8���mr�+�y6���ʙpd�܃�]\I�\�{{��CbMD��p��MI�X;Ê+����2s��!8�D����Oɽ�z��ʃ��!@�:�&/���`�_��E��U)ٳ*�_��+���&h�7}Yn�w����;�y΍:\�+|���9s[;��U��Q���)������J_$5�5�N�����ԯ��@��ٱ�7��)�Ug��uć�����
��5�Ұȯ�XTEAK9�O4C�F؂�M��!��|�k���4ܸ�DVC&>)2הx��4�@���!����f�,��u�tKYbEL�K��ϔF ɤ=)��W  g�X�Xz��F�����9���>�]�V�L�E���C�#��-�J�ȱ�f���o#��oY������pNHkn�z�>��Z���;g"�����$��o�����~�>��.\���ݬx�MP0�̨
4K����7R�h�) ��.��8�?�T²��'Y��Ѡ�5�e�w;�j�}ܿ����Y����2A��udx"2Gw���0aO5J(��"���/-nP�K���vf^��c	n�mYQ�%�3ͤ�x^
ˉɻ�	�8"'�Z+>vU�E����� �v�(y�΂	��H�Be�̵q�|H��~Y;v��w!��߯�R7�HQ�Y�-����.������\���_Ka�ٙ��d�zh���",�i�ge��V؞�#�='J����`O-���\�tiR��sFA��_o>?�$ҕ���F���,1�r�A�q�&cr� ��&!~c�����/2tan,��]q�����ړ��!�H�0���������dUzΎ��o-su�"(܈9�-�!�_$~y���YF��ˣ�1c�Յy/�.�Rd2W��6�j����0L��8/|�z��k�l�M�Ȕ�*�S ���v�ϛ���i�*�X�1���mZ�����3i�^�g/6��w��Vi��se9��t�%�m�8P��>���_-3�o�+--Ut����<1aD�����E�^��Ij0�>g���l3��`i,`������&Ou5qO���Bq�CAD��9�$r6;�{�n8I+��'^����"}���❉#�6���4'�����w�ق���� -<9��i�R�ۻ�=�m�p̉�������X5��zA jR��h~p~�r�M�JĒZ���I+�e�m1Yԁ��7�]w���M%�����d�~���&� ݇���u���|=��Z�1(ny��bبk	�_ /.�vH!�'�@d�h�IO���2Ww5Q�sϰ��jt���Y���*���3���)�����C�ƅ�� ,�$:W���E��][�}���F��;SΓ�Qi�6j�?�#>����]��52���t׶A�T�h��Y)Z�Ekև�\�,�n����w�'�e��������pU�),�m�XX?�&��wY�\����w��V!�s�Ƕ,N�hذ^&�Jx�ȹ��d ���%�F�?s<��WXM��MaR��;��a��j��a��1�C�T!<t�&�Q�Ƭ+�y�e���f�)[C�h40ОH��֐��@�i�ǧ���1e�&Ȼ+&!t�$"Q�q�p��ڵHkgQZ�X�%�׫����,�JB��PS52��K���P?3?��a�<�%}^5X���Hs~�&�7�����9�Y�}�2�e�*��JޝH}?��/����s;��gH^@.Д���5�3�q�{�i�'����0J*����l5�Ka���t]�AC�8�i��VmRq��!5��aڅ=���?3Aī{�Z�����eCy�v��󼵛��i�̵Wv-�T@sj����x�ͬ�o@� KȚ�f.����B�y�YQ}�y �?��ی�+۫�W�)�$��N�[*��d=���~{��h�l�X�Ч�X�}r��u虂t���寮`UY,۱`���_9)��'{���ḳ�.m�c�]�`�m�|ժ�m�Ū[s���	%
���iVm��8|E��n�*��h��s¢
39���k��<�/͡勴����������x7O���4ie��'$M~�����)d<��Ot��c�LO����l�x	����Έ��[��n�e�y�&�6>�h���2�
;\�,+�M���M�«�T=�:�Qj|Nm��=|JKZ�+�c�
-pj���Iu�P��Hp�4�[�<;?PU^��q��V�>�n�9ߐ*���pyTh��b�����n's�C�L_�"�&��qyJ��Y��x�ŋ7x����U����JV8�$R��^q��X���a2��)"��\SW�C}ZLxw���ޫӂet4D�y�e�B��d@EXm�.ï�5��F)H��)���7�.EȚiiSxs��G(*�F�p����}�l�%��Z���:��q#�R��%�;�2,i�<|##	+n��6�v�����T��N��K@�Ňo�}3-y=h�J���yk�30�atv!c߇η�p�����yQ�.d�K=�����EW@�T���x��i�~�Db�G�����KL�[i�$���D��`����W�������($E�.b��c3K������E��0�2-7� �:�.H
���Ť?��jY�� �Zh�����d�}�m���['�m^������d?�Y�I#J�5>���{��_�nQ�(��մ��:��^GB!`6��m^�9�
�ۄ�%����#@�۔z�����Xk�>��ت�ʞ��*Z���^M���̈*���`����<Ǣ�L3�����HxM�q�6s4�X���V����M�	 ~��K��q�δr$�8����/��(�ai���<<�"��>��AR7
����pD��C�\[q ��R9�6ZTGB;FE�����!Z*�~V�u�A����GX��\RNP]Ӳ8�'�3m.}fS��ذg8���F��(rF>��\���<Xx&	���L�����j�����f�ڭ�FBѶ��'V�
n=�M�n����������Y���P����ו�5D����8������IO�a�S�,~̵�,eD�g�d�A��V�'%r�(<Y���#˫V���XJ�:���:���ݗ̝�5zv%{r�N@n۵�+�[5	"�vG߆'��������b���b�.-�ae�z�t�]�i-���j��υZN��2��	�E&�mNH��2un�(��)�j��#/v��ƨ~;����;rƞ��P�
�!;x>`m
�(g��xh��Hڳ��)��J�%_=i��������4��̡PY�o��Y	tߙ�ἔ	�ه�:!Q�y͈�"��;"���rI�D ���4�U�#����.��<���&]Ǧ���w�x�9	�:t��+����/	N͆ ����������'��¼E�?|Ù�t���@
�C���KUYt�0g����ӫ�����nC�����ĠT0�ҋ^�o9�N�`���£��^�Ԫ���b�i��$k�Y����ĭ�:b� ?�nP���o����#!���������ch7�`_�:�,��`ՁJ��[�T������"�����Ә4�y�(�	-\�
���/��'�Q6K&�J�����oY��L^b�W�%z�-XS�~��F�8eii�'�)�*Fۖ�� ��E
/	9<�>gU�מ3ea��`��Ҭl���*�.)[4WU3���)���"�{Y/_(}�C^�_���
g���ms����ᛰ�B���^�1x�Ro�N.q�[W_itt+��]7*Lg`b�)���JǤ}��W�zSwۂE����@��8JS������F�R_Y(����r��I����h��x����8�(3:�2Ŀ6�����וY4�GJL)D�5�j��C���rưwE<�8ȦB@l3��\_R���Ex������B�}��5�H'J��&���68)����֡��~ͼ�����OI[�IOi���|�"�S�z��z��sp�TSV�����s���'G���u�����D	�<������!c�؁�����
�2��%NO ��م��� c��̨�O��ꊨ�Ʌ��w�r_�����@?%��$���;��g���j���5�:T�3�©��Ɗ��1�q�C<O\ލ��i�� <gb�DO�O�K}|�4��ֱ��Y�B�M���I�7V�A*��qk����<�&�[�|d�y���J��j.^�PH|ۋ(�iP�<���UTm^�TU��g��S�M�j�M7\�T�J�?±��5`��3?�.4�/��ZO� '��D��*��������N��3�D�W��c�ڽ�+'�tX�l�pG$((�K/�v�\S��7��Gv��Q[��DmWѮcU�_�M�(����V�Fp�Pԏ�E>�$=<#V��#�I�k��%W����E��tz\��`�aP�BМ�?�h�X�8��=�<!�3מ����w�y�-9��n���kE�6[�%�S�p@"� ���(-N�e^_Vg����DPøbn�zUx%�_(�Hi�K����	g^Eφ1���s�u%H�Q3_�������}��?P���1��ko���^��@��0j^5��CA�x\��,�4U�
(���i���8$��c k�.�u	R��{L����&ob4��X���0`�/-R���]��ƫ�"�=���<�vO���u���`C��)���s�ӗ���+���x8�?�!�����:�[��d��1,���a�	I��4�E��
u���<�FuJ9����*MC�g�.ja�w�Y��g�-R�V�8�\1�=(ֻ������G���F��U*�����f���3L�%���z�\a����z�N���)+��*�~��n�a	��Ք[cq�<�=�F��D`����bZ�xK}�G ��[Չ��nԎ4E�f$(����ߓ��.w�$<i�W"��>����lXe4\�0��J, �����t�_�Ko�9�����O���)�0XZ��g2�i=kז�g6}��G�03�đv��aY �sS�z8��qؑ�e_0���gӾ;��]���E��P@��U��גߧ���<�w�O�$^�p�
�B ��[yZ7+�j�)�N���H� �mCa*s�
�}f_%u�f�U�	��++������m}rR����p9*ET9fF�GӔ��Jr.���dE'ho���/m��N����t���hi�N���~��[���<!i�}�4��KZ29��&��&�4�33�Ggf���~��������秮��-9��;rZ������e��]�?���i��X3�'~,�oc�*� �t�%��hՅ�ƚ9@�b�b>H�z=��(�<y=l��m��(�*cY����[G�d�s�5=h�`jJ�=h�CH�4�h�G_R'�*T?��H�a�<f~B�&Zкe���/R�-�&,����uVޑ�/�Yxd�'^|(��-�)O��\84�:NPI=�7�=묪+���}�̩����l��0
~k�Y:��_�Z��q����0n��?x�U�5���٦\-ư�@�̳���z־ݎy,�5�l
[��W@+��h�N��-�2%\��6��K]G�Y���|��+B����?2�/�`�I�]���^~�RϿ�ν_T��2X~x0X���� F��E˞7*⩴LK���mVr��S�K�ơ�T��kЊ���X�͡�DNl����$t%��6�~V�����Ӳ	M�{�0�`"Y�wB.�]f�(��^�@�K�j$(���W�Y�������Mxy0�r��������gr�ms�ȷ��pJ{��l��;����пL�߃�o�h#N
�} ��� ��TZ�:�L`�Y�9�H)�qְ���8��jZ�Z�����k��-|����v\�L�n7��݉p6�o%� ǽ�@�Z���(~���(������Vb�F��z�����&�1"�Ƅmh�u��ג�;�OE�!4�bV�*8+u"�g~ƃ��9J֫�$1c���Ւ�C�����௭Z��a��p�&i������϶Y0��7T?�9���S��G�
�1�'W���h�������[��_�8�յt���uz��m�����fd�}�������Y��==5��0G,f�`�j�d�;ّ�v~Ô�*��V�\�/��}Ѕ	�*��X[p�l���.�g8k��[�~߼�j4�"����M�p6���l�u���r�9iUa,~��K:4sX�m7Y��t�2)���r���ҧ`��)��<1�h{�YD@[��&�F��EKA�0ko�k:�[w��7���> ����Ɯ���9�vY�S	��Z0	Y720�%�e#XZ�(ރ[�{��� ��i�@��"?
'��ez���_GD݃5;.wa���+���d���P�����e��>PQ�X�#_J�G�].>���꿼ޟ�߽D��x|Η��K`��4;')�8mΧpN\q��I�J93<��R��}�+vǫ)|O¦��[�����o�Q�mꯩ�ˎh��	k@��ƸϘbR�gYT-Ã��bn�ÀG���f���DӬ��o��*p���qZ���f(�O'~Y|�)'Ƅ��/�*BA�
О4�Z���2�]�zMtf7�M�K3o	�w�|���4��HS�"#k0�B�>�Y��ɦ�����z��e<��8_�� ���)vɀ�YV:���F����a�?ѵhFy��C�y<��.$>�
7  d�q�[�$h�ϼt�0/$������G���E?�8)iq�_��jc���h�ω�]v��_��|�UQ�{��X��N�=y�̭`,P�U�CQfе��&����IJ��gC��g��|�f�<9�B��bo׬/K	{�i��nR����D�"�@�ȱ��M�hdV[
ț�)���'�	}>P���!9<LZL��K���O�?׫+�3��v.��i9M�5��,'L�=Rgt��l~�����'�i: �'?�z;��֔-�y�cW1��%�E��p%z�g�9LJ��< �=_�NY�/�
�#�V���'��������rX���-�^��
a[�U�m�b���l��?���w�������&���y�ch�J��#B�P��ӘN/J���\,�TcQc
?v�y%򞎊�4?n�+p���5|	N-�k@r�3��� � �a+�5C�oHnf��h�v�V4�������l�7j��Oϳ��
5o��[���9��G�C��qW��81V���#CcB�@��ԃQ��r�bVWA��1P���J@�t&�lX)����EYwȏ���ELȈ��Nb�HWX�%5�C��֝G�홾��ۘ����>D�{d;s����c��,����<��	���.B�۟�W�F�b��Ƶ#�uQ�&�|;�D4ß�ؤ�kw��I��[��a�&������Jd���!�>@*>d�$��e�����%��1�7�x�m�ŋ�U/ �´oɂ��B���i.��;�}�Gd�l8^������ܮ]�-A��vT��ګ��1<��J�8���A6�}'��!R������2D�D���Ƿ�*�X�i4�|g��&�
�#��a��Bry����ߠ�-Y�,W��t���e���4@��&�ٱ0_�鳚�5�������>��u�PP+�� a��4,�1�T�����q��= �FU�EJ�w��6��Te?$��R$<:�&JY��;�n4���q��CX��.dRN�&�Q�d�ՙDf�_�A h����-w�	]jF��354��W�Sm9�����<�O��-%M���� E��]!�:<�B�%�S�5g�N�"�IH�j�F����U��i2���bq�v�ri_,�h�*y��������P�)�F�UFp�)i�=l%�'\.#��r8����Y$EB�ŋ���$�N���5�Gm૘���Jf��J�=ĺx��"!`R��%��-C�Tj���5~n�К�%6��.5)�Ԛ��k5���Ͻ>�)�0�>`�e��xG����g�&���M���T�;T�#32)���z��EJ�Dv��s�>�3�u$�G��Hu�bKϑRr��0���_9r���}���u$���7�P��2���ji`���(^y���,=p��G�q7��WH��jt�1i�D�.�XKT�*�$t1s�(�@JL�,�@����'dP��S�b�jo" ��C�2�����r���4h�}}(�<��>����f��3P�\/��k�4.������+��;"N=�\��7�����2G����"�6�)�֮��G^K,��v���ߩ{�~�8�r]��,Ow���f	9�R�J�Lx| �Ӳ��G���15����]S�[3�-0]�<����k֚A�j�C[U��rd+��>�U��zox��7`��J!�.���I0d$S�%7o�2rl{���L��8�K^i�<���	I6�;�VsT���	w O<�J�-0���	�hP-Rx\���e�Dj�~ځ��}/�:F�5��D��G\S3��Ԧ`3x���6"Y�d Z\'�������,��9��~�M���19���ݫz��D/�r��J��ā�w���@e<����'�KJ����<d�����9��ފ� �����͸�U����D�>؆Ր~7��*�IrL��J����o�08~S�'%�U[��q�%P�<�����Y�(L ��H��(��7�B�(���z�R���� �و�0�����W��۲�m�d�Pa1�)�^A��C��&a�ad�62��x�C������h����#��{]�?=���o� b�oS1�{�O���+�y�3E���vI[
W!�3/�Iou-	ѳ{KE�8��/I�1ԏ�(�_@����n@5��x8�ȍl��R@�fS��mӌ���[�[�(鉨��Jv��HW�Y��Ƀ�s̐R��-���J(�cN��O��B���S�BO�����hV&��!��2���p��		P�x��)��ι� kF/+�"���k~���.�� 8Ѿҋ)է�/2$����ixMb��E����5-o����arٟl�*"�Ch�TY��̆�n,d&b���ÿ&a�mq>_����+8f8> G6y�m� ���#lx���P2�ǬZ���Σ��N�ea\��_��!���%6ȤR����L�p��^��"�t�*�_w�8d#��"y�.� ���5�vE�" gկ���F\�*�/Co��p��h��C
�I/'3��c�樼�>>�(��X�1�-~<�l?���
&c$Ӊ�h�9���>��(g�toD"��M�s�h�C�ȿᩉ]��� ��|U�Il��B=�8��
r���]��Ӷa������E4�%�{�Y-'O?���i<(T�?��=p�J̯>��_�0�#_�<������d3RA�������{4�oR�߳%M�ƁXz���|��!��mXV֥�$�;ڢ�e"sXt��ʭQ�l]~�H�������h����)�с���HSܽ9��&��㍇����w����˹dmk8���h]_j����CD���&�aJ�1l_<*��Z�_ْà��=�a�/2�*d��� ��ST��xR_���Y���	i�X��� ���L�SJ[o�KQ_�Q�W�+�+��]��x�Ɛ��uE�G�g6�I_�<{���N��q(���7p ݱq�L��\؋�g����z�_7r���-/e-�ļ>��Ё�Ï��Z�N�~��;�5�"HΕZ�?�NC� -
&�]fD�G%^R�x}��F�O9��KY��Y�펃��z�=_<�~��a��0i��r��S�?�v��y�~�M!Ь".MM|��݌,9�����w5� ���(Td��8��+$v͇bfg����w�?���<˰�1rԋ	���z�����P�p����G��W����>@T<V!��V�g�/��|�F(����.�&��,.��4גK���I��
iߨ�/R�U�J02f�O�8h2�iF�ܪF��q��ŏ�5�M[�jfp,W���0���A�D��XS\Y���k����s{���긯�dŽ��}�Z��gA�r�W�c�D�|��)�{.�&&��Dˋ�f�����;�&HϨ���C5���^�R���H��r��w��-�N[���R�ko�jQx�-J-K�<t�ð'b��c����fbE�UB
�lcx�O6 ު<�u��|���"��Q$�����V��xCNj�A@Q@.2F���Ư
�Y+^a�޹hBC<�v`�f�i�.=�e���u����
��6��!�\���I��^�`l
*Bi!QΆ# Q�#�~]���� �m�I�T�WB�XCQ�'�ј���5�Kq���O�\PA�؆.)�js9��FY�RK�GK�奰���Sx�I�&����f��m�c'�.���\� 1�K!AS�������e�x�����t3����#��@���J49�R~��W.�ڹ��w��)��p������Ad	�1 8
���qѼ릇�$�M�����@Ą[nC�+`Q���
�Fͳ���7����'����%䭊�r�!�e=JU秐��������E�2�J����y�sL�oɩ�i2U|����j���he!�s���pbr��0	1�{n �/:�`[�M��}J2�����@,K{���3�-v���sH	z���Ҧž�i(���C�,�� |�w��q6-,O!���dd��{�3)���3��
1���_��c�1�<t�T�662���_П\^�9t��2�!Y�����UiUtفh)����m\*���_f��i_��4�	|��:�����	��T��[�rz��X��Dv��Ǣ ߟ�]����+*0�#�)@��eAxE��wB����N�{C0(�A=�T�}_TnM��)���M��A��b��.).0�D m��=��.�)0��l UۨLt�5�_��[��e�^Ύù�S<8|x�p�����uWo���
&�t�ȵe_�C*����o��)�)��p�y~�CE�Mb��MXC�sf0�9:�\�5!�	--�[�{.�t�O>N��R&t-49���tnKb�1\$�uX����[�h��">1%�|��
�qY��3۲5���Q�� �=��@% �p>n[�jJ1o�#Рm������ջk�@
�<CR�4/��c(�bF��������/���a�J(�� N�� Xi)���ڶ���i@�j>@���6GSP9�9kSx�@� �{�X�(�ߐ[����.�,LhJ6{@n�K��'�:�Dc/�=���_-V�oSxu������s^j��j��1��W���W����o	}M9jqʃ�{8��E���}�6�g1�-�@�u���'��R�t%�i�=� &�Q}
4i��5dG���_��ӥ���;xB艃q��d�X-�B�Ps*�	�N�}��S�"���f�R�]; -���֠*D��FIfO�r��ſ���DI2�(Vj�Ŀ�JQ@�J�`�7b�1/ݧ�a�&�!	]��\m$x܏�=�.��GP��8BTF��%q3Cj�����xy��W�����Kmψ���Е���k՞���ظ�-`��l���"����@�����_��3cF��4�yI����ۋ�!�S��(IF�2�����*#~*��i]����_���=�0l	���l��v�#=B���tI�V�J1\�u\��z�O�$��e��/C�����7���Z��{��r�Et&����?�Chi���"c�R:�v;���\S.���y�/������`�/U1ݭ�glE��D�im+Do���iH��I�{�a���wUΑ���^���i�8<� ��Mɏ)+�#�����H��5�{+g/V��g�,��E�d��EN�C�h�,�6�&��c8�Sƿ�3��*�rt(��d��N�F�Ο�Quk/�������kb3<1��V����L ��x�;?�KU(E�����	�d��d��bɱ�P�Yֶm���	כsF{������dC����H���O)2S�l�O��Zo�C$C����v�<������A��b��V��վw񊛴��/�3d0|��!�61#���ʔ��a��8���vb	�G4�7����&��k�'!q-'|�^\�@ëD����t����M�=���r�����j~�N�����sPjq�L�Fu��$RI��^��9+8O���ov4��h�+d�'�i�"%�Bjn��4-"�vJ��*�uTɼ�Sp�x���u��z)���Y�1�
c���0@l�$sܓ,��������ѴeY2�#[6�N;~��/t�=#�{h�|'`����&����kˡ���LLNc�Hԕ6�nY�Ψ#Z��7���zu!���;���[\n�\�|��`W�ym�;�%s�k#��hU.�� �amT������{��>r�VB؏⛫�$��mX����q,td7���k�.eY�k	Ao��6����R[a�Z�4�����睿�מ
����V?d��v��V������OE7�n��P�D�I��w�Ϋ����T�;�UCh��}:vA�J�J'm�Y�焮4�,;�=s�62��P��9:Ik�c�x�;ӭ��΃O;�Y�@��'GAU���,����釾���SnKL�%�Ե��r���%��J#���L�RD]��^{��z��u��g]!��]0�q��� 2^׋=��������Lr���6�^�d������`Q�C��b��֭�� @�8�0��}`�:^i��ؗ�8�k,��|�V�<�$��v��K&d��[ CJ7�B�?c�ò��Z���(N���GL�Q���"�R��8�An�?��da��R䄧IZ��y�e�@���-�B�厜��y0�(�B�t�-P��O��˼K�p�C���Mʐ�ݝ��y����ή��m�i��V��F���Jh�7����F�Y�Y���S�&�z'���]��tj(��_MU��w&nٻ��� )Z�\�;ܰ��JK�6E����uۼ=,"{>[�l�A�����T�yY`2!	�`F��3��N�b	.wq��YL�Pm�����@g���9� �\�9igl�� �,�Zn�� �ǿ����fz>�|�K���p�˦Q�I�L�w� �����a�3�R]����������1=n6�H��J�ƹ�?�
UY�,��q,r�:�)����ro5E�7c�cS�+Qu�{5�6��g0����7ז&x�7��n��cy��m�u��w*��<�n�ܠ��\z;&�4)�W6��V�b��'`O�����-�,�VoEN�/�#fM-��4�A�f�ُ� �gm�ߚ�R�?�?���<�5O���8l�l4�����q��ٜth#�����堵V� xF�]���O)6�e��
i�z��C	BB���ն�lw�}�6�㕥a�
 �4�,���VE�]��!˱�۫�"�J�=����e�1Ē�
�=yq�uD�&�>@��x��+�4&s�֞Qd��8��� L7ʎ�J�Ӎ��t ��E����#��RZgm�Y=Q��)<���bX����܁��6R@A�#Ѭ~���;��w!qجLN?��E���P}�j��q�P[��<V����`��?�[]^D�g��y���3�;�g�f38jR� w�!TC=��yED���W���VO������IMAX�C�P�u4Ob8$M����Y�-y[��c���y�4���C�c}Ad�w#��@�q��ث�W ��ي��q�1�Ba�8�7��ъ�M��nBa�� �=1Ӈ[BԲ��#����L_��K �����\����?�k��	�cj0=�)��I�픏��&+� a"�L�ϓuUJ�!e��.+���q/��x,�`�lp`��t���]hi�'M/��c�J��v%�v��@�Ud�F�Xh
���i��l
�yu��s�
l 9�2���&t4�h�1}����`�]Х��M�_!'�[����99�6	RN�[|0�X�d��_xSU�'�
D$�W�JH�����'�-��i58/ԩ��ɜrh����!�TV"����#U��&p1`�?����:��a8�U�"m0�[�J�|�m��}u^kwi֧C��b�b�m�Xs�:��ĳ��C�L�A�XmPi����}J�-mT#9�պw>Ā�r~V����*��%W;E�jC�Ȇ2[����9=ݖq�݇�7Q�h �C|b���>�d��F��P⌽�bb��I�w���'A����4V��A*8믷R��R�J�t�"]~d[�sn
��']c"���Ӣ��j��=7.���=p.��H�܈����Z[��UY�]{!*PS�20��-�D��'Ɖ/I�=�h��2iM�Q��C�m��ـ�cDbc��bt6�9�Y��w��ߐ3��<��ݵ��?�'��p6�;��H��SU՛D��
��7e���6�+�J"/�>槿��^�ҝ�0�R���`�pQ2��B5]��3�en��0=Ʃ}n��)����(:�N�R���&�?>�m\(:��*b!~�� )�/~}�ͬ_B��_�8µ@i��3��>Y��}^���eK�%�������3�R$/���ո����"_s�Y�J�K�<�A]=N4
��y������G���` i>�/w*9TW/�x!3I>����'��x���A�!iޠ��:�0h*���}>vUv�V4e���Oy}�,7i!	��0���X$gF��P�<�Rٺ���=٫����b���6���T'�����5�K�)�Hm�Uf�g$��� �	�Xu�'5��-A1��	Y��&>�z��3��dE��-��U>�?��_߸M�Z�o��ߘ��-�)�Urג��[�8���.ҫ�շݪހ��SӘG5�`��u��Bm�(�Y�{lm�"6�W9��
�����g��@�K���K�-�q`j�k����+V�|��<%�d��tʊ�JVۣ��� �#��?X5b�K�yơ�[PW��_XƮ�\fyd<>�N]y��'7͸3�`�����"^�5<+���X��v���E^��`l���G���d�i�q"	�ޡ��F%>ꛮ���⃟������)uj m���I�Z)ݙ~\y�p�?jhAL	����4�JQl�c� Ϳ6Tx嵛���*���Д1%���B�=3h��d��z�e�u
���8@p���Zph�����B�n���$�
F
��-� ݶ	���H����r�ݔ𖅶ˉ�@�,�\&�]��P�:= h�3�<����1���gY�;�MP�B�\d�Ž"*���:��E�i�փ.7�2�O�3 �d��v���S��N;WY��p�chU�!����G<��6�>-�_��E1a�����`4ڶ��=����;�ŧhZkf��ƫ��[T�ě��v�����j~�� ��gle2��d��v{���4�֓s�4�8��6C�M7Lm��c[��݅���ݿ��A��H���h�}�-RE��̉͇����Ҟ�!��E	p�"���j��B-�Ί��;QL�����=�� B�
n�&�� �&�i/����� O�%��(b�'$�1�B���x�˩������,��q���0�� �S5��<�Q5&���I�>�� t���C����i���N�muN�p�]�V!��a~8[U3C��Z��V*1'�_k(,�G��	�/�$���W��a���s�ݫ��� G�Z%���И�}�<!`kd=�d�Q����J����7�+[4���;�D;!]�m����&���s^ls��S'�Z��E��{�#��-�y�{��h�4��1["���p_���yY�ӝ�RG��Q��r ; �,�u�P�*���Q���d�ű4-B�����؂���p��?~�VF������B�K��>�f�G�-�l�������ǆm�[����~�A�K�]���e?V�M��*@H��U�wU�Z�w��!cI6:�M����%%�Ӱ�KX��鳰�cɍe��5?�]B%��Bbl�eP�W�6;�+�ǽi��3e< =O�$��ҝw��h�6���*O�,�@	��q��x�@:,&�C��	bs2�1*9��0�ւ=\��䊫�]W�+_�J�Ks���ֳOh"�Z��z5�*���V�:��@=XnP4��"�k��9�J�8���+RVZ���	p�G�n�S�H}ݚ Zz�#�}U�Y؋��O��2p7��P�0�@PdO���M�/y9����>I�ȣҠ��%��6���h ��yΤ�]j>G�6@��Y�ԗ@���:?��1o]IB���Dm��0V�YvFW�H�"�㩺��p�!��]���L�������.N+���dF���"%�r,~��w��	��v�7��������W��n[��Q��)	e��Ud'����sӰ�#���1ԓS��fYx\u ���@m��λ�� .�g�	�E�Pm)�*�m�]��5��ˊg�n/�Nħ�hj]�~ �f��¢��F9!PO/��ĂG,�{��1�|=���4�H(�H.쭇{��$�U�������6�9ff��|��^�F�8����Q��p��M]��wk�Č��a�x���41�!+�{�x�B,4��U!�@
H;�:����p��������L-]n{���`�!��q��Y��5�y�i�E�u�[]0����R	�%Y���������^u+s��y�6o1:Ռ�ܔV-#9*��b������`��#�"}�7�*�e��#�g���z�z�U���H����� ���f��V`�3��uhп	^(c�̻K�����@���F��\Wp�D	��Y�j_�d���NTG`���K�y�n�Q�D�Ÿ"�]�S:!�����XM�6l��:��|js�����H\�_L�	�����zSi��&��_0���0�t�6�l�� ��_����N'CW@fA���Wo��Éy�BK�Bp�b�	��LpQT�L�d��܇�z�8imBش\;Z�ߚɩc�[��U ��1�9�X��Bi��F�4���!�y�
�XX|�!���g,p%r�S��В�X�2���E���:��KV�C�𖇂��XGH�bD���j�'q�����YUyN�3�����.n����埜1X�����a[Ÿ��sM���X��/�|�m��	�tܙ���bk�16���l�71�(W��:H*&O��z	 ��v��L¯�º�d_�jj{,o�V���x��_��P3�W�F
��;c�˯*~�����'��@9gx���4��|�5�#[�5)�Ta����]�a��NQY6ֶ�����%�?" �%�~a`��q�_�H=]j���I�Lv^�s�vٮ�*yOU�T�kIҞ����{��<�C�@�x��S�jsW��
��pG%�@�{��#ŧ�A8b��є��U|����}VVwPrr]��R�ț�f�4[ux]��qs�;�p��|l]\�u�eR�yo\�bn�d4��G3K�<�!���Qu�Z5Y��	�wX'vG�����@e�n�Ɖ�(a da껉��) �����f��X�I�f��t�Ӓ�����O����&F(�l���$��Ѥ���iK�*M��ᤉ���CnG)�����k�T�U�8���#���'��BI��X@�5Kg��&1РO����-P/0A�Q���-�V��n?�L��B�����ڔ8��=ht�Cu���3�$�A��l1a�m>�=ѭ���En+,"��j�A?U+W�`f��7��C�b��2e,��ƅZ��Ѱ�!+B8D+�α܈��-6�uK��[��6/b�@Ss$Mi� �$?�X�Y��Y?�+�:z>��(]�K �#�/N#~����W�FD�~蚷u*��G�x��U=0]r5u+y�8��6�W�dx��s��w�`׻I��\�(#|rOm	�8�
;�	��Y�eF��i�b�%�M���f��*�����2��. �ȑ�1-O?���
����#�x�޾�6Bbn�@eO�\��m|K�<.P[Xb	�9��%�HŊ5��7^k�e����w����C;��.����}��g�X^�7��3&n��g@�*5�G;4e�Θ�BVn�EJ|�c�9wq�z��\I8���M1���l�i���ǫ�	��ӧ���j-��׈HL�d�xx��%���{ r���4���+w�G��Q�/@��˲%k�ru�H�2��V�h�'�b��L�����WTz�J���D��q��H�rY�@6
���2w�mw���	;�%�^���7��c+�-�7��6e����{��7F�-�D���Ն��-ޱ�G'�G�U'�R|��*eX��ɰQٮ�JѧZ����b�z��dT��7�>�����W�.#_9���M<�JWO�d���N�"8}Jf�'��	�᪽��A��6�W��i�D�ݝ}�0�/J@8Eg��w`�1����?�Xr�\���:қ�$+�N������&���.�}��nv�6�������7�K4���B(M�z�1��u&�u�|������R+��Z��ް�_G����	7�j�/d��,�3RF7t{��� ���fO�u�����4�s�P�v�KI�c[���J��AEe�����=o�Ϭ�9�$�Ӣ�3�r�� ��bP��'!B ���"P�J��o'�&v4�2�jZ6���9�MC��DC�<5�|W�Irё ��Kƽ��~�8���������d�������26��<�8 oKK^��^ ����{������&�'B�&�"�oțN�u�����Y"�2�J;�(�����2`���D^(!U�i��Tb\H��o��d�{W_��7�DN�P-Wy��������x��T��8��)���y�v��_��f�e�� �����_q��5n��Ǡ*�G�����|׽���D�cx�ar��W��>�l(ep>�K(���7������h�Z?=$^b�e�Z�V�d�5�Z{p_��x�I#3TmV�XZZ��G�7Iο�q�;$Bʍr'l>R�Ȟ�JL͉%�q틮�遥��X5�o�	�o�����b��Ʌ�qB*!LRw��Wy�����0�t���Ru�L+H�����.8�a)��{�`���<�R��.#��")b?�e<����H�H��UL��KmG��y~�ɡy�_;2N�]�uj=�Jm�^lo
�A�=��ط2�g0Sh9���\'�L��r'6&�a�E�X
;j������$ɞ�����o1���Cn�O��jU�������'1N=rE9���� $R8�����7�]����C�����6\��e:�.	!��Y�7{ژ���5l`s��%�X�ӡPL.�O�(�-���k�VA�R�4�%
��B1m��.I	4��>�*+r�@�	h�J�A��cX�k�E�#��$�ŹnQ)�ڨ�e'��,|�U:I×��誉׎do�=凂p���*����	C?G6����[�@8%^����i�ѕ������ �=���@���mE0�[T<�]��	��`w� q�q�fՃ�x�x��7t�v �G�d�
R�f0to�z3�	wE�F��츘?�C_7S`^��X�4�'��?��ě��5��k'��+��)�]to��O���W�Ğ-�\�	n��/q���s ��R*�����Y��76��X����_��� �mC��p��cR�<P�Z��$���̲	Sw3����}l�9��v��2�͢[�y+Y7��}���yv�I�f���@�!�e���T�`XF"h���M6#�T�)�O�j�w��Pݲ֧x�F�:�����=�Y4B4�ӢΚM+�kGĈ���D�6����SaI"+�D��58���8քIwfjV�Y��*�ַ&����J���%�aR�qR��ܪ����5��D�l�X��tp�o�A\W��B��7I����!I��;�i���ߔ�h�+��2��|��t�Ɏ��KU㒩��D�j�\oL�'H��@�>�|T���������Y(�X���7�[C��T�??5���z@!����6����HD���)�h�m��U��mV���1�h�8�>��ՍPFi�/�jh�"�Vyrex�`R,e# Sږ'j�zk�a��� ־}�6#�?ʯ�h�G���x���]J/>�9K@,�?\l�5�l<��K�m~s'�a �2��k,?�Q�GtB�E�*[�&n�}�� /�OSG�8��#yY���u�k<��vX�oI���O�-]/�.U�Sd�T]b�%5�����Q�B���-��Z�ᡆ+o�.�3gdr?X��
���R����s��/S~ â�P?�H/��׸N�O[����A��oWF��!�*�h�ES�4?p�9�*��@T��EU���A�����(oa}���Í�x�P��ݰ`6P�/�*/]�nw=P���f��9"�.���S�L�\v��8N>S���1����y��SK��&�bE��o�򸬛�V�'!�'���|�%H.C�|8�+�ꍰ6@Tb�8&�X1hd)�|�H����֯�ތ6*d:�pXu`Oh\�x�~�s�+M�ͣ��S��t��Ɏ+��`Tl��:�, 5��+lF�6�im�+��c�"�G[١d�q�Ǌ~[<��@X�^�r�J��Q9��g�j������b�/�ט�P��'E"1�oM�q2@���������p�ҡ�*����}8�/lJLίW)�L�p����Ƌ���r/�;���T�v	x� ��+]����l�Lp�8Nz�65��MF_3��f1���`��[x�	�ݎ�����$����E����=EY�sĹiƩd=�.���W�hf�����y[w���昌)F�s-���U`S�K��!�Z�s�-��eʖ�~�=��ߠ!.�>�8�x�x{���;1�h3�̠�)��H�B��ENZ�p��7��0����k���Okè��l��d�d�FW�@v^��5|-�|��	�]�P`Y�u���mX�ŵ7���C���Ce�w��^+�����C�6��7�R�dk�Jr��J���	���Iì6Q�xn�K�l� ��%���j�ܮN�eq����ÓD1@��υ�������Y`�e���5U(y�%{�]Ιg��*?������f�v�vK6>�ef�g�vQ��g�����#�W��1*C�G[Zi;�H{�|��(�F�¥*S��������k�/��w�v�}���3j�{�#�����_!�fi(6r�&�d��j��Lk�t�H�n�����3�v�1�e��hږ/a�P儷�;X�T���[A����J�r�T����P�eE�
x��/Z��t����y`+ wq)k�~I��Ԅ9?�T�1@��x6��g�����͗W��9���'��FF�� ܑԀ�D�����c.p)2�@�.���Ɏ���k`�lwb�`�`�:y0���%��Z�L����d�NԭӳqbQH�5-O�98��,�mr�	� �ω���KK�������)&Iꄛ���C�D���^�~���{
k�
Ж�0�Gݓ�f��I�꤫�B���j���������1���R�D0��3L�NS�g�
[HU�D1�A��-G�4jkf����616Yy5�2�����m�Jf�/�g���r����~�Xoʚ�pU�43i�d�.M{�v���7�|�ED��������7J��0>q���0���U� �^:�S���];�T�_�А�H����TO����7� ��^>iu�Q|@��I�al�����;4�U���W�\{��\���-o��\�>y����j�&5�n�=��Ԇ���=��(�@���v�d���Q�r}�(�
��_���/�l1��{���HU��0ࠖ�W�V87D�	,<��H|�d��u'�ta$d��D<)	k�~t�����^M j)RLp�xYвK�Z����>	S)h�: R]H�}������28��FL� ��)����cu&ݏW�X��p���(�e5���:���w�|��;��}�ء|���R�A�ཐ{��l�����b4��:��N~�����&�H�İN�>�=�G�Tc�߻e�X��i����"�����2"��;���/B�:��«��
��	�J�E���"��7�iϡ�N�L���0��q��(�Uy�3c����?��}�2Օ�YTV�i,!x�oh������}�PΨ6��u����0���]l���&ǳ !�b��̣U����� 54�cu��j?u�OS<L�V�g��N�
�R_0o��;��1�R�#Y�2���-:��8�&�	�D��4�0e������2���N��Ჯ-�M\r6���1��t�B���,���?�&0ֲ���e9m8ȥ�0ƫ���[Ud@�2�Qcx&�0~������N���g�)���I��MJ0��-�0��Iˋ���G�3c=��.aS����]-'�����g�y\4�u�Kah`�4����������9��~��9W�c`� �0�P�@��a����;!8�)Mӣ�܁���	���Ɏ�� ���v^U��^}LY����.��}�؜h����;k�]�*�ޠ�X+�2�1`ZLl�&����PhH� �V��$����jU*F����g����Hl���H-V�E�Z��j�����Q�+�E��u'�*�ņ�Eh�dlTF~�#Q���� �b��I� 1����B�|K��J�K���5+x
I�d�@B�eT�I	/8����`�g]��E�@�����c���uPG��Y?E�/�+1�CW��#��%Q�pl��Ζ%�����tDH�Y��@0t�ذؒ7&��H�'���V���k=���E*ʎ{�Z��]�x[wE��Zf�}9�l��Nm���u�S����EJ�ZQ �H�~����|q��3�%zlxr��g˗�!�:��8]n�/Ӆ� �d��>9췮f�}2;�[����\�?S�ñ����ѸlEiX�G�/q�\!��_$�eo�,�!�����s�Iq�u��v�|� �cF*�$���@]+���
GE/±��^ք��EF�;:O�%~�xR-�;�S%bb�GJ���^0��%cb���C��{���P�I�%�'��/�ղtc���(����@�mL�b>��-V��*�ߺ�W��@މ��vZ~�`��t�Qa��2�C�6�f㢰J<�~�Si�MdJk��T����%�B��w�*�`'��6Ƿ�"��]�ݟXYYҢ[fG�SF��/|G�"%8�������זZ���u�䣤0���R�<���W�-׉�\l�Z 
��h�>Q楪��%��-s�D����J*��w	�8}�C¥�����Uryϖ~±/��(�+� ��+׃��
Vw|�6/�QQ���Г~6ZGҶ��a��rXH��?G�&]�EZ��G�,��IepV'֥|���G0?��C�h?ca���3��,�QL��:��}�^�_�i���IB�v���}�tF����s�m��Bݹ݋o ����-��/�|��qd�,h2���+F�.<R�!n���ek~����vWs���T@�SR����~�2��*���aU�\��<��֖���$*���z�ݷi,��>��ȽaK�!��`}�MxgΧn��7G2��E�L�����Zx�=�^�.�$��vMg�7�8�2�K��E�{���޲�*��T�)Y=� ��}0W���;|C���Cn12
�X5q��:a%Pwn�Z��7����m�ѳ�q !B�����ב�&`�-׹�ߔQ�T����j�@b�丞G�ҌS�	ԒBc�N�7
ڃ;���u�[�r]��!�|�t�?UO��W�-U#5r{�Y�`����
@�!�h�b���V��,�rۏd3��K^��L6�z��j6�	Y2�,O� Ҟl�+�9S��
��L��O?ރ��Lu��;	&m�!PU�p��<�φ�+��|?��J�i�Y�Q$�a�=��W��9�h>4�q�5gj^��6Z�$w)�.��u��{�<��p�Yu�S�l8���q��S �gW��:��gؖ�MW�	T��/y݁T\��^
4:}���
=��K��eq3	��ZN�5�:�kɅ��ൢ�Տ�q�4��5�/��i?ۻ"sC�ha��	����;�ӪPcADMHΥ�H� [�#��-�_}ǁ&�����h6�;��D��K�oV�@�C��*Kj�������P���wFu1P�p�Ǐ���h��>�����.̶�p1*a�O�����SXh�X�<���V�j_0�8�
 ,�:5$Ϳ��c`C�t���T����;���1l��T�H�3�9LC���<�"T�&3QK *V���'���Չ�dl��.~^�������t��8Hd�c�����
W�V1��#-٣��S{�V�'H`(�@ʈ�޷U��q�0J1��@�"�,�s�ZwkH�������X[2�V��w�e�^ �E��u��b����vZ�n&�(@��BA*���h|�F���r@1I�8o�a�r.� ��e�Z��c��(�uO��f�Rh�Vu@G	꣎E�Kh�i��d3��xŁ��wY�ىWD>��1�G~?�I�K�3����� �5�\s<���8'�hx�]�3^�+�<�2�������+���dP�5˳�{C�ń�3�-|4̦uK
�����Ꮒ�
����=Y�Ғ�YW�J+�\5w��)m��tDDǿ�����nuڑ�c7$kM�,���'œ0W��ځ��k̯L\����#��x�0�-����d0�J*��t�^����1tkD8~�fo����"[���^�Q{�t!B������ ��{j�͌'jwqBG��x��SD���:��WHˉ��-T��UN���KO8jsB����	w��nQ��������p�������Q�����yZ^��O�����YA��_���@�����|[��h>���K:�<6���S,��M)�Γ��v2lE&�J �GS��GҫH8�#�fC/���`���l�o)9ᶈ���`��:
ԉ~�Mf�^�a-l��G���	ɡ���?��"�
9�����atͿ'Ѱj?"�Ś�˲u7d\Y�yvjy �A�}	&����f�����͞"Ƙ5k[d��L��%�����)�U�/�,h��$~Bo�$�'�:�p�7��着����8	z��4]����o!��kF�I����H���o(޾"���4��JϨlOWaN+��(��f�3�2�=*^�spJB3A�_�	���{m��6��/R�j��L�+�U3~�cz<�������0�?����ϱ�F!#�<Ys�0V{�$T7��MP����z�!r�o�E�*r:��j}���|4?Z�yii;?��}
������5I�;2� '>�@8b�u�R�����"71H�ꐴ��ǉM�����B�/��
tr�OBQT��;W�bcI�l��*[�u�r���_ОӁĠp�R3�����zm����2K�ʂ�9�U�=�S�~["9K4���?ц9��b;�� ��Bv"�q7�/�����]���k����Nd��B:��J���W/e�,=��_l��ҹ_�0���=�}kfElU;
 �MҾ�)uD�x�X�5� 2Y qw4��{�y2���T��۷d���;�H�UR�M����tD��;�k=*!Ӵ�4�[VL[�%��-�)"p).�����ܳ
U���U-��0�$�� �$�.-av �*q3�I�|(�X[�k�\�zV��䈞=$���l6(��Ăbc�پ��i1l����}�k��w�*�gd)�����|ΰ�XG�/�2����$̔6v�`ЯZ�|f�o�Ƴ�"��8h�S��Q�
䋄��z�4O��&�_7���{�:�.��7��w5,.m��+�J�/�<�q���.״{uD��r�m��`�6�=>��0�GG}�Nq��[<��/�ZmS#��b/�*���#N�-z ����ML�}%��������U�S�I���{g����[�t]���{)44��d�0�cξc�]#1�P����Z�Hr^�G��0�/-7���/�=W�:�9�Q�/Y��4��$�ﾽ~n[R�Ϛ
+��zb&MP�+ޘ�t���f3@���,�N��7L��)�ѓW����g���3?'b�����������k����l�ԭK�!�vR�jo^��'��|��6"������6��q�$�'G+=�qi�w.���	�T�o�3~�Gd�0|�c Z�D����D�1�]f��QB{���:k��B	Ђv�<���mn<�%��?�v��	o^-��b͕t�J4������zs6�H��0��� C=�U�v�'�L�7�P����4��񘥁��XUg��%^/q�қ�4=c.��t���}U�1+���ae%���'o�w���	��S�۩�;�KX��M�W�Z6#9�b�m\%���4?�B�����=h�|s`�Z-ܓD�m��q�u�HV ��`�=���Z��}>,�q8_��>���\bF�y �VA��kJ���dY�Qq)FB�'���� ��wd�l6�-v�ۣ( <�r�hk`�?E�H� G��>b!!%h����|ᙙ�#���/�MC08q����h����;fp��4{��]S�h��߫C���2���^���8�q�p�w�:�*��#��Ҳ��#�g��*b��%"D�c�i`�Ԥ]�G��g[�鈬�s�� ��[�r��[����y~��=f�5��<��A�Q	�m�H����_����z�Q�Df�4S/Ň���(1��P�g0��𻌫����ö�4]0�,$�%�:�7F�/��=����8a\U��Q>9�ЯLr����
�r���x{���Q�#�[��x�%g˵m0S����ٽ��y��9E�/���^��M�sc���6�|����[miG��G��=-.Ѵ��(U��ɦNvA�����4)bZZ��E
�͏,t4 �¸n�_F�ֈ�C�����	ۨbl�U�������jw�l���ς7>4��	w9�-q<��B:B��cv����	���y�IV�հ���zn ���7��O�.1+����U�R}&\��	��.��9Rr�E�Pb\3U�,:���ļ����E\�d?���p�3��>��������qy ؟�z�'���|��G��b^nGTc_zwH�>��G�7�Q~C�3����!H��z��c;5�9���Y�ʋ ��'�+���]F�|��������q���-Y�Hu�\�٢�pp���� �w�gq$�̰�N��+�jD�A�a���.�،�zv�X��w�%��S�
�<VL�]�A����DSU��&�UbL�P�YV��m�g:�7�����Z��r���?Q_�u�E|�I�)�u���Q��|��僮h@.��k ��ԜyzV&7Ő�q��U�l�j�BG�XQ���<)�f�]�U�T���r�"@��\.q��`V�s�����A_<����ա�p>��a%2����Cn~�Y���n�ѽ�W}������l�mN���
��v`�P�A���y�����^23O�*u���X��T����M��FE�]v�`�\���5���j�}�ɐ�`��ٜ:��Og�7Wnx~׶�SgTwE]JU�(�H<�
e>�8\&a$����C<|���u3�4�I��#�Q�9wߗM�Q[�_�@F�WY�S�,�Eyp�3�s���&����n��_,����c�D�W	WW�Z.�»�h�K�O��j�녯���l�OcrM$����Ҟ��!1���f�~�yy���^Nv'̍궣�[���h0����ʢ�
V��b�S	p��(�
}��W&@�5,��� Qŗ�����ৢT��N͑M����}�����x�<��@O���w�^}�hh��Fl21gYǏ↠j��X[�[JA��>��Y�����ǫ��I9��O�������E���8U���\�Dc�������}�U����U(�1*�-s�KuM)�c�-����(}���џ3���)m"`�?��T�}4_��w1���ĹF}<8� ��Rc|O�g���E�m=Glؕ3�g��V��TӰF�B"��P_$} ��&1rW�7�����KۘL��k2�O<Jd�E��q��%� O���N�(QtD�Ӹ{[t	�F��~���=��B��,��#��cP�q�n�z�{]q$�/Ø�0-�׃O�}�~�i�4�����!>+{;�[�q0Fox���$�@�Y�_��Mc)�3@ m9A`��(����yz,�O84ΫZEO�F��W���R��޴c���*�0'������7Ȗ>A`��Y�����|ғ��I��gٚ�1%fen���F]e(;O���~�;_b$Cu��U�a>���гT��b��QW3����	/��M/��XG��oվ��i^��a&��0-���[�.�1��*/v�����]����|#b���{ C����t��A�����>;�=�����űm��R�a�3Σ��$)����J�wW���G���Y�����;m�xk�l!�B�7����9���i�-�d�+?�q�z��j������xyaUgK-�?���nH�Ѫ�o�jU�Y�)p�}GO/ŗ*d��>�W17+/0H��S@���떁۶��P�y���jM�=eC�$���U��X*�!�����N�aP6?�2���65�Ȍ�����ƬY�Dt��kP�])�+�S�"��cj�7�}��Cӡ6�57!�8�R�ںm]��_;�N�����(�����"�g��c�%�c��\���"���o{0���oC}x��#jwُޑ��6,`����� 5��������\{S��;Mf~A�%��:��Z����}��]&,ޑ@�|ŨF� ��Ğ|��S�$|�t�EM�	|����ܪx2"b{rQ�� ������?#��3�������`�rcd����☷	q��M�v�8���:&}!�ZG2K���$��y�Jd?�.<e��
��	���
�9^띳F���|

�x��M��|4��x�\ 	C����5
����=VD��M�p�Ր�1�xMMک�Y��՞���4���<�{3&y�-�{�ZK�ko9��Iq��I1h� �$r�%'�M�9$�"���Sp��.j]�n�X+F��rs=j���ɉ+��,�s=�i�Sv�_�v��4����=Mj�^-EW���s�^�; u[O�<k����3U���Ft5S|�ӞP*�_X��o2�H���+00�PX�����*lV��}�?�]տ���c^�`�)���������'��Y����$��W�o���9GO6f��2��	д���("�B�p�
J^�����5w�JE�팘�0I�;&�rT=�b[7���e�ը����~&M݊~��%�&�ۭ�"�32|��c������4n} 
- ����4�r0f#�b�a�Eu��f��_��h�b�S~k�ʸ��w��h���?�Ȥ�����I���������՚$�����$@��"�A��*����Fɞ�ibv�Jk���P{��JX�Ņ垉�t���s�:��Έ����i��ʻ���-�q���R(�lJ�j1Ы���/����4����v���W��;G�%O#,0�~�z�~{�Q{$�fH���3�ekD���6Ee���/�t�rO]��"&�c�-��s�&�"�������b�~��`_`i+.lC�%��u�4j�J����د�~���W y��`RD�vT�o.�(k�s�o��,KJ�j�?W�q��Z��Mu��W�%JzT�����;��N�qg��vͩ(�"L�$�!�
�T��B_я�?�W����>��_
@��^sQ+釐j�$�-O�!��-5��0���<��]�ݹ����bE`��.�6��*ԭ�.u����	p�H�˨�BO�g�
f����s3�~f��y��$���2�fV7��t�=f������"�	sG��ʢ�Etە�s1�Ɍ�(}Em}��qe�0�%'�	*)]�tq�d�p`�XU�'���W�FC����FY���|w;����=5��8Թm	7��hN�:q	��u�fKY3.�>70�ҙ�9�������ذ���O��8D>�饃����ė�6�r�z�T�V�CI)�p��GR!i	,OkU-�HGG5 VZ�g/�O��u2
i�8@-=9b���o)�9���2bYW���&��,`M�N���Rɇ����U.�~����P�h�9Fg��Ġ(�攫(y�����JB+��]d\=K{8��.�G���J�xUa�,vUwx�%��66�})�ģH�X��ﳫ�A�撋CnG�}���/�Y�;��\{e�`�`a�@�kX��Ô���A.�.a�J'�k�AG�7��Z��|��tf�៲b��G1o���DG)礔��8/"r�t���Z���]J��K�^�f��c%�TQ�����KFH-��7���Z����wYwG���Ruc��^�ِ��}@��Ϝ��ѝF�>����꿺>b5v+�4���u�jԈ���z�8=�T�A�"}㥭���؞4����NU�k�v��N���n�zy	��(�&r\��杵�h,}P�|�&��<�jB�T�}>�sa����x���㐿�'����b%k���h�� �����Yq�@L��/�w�	;��D��K����z��4Wv�qG�HH���;�de�����p{
T�]�%�Ѡ��-������s^A���ȵ��B�0\ê�����Sc�m�!f�������7OD�Ӥ������(^����XFC3;�(������b�ر����uJ�_Q�v�߁R, %k��ۘ6�>�yA�]sh�I�h�o��r����:&sx̄%9�4����Ȝ���c�/54��|�'��lm��c9���sэ�
��P�� ڽ��^GA<*p%���2W�����>7��_P��MQ�F�KB&���r4�H�
�S��{�iB��M�J���{�d*i�PС�U?R.��]�v����#T�ǐML�y`�D%�F%f(]2*9-�����{^N��|���Yp��KV��Z����*>c���Zvv�
x���km�v�DhMw�.M�+����[-|��1���8�H�ɳ4��_���"��n"�P����O]L����(n�� ��:Ö6'o5W���m�B/Ś-> ��Ib#��B��0S2��D�P�Bq�Dߍzd��ϥJ�ix�-�D���D�0�ùU�R'Wv/,*	�,��+T�[����� d�� �$=Q��&X����J��J�8�QG��%�>T
��i�bo���������ڏ?V2�cv"Ü��^|��3�p;L`��:K ��ג�����,��9�����%�~����s�\��� �R�z��3	~�B,�ߤ�HN�ǽ�Y�3�:�����X��s����2;~H����H��#;"�X93��x��ǮS���0r��D�W��|��i��G�S����klw՜b�ഏs��(�@�fc���f<�kM[��es��@��T�f��zln,�H]���@�P��X�
9�R�tIqv�.�2������$���k��Nd��Ɖ\����u��@�hS����a˓� G���f���N���� �nѰ�����L��L|Ϛqʇ������N]��>�#3�O5�a%7�
�8�׶�>�C�Q������R!O`�h�|EJ�����&��.�)���̻���k���Jt�s��@}���d0�6l���3��� ��|�=y4���O�0� aV��z�	�D5q0~:�[�^���"�4����=K<{�g�42x[,�
�UՍ3y���Ԥ��̿������؏p�P�R��t����,ƍ	M�``&HN�l�Gm�>��/ݪ	SL�G��X�����`G��lt+��N�w��e���I��kl�;���?.��h!�����ݤ�ғզ�c�[;�[��/��ݔa�����6��%J�L�,XC�Jگ�rN�RS.�'_5�;U>qO��nc�U_��赑3��J˭�L
�B�k娑�O[+c��|�{M��9��(	:,Ji'�%��Ƨmr1r����D���Eܝ��j��
���~~��Py����X���L�2-�=G�e�4�R��_x�8Y��'*Ge�-"t*e�*b�y���c5� `���F��t��7�m�Qdo���� -����E�L�����������/���D�ŝYd'0.
;���jR٦�NЖ���֕B���L1��x���evv��k=1zy�-\�@z(�~&.�b.a����@]}�̯�$GϠ�*2�ѵ�d�x�}7�ؗGo9�^�6�)�:�vL$!ײh�� ���W��X#�� �*�-K_AK�׿�Y���~�3'K� _��	J)��@$Awp9�+k���D�$s���X���
Px��X��r�Z�@���U�'��|��r׍�3t*#�zԢ��.)Ik�u_�\�5��Bg��@��Tf[{�<���*Tʇ�'�î����Oƣ�ʕ[��'�7�S���a��Z�2����|	��d�`�,{4+5��5���* \&����%?��z����@�� 4
K?�g�.�<D�,�|U@��:�P�}rX�h��J��&��G.Z�W�:/��}k��@��kU��>�"?��J��8[���L�����sv5��K�C��D;�h3�~��o6�G���&���
,��p����m ��#\[�*'�L��=�g�ş����F�N�'�V�fL#w�����/
���%��nU�(*w;5l6�W��������U��}��Z�����L �����]t�ĩ�eHc���n4:�u�Y�X�52��{<��)R�c�~˳�|?R�c,�o�>�8d�(رK����{v˄�I 	��Z���ϊ�ǂi˙>�zH#�i�	���i�Rg�(���\�+_��pi�X 1��V�;~Վ�*Qzk^7�M��%K���_OL�Ov���.��F�/r�wP������%��X�5�X	�`f������d
(��P;FI�ۇ'c�*�HWvbl��+0�+M`�h���[.�Z���x4�(��"�-{半��\�!J���A�NTa�v
�st�u[Q�T�<��&d �8�f�ș�;��R��Cy,49 �"xp��B<򡅛�3�Ҭ�4 �����cw�O50?m���Me�h_5E|���ݻ��k◔,|��͏4i�����ϧۍ˫m�J��B��f����;�46���u��0��:�q{{�� ��@x�g����0����ɇ=Ș6�y*��r����7�;�����{Y@(Ad��K;>4h���� vnJ�Yw��*#1�Q��e?���T��p0��X�*��N�h�He�2|YǚN�:ڇ��U,g#��|�mxo��q|�"�g�)"���ڷ��x�v���>�=�خP@��N�I��1�+
�\8y�<�����a�Kg^�'.Mځ�쎍A��Nt+;wu���'��+^i��r��Ĭ�x�)��0�����~���H�Mċ�v^�Ou�����f�I�Е�L�>������=�B(>����:#�L	-���������׼�l��۲3��E�=q�) �
��꥙�m�:(�=������F�#�8�u�FIjl���#�(}2�\1A�*ŰWANmN�yPh'E��5?�4����z�5g�/oV$9�S�j%eS��K��,b���b��C_=���0&�
� ��P?8����2�}��qk���s��E��j�gUa_d��qI2�@��D�����	�u.�.l�篼E:�
�O!:ma����K�g
ֈvz���}6�>cM��5oNw��uʚ3�zP�K�{��YwcZ�8 2:w>.nk<' �x�����bA��~5�K�1��h��ry"^ٗu�1V�Ċ�� �a�lw���)���?�_9��r�����j�3�ʝ���+I�A��,�d�&[�����=���!���'L&@2LF8d�� y��dS龭�XСѬ~L
v��h�h��	[�I�jY$���e�2����b�8��p����twI���޵\��Q\3��jv�LDF��LG�U�=�����nd����=���g�娓��f����.�S������0�����[�����>;�Q�{%x�%��+�#��qHt�T��n���O�|�2�Y��]�08�Ncm����B\�=���u��R��8�Us9,�SC���}��X�)7�^���R�}�I��%�agb�4]@Y#�̬8�fg�.X�pMv�ғn��ۄBƿ�b4'��0D�	�_I��m���,�^2��}e�9I�:�s$( 1ʕ� rp��l4�7�^���lm�hS\�����^/��x[A,���Hp�-3Q]��(�te;K��ZZv,*I<C	l1�l TR �/o=��l��1�=W���8�0=9�"e��+WE�囒Y�� S�@P
 D��]����&�;'A&�Ys?a��������m�`������Q@#.*���j8�3F��i�D�t����G_h�()�3���+@C}��;�K��9�?���o�,'������d����<7=R
�V
j �c���Z�?�%�:�?B�ڊ�����d�0骑�e���D�j��-=>�O6I�����/ �믑�:��[�X�x�Z#�j ��|�0�ƀ��Ȟ��:���N?���C �(�;>�q�)p�	;}m��P��n�R��_���c�� ���y��C%B#w}v�ꇷT�o��Z�޾2����,�$s�<ի�G�|c��5l-�pS_��5z�5;�k&�gÞo9�}��G���
JV�rN����}��pEC���z���}mqF|�ay��+�]���[f�1�N��.XV���%�w���x�
E�����N�8���k��CɰP����N+�%����P�j1�:FЇ�t��nN�����ۦ�I ��2@���F��j�i��Եţ��b˖<���:�ŻX߷�t��r~�=&rv��R 	����í�rO�T�`��s��P� �IjxsPA% %8�ʬ����H�yD��נN�nJdX`5��EU���zq�杔�*��O�����F��6�(�~��t��T]k#�ܦt��K�&��!�[ԋ�n�S7����� �ѹ���y|�L�ԇl}%�<��r{[��-��k��4^���ȷ��D�,\v�LO=;]*]�"�w]��v:c*��oN��~ށ�+� �4'����¨nIG�Kj��?�O��8�|��n�2S0�(/F��A��0��7��?��xĔ�\*1M`��bJ=J�� ������<h��CDN�t,\��� 9�+�+V�t�yS9Q��[�6�ǌ^/��16���u�����\#6 �*�	t8!�<R���ĮTw�S��.D��[��#�dbv=@��~�|����o�Y�!�t-�2f
fk{���)��c�F��~�v/�{a>� ߌ��+�٠Ӂr	p�ȶ��rYs�ҋ+5I��K�l)Ɖ��=5Zk�bB�l?R�͍�n�fq�L?��_�ׯ��1L��`g�l���੭��I����t
O�p�g����[_�� ꅁrzOmׇ��z�St��v�E0����k��9x�*j�x��vc>H�6ᇦm2��bs�g��~��Mשg�`��!r��D�@4�.���\y�Xa+K���4��`�9H,���^�~`'R�i���C�].���{�P0Re��w�Z(Kp�d#��%�L��mK�KX�Ń��_�C9ޙ�w���&ވ��z����X�tA�- ���k[.�(eqչnE@��\��V�O��/�~=�J6�Z����iR��S�m<�:8���O�o	[~f�C�^�ub��BHC`��Q�9-*���W,2Q��J�b,�MK����!yQʜm��ռ��e~\��Tx�
f`��1
X��lǎ�����f�*�K&VkF�hW��;ɺ%o5�s&�u��wԑ��xD�AG��<UCQ�;�b�tu�(�2<�W+~7�To2E���L�J1H�ӌ�&�

ׯ�"P�`?�i`����
�z�^F�� ��]��θ�:TM��S��"�;'�0�dv����3�+���d��9S��sz�C-'������2�?�": �	��̳��7�I��Z�1��"��A'�*.���B7T�EWҨӨ��[�)m��ǓۈU�k��^�z~A���C��a5���nH��Z��A���	���}�\*D�����߄��5�65a���k����<J�Lz�ŨL�{�!��Y.i�kHmJ���F=�`��>��k��>b*�$��7J��v��-��_b#��Ap��-�h�"1�ߘ������	Y�sdSC��_����^,�
Lç:p?��vF'��7�	UHe�p(�9Z���0����PE#e�2|~��%^���m	��m�{U�%zM�G�S�U���g�{g����5bx�:��	В�?q��N���$��(|҆X#�^�\���G_�j��OyH����,7}�� ��T�\M�`$POP�P���;K�c���/����a��*J��ns�Q 3"Y��}��;���?{1��^-�;ft��=�CY�n�Py���Q*h�&t�U��8��;_ss5�$EL;`�V�����d�5="H;ʱ{�~�@�������8FW?���q�9����9�fE��",�}WVPAmO�Y�"8;?D��%����<.Ŝdi{v��*;��'e�+i��|N�$	tͳ�"Uh����y��_�х�G�b�%Ϩ;�IQ�i%��u�D��h;!@
x�R�:P'�H<ߩ2���9 ��J&�cZx�ٗB:5�팡��I�|/�]�����p(�6wk1.�"S��BS~�]�z6��+�r��<�NbKL�f���å�v��
G�WjC��4[.M�^P��/9R��.f�q�{������܇K{�v}Lx��5��s����u�d����dk��_@�2J�&��KP���k^�8��wT��O�:��a�J�	����.urz9H-*@�L~��B�s��s�eR@��"/���?�����9b�2,��m��\мh�oBj��VC|��ڠ�s�?E�o��/��j�p�IA�.�����h����`��=��[Ζ1� 8����A��fg�,�+z�����p�b�ChDm�$��?�.�t5��9Z�����*�[� �t��q�8מ��̽�A2�W��!^�j�����5�v�T!��F���"
ٶ��K^�6�#���7M�p�œ�Ӹ���: v��vQL�*]^�}D��Y�E-�VFG$�g܂]Y�k`ZT����h���5�{W|ά���MW~��<�۶�&"�������˺b�^�c�g:O�d&��h	�y YqG�/��&S�w4=��R�������ѳ+Sl�͟��Ơ���Js��P兒&/�m���#�N��~�k%�Du;�L�eŚ���#^���ѻFf��Z��_5��O6?<k��I@��i�#������jv�;7ыՠ�?�u�b�u%���Kn̎O]�QZ�~e�f�C!�nBrm��g5����1� �*>)"��4+�$#i�>o�)n�kqv��WBΑ4z�8-������C�����[n:�/bDJ(�{���ib7��ӧvsG�6c&��3W{dA^�%ˡ��1}@~P�u��٭��q6|	f&�w�Y&Q�'�ڍA/�~�94G( �\�ψ��qu\y����2�����z���w�h�1�`Y��@�q�w
-�/h�]����%�")�� ���.Jr���G�;d�:��� �bq��`�0aUL2V= �0"ymR�&���s��iOjύ���/�uܓ�\��:3�އl�Ww4�^��C�s`v�%Uxh�K�	�a;#��樹�҈�=��e#^��ad	
��l���3L���v������I�g1�]��\��z�:����'Yh�u6�Zs�фbl�|�{����me�a	���Iy\�<59'����$N����w��NJ�g�k���;�F_��S������t�U?z�u���}
�&��T5���Tjuw�����3O�$���qf�^����� �=��O˯/�-��c���ә:��s��ŐfQ���ۀ׌8�WU3�71HwT��;J&O��S/]�%b�-,�9�	�7�z+���.C�����泬*0�C0Sorl���u��Iӎ���7^��փ�f��O_�+��̅s�H�ft^�\)U�t]��/��hq�/A�n7?��E�MP����, /1�$y�F�~]�!vF�	��2�߃��T����N?d�Y��E#*`�2�m�m1����[��JQ];@p������鹢��#V�ye��Ԯ�u��x�˶���W��!�yW���`�-���%��y�a��^'e�(��8-�1�s	��* ��έ�p(� tD�.䛠Ĉ��s����׏Pe��N*�ah���&AK~(%����`:#��Zy͐s~y��{�d���hJ']�k(��D�Ta�N#�	���E�k��Ӱ�C� h �AQ6���b��"�Ȼ�U`FF<�?�W�0��-*�_Ck_2q�"�0i��$�꾑!��S�:���0{����M��Xj�G���oa�q��8�}�v>r�;��qzʛ
���|.5~������}���L����'w�΀��YS慄�:b��|Q��#����u���IS2�f����%���U�cw�Eȼ�)]�~��dj�������d)Ozڀz�вVىT�
#�/��r=�~a�R`\��yҢ��Bh��d�Fgv�u^��X�mK(=����$��4�]� ��]k�2w'c�\�Kl�rj<S��3�2pY���~���r��A�VB՗��6�I�7�Ɠ�^� ��\�/��/��>�� tF�ۢ�dy���C@3�@ĘH����'~,' ��:�o�Am�Dz �+d�y:��#r9�Tt>�tim<b��K��j�0���;	P�/��mI'�I{Mk�&������`T��-%�l�'U҂o_�4�+T��PI폔� ~���]9�
u�TE��L���`���N0N=l��٠ �q�v��~����]�(ů>���4ռc�b9G��MPy�":�ec��ʯ���5I�_<�*G3�x�=3�^0r6"�k�Bg��2W��g�2�R-B�U)o�4\�i���"N)���Gv�.Z(�h��s�r��2��8/��݈����#+�S��7{4�eL����ez�os���=�>W�"��D�S�t��3�����_��G]c&��Qָ�"��@��8�	���!�c���$�@�4w���x��CET�fo��On���o�N�ȍ���A|���S�0t�ix��T��0�va��&pS�w��E�gj�bc�P��	��	�������xV�_()�Y�����g(�)�.�d�ߺ��vj��G1'�*g;'�y!
�E�]p�q�5:�_�?�O�h�al����F1�zN�t���heR�n �I��AZ3�z=�����jؑ���j��M��	�9L;�j�pß�e�&���uw@k^��������w
�^:�yj�@�!]L2�Y��F#ؚ��)9/2w��uPz_,���p;b�t,h�c�	���� �$l�F�1}�k���FX����7���M�[h�#Z�dz@��}��UugYߨ5��I�P~�PAht��cO�ҹ#Wz	���ýH���
��;���S�����,n�x~/w��#l�^q��geޑm��*�h�$e[��\�bt�|��`�Ҟ7,���G!˺˔��/Z����W�U������	ܶ�Dp��u�f�v�$���`�r< ����J�c�d�3��u����I����Pǯ�̰Zz�sjHw�D��ظ���� �1\p��/�'y��^�n��������6d胒���F}���=랑6E�/31��pK�Цx�!d��6Qw�� �@p��"B�h6��n[폰����sw��Uu:$���IuY�NgQ)��L