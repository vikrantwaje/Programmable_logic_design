��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&�O�}>Yo� �s�:!��H� �/�J7{^�K܊���.U\|r��)��&�ET9�=�u�����	NC}Q���hj�'S����i���s(��
�y��3����O*S��>9}����M�)Q� �j�d���|z���Z�a�"L��+�/�����y
��]r���܏�p��5�w��)�Է�k_��[J�`u��]%�����8ַ.��(���#Q:��b�bˆ�w�z��o���l��i�3�h�I�p�>�)���G���Yڞ|Pf�nA�/����z�:���g�F*{h*.��z��Ax���2�y�u0�i��1h;�CdQ�vs\��F��TF�)kSx5D%�K����3S������W���.�Mwm��1`�1H۵$�j��}���!���A��O�s/\ss�UP'� E�َ�%��`tr0���1#�+���S_�+���/�� �"�1�C4�����2�h؜o�f�Z��Y�X!0.J�xڿJ����de���e�($��c�,���گ��)xb�
���f�3x��&٧g?ڷz1&��衸&��O'�,�.�4HN����$�� ��\5�CjE�@�񚳈%����Tb㍸��� �L-z͇+D�e.�cӉ`�
�ݧ䫴}��h��M�¸pz�9��.����"v��Ȏr���C��N2�)!n:��%I��x`��z�Nxq)u�<��i9��ij�%*��$I���C����������.?��n%��@�av�QV�|�ƪ�Bb�'��@*&,4.!ܙe�SG���#㈀������� �w���F�C^o���t��UN�ܼ[1�`��ڸ9���N�0�lR�C�R�S�2�h��v{q_�
Kg�/�wQ��m�u�)�Q�tf#�hX4���4�l���| t��T�����z����9~V�F�c��v���QP���ơ9	��R�'L��}��XS\!�����{��Ec:$P��7`�d��h[��]o�MI)�DhC~��C���{rN~m�XF���%���/�U�ԓ�^&.�6U�q�D��
�4���w��g0w����g���D�w�êD��jO�;�?�7�� !_�����(G4:�/x�O���j�k+=9Q5WIw�f��*��<�y���p>��F~k��Z���)�6X�VM�]�U���B�X���ܩ�Z�`�p''�{��1�eq����4�:n��6�+c/Z6��M��Nc�r�֙��nƟi�4iPN����/�M��|c|���!#$är�o�]����W݉����T�
M> �L��?��I���_�B���5b\�;�x��d(�q7W!G��r>i��C^CWMі��Hs��8�Qn6Y��dH���>�=�*n��ѿ�y�m�c�7��Q%�Ϥ�s�F|w,DI���H����Ɏ|k��P���5���\��#��}����6ΈN��lW�������m��5�mx�8!�>Ȓ�B܀������V֓��`'F��f��}� n$�:W�aaۜwJ0�!�s8�,�O8��/k��/�q�K�_�!���z�#b�ʺ�y;h�KZ*i���)�����f��@p�&�&"p=�B~���u�";���*wm�o8_�k����`���&׵�ciX��#�W�^�W4e��	|Dz�l�xu3�:R��v��?V���x�l�3�M����a�
�'l��煀����	��-��)���Ѳ]{cQm�\������?"d��_� �K(�y��ܛ�kH�8O��-�<R��e���[�CQ���l�@!�UJ0"��2������������u9�������Tw<���
�Dֳ�xQ��5���Mc��J�I���4�.��d�C�$�5��v�.K�����D��ެ:�ƅ*�s�ӶjJ���^�n�s�c�\�}b�>�>�ZB�6|F��UwXηa�¼ct>���`���r���{݊�'��d<�	�@푗�g	 x�OА	O�T�VI@+��<\{'ÏǍ���`x-��\3t�$&U�O�w���3��	�fة��X���g�^�F�G�vD;�퉱.�h��� }Z_D�ݪ'�M�[��}F���]�%ަ犌P�AW7�G�l":S����E�R*�|P���G����:�bM���ې86@���3<����'�-�@�e�}�r؅���33��*�&,�X�6�U�x�F�W����-*X��n-�&P!�=<�XS��jc�^�sc��H�+�4c�5�B�wyu\���K���}�>�� �<;�1�+�bU��AEZd��3Y�a.�: =�P�CJ�ǝL���O���@��%I��R�|��2�}ص���uʇ#=j�K�1��F�` �|H�D�b_���-IX鍭������t���_،�H�>���.r��ݾ%��S��ף�o�LrQD43K/X���e5䌶�rQ.�D&�ZQT��/z֖�G/'&�E��Z��g��9�ʐ�݆B�|�O���ګ�2
���m��B�i����S]0ز�4�Xf����Sd7��S�3�/�aT)@���Щ�6�}�_Ͽ�NJ�#�gR<4�8h7Ro?`���-c�.c�i�,`!B�B�ҡ���	�&�pqE%�:3+LpՅ�ǩ�b�Ɲ�;~�+��fT�"5;Bc=�[�jf
cB�a����.@_4���}���D� �o<��Mv���J\�h~����	����,7����E�Ay�%��j�Iʥ�w����y�mYmp�,d�$��g�J��-��eE���WC([)д��=��;Qm�CH"��@\8�د���]h����Ի�J+�Q�T����D�|/�V�h�7X�-����GNag!S�Pܤr��C��[
�To�Y۔���]9��\�ʗ�����7��R� "���c�j���w�Ҷ}G ۦa^]���tY�_n�_��E ��3��D��A�z�m{�c�;��[<�+A�a,{��&{H!#8��ʋ�+����*[f�i��e>��Y��{���������]�8����Uh���̺��L�Y�o���DY)+��7R�^���`��E:n���D���K(�K�Hcl{ʥ6�E���:�zO�b:�Z������	�`*��kֈ3��u����KS��❫����(	�LG3��@N�(^���P�/9�jC����U�C�Ƶ���9ogѱm@l'xU�8��-�e�����wz��6�ˢ� ��"�j��7��pi�?`	ˁ��H-���egL<��!s�}�����0M��r7%:wȼT9|ֆ�]��>ESPx}���#C(f��C�hs��)�[����-"@���e.�:�Z_g�]�FS檩���%r��ԁ��e"��޾���9Xi�ڐ^p���8�:7�{Ng�oA�BH��Rڱ�A�"�H����X�LK�Z��s!)��~bMwL�}��]��L����{F80�(D~�e�=O����θ���UT��I�����QP��+^uq�Vn�3�װb����k7��կS���g� �����!DV�O��c�zR,LQ i������z/^�l��7�,�I%?�h�u/~�"arh=y-�`R��O1-��
��p3N�3c�;��&��Н�8��w�5�`�,]d��B��7���W�`5�l"�3m�W값Q {묬�
���VZ[u�m|�q�� @]v�����d��3*��X��j�$�r� F+�չ���j�
����Tzc
7о��I�5=/<X��|����Ʊ9��&C"/"|kJ�[�<���\�}����L��'w�b_��7�9�Q"f��pK���ia�u��,�kH�{�%�Y�w�x���c1�ϧ�s@va�-,��T��)�nu������M�G��&<�S�/�Qrr�s��xk(n{�e�x��|�m���!�WT:톐�����m#�>E�)r"�g�%���m����L�����>�S̤ʊǕ��7 Sȷ��:���"�pǛ�l���?�h'�J��9����S�6�C�m�_47&Z�ݫ8�8�^?�ɥ��K�{�t;u�f	j?vB��`BHކF���$���]gNR�-�蛁�h��n��8����� c�e�M=Y�R�\������Պ���{Vu��4�A':wɑ�I����:^q�D��v��RP�zl:�����&�ж$q�T~�w��ݶՂwC�#���&�YBJ��&��"�lT"�Rc���TI����3(4}��ڹ��p�T���2 ²3�"E��Ucú���麈JD^�,�}�ՂnvQ"��A��}q�?+ۂ��P��ë�4 6t]�[�����\v���!\��nn\	c�v�W@��[�H@�i��Hs2!��=���b�el�+�"[7�����
Vqof��񦦽�����M�A�YO�W�6�Y�[Ï�lLF�p�Ĕ��-ͅ���#B�O��T}WŻmY���R�� M�7��
_�����]�b�����/X�i�8�������I{{��4�2lղ�5c�Sr˦о�t	���)�?aR����']hݨ-'H�;�_��s���I�
sN�99~CRs������>���P����R⑅��E��R.����0-��M�󻮅8F�/��>R����h��I��_]x%�hf0���dR�͍��!��e�dD�JW�n�dv���4�u:R?�`=�'z�]B*k�^n@�5F\��#	E�3K�������n�#�]G�.�q˸_��غ^�/0w&6�^-�l�w�HG�������w�tvLշ����KgȞQCS�=)�亳no�NH3��u�]�ovŖ	PD��\ 4��
��]C�{�ʯ��.J�4�"�E2V4���0�[{�q�,��1��ZE0J��JjW8���Ǻ� ���U��(���v� ��� ��7���0x�!L�t���@f��b���P8������'����� wb���^b?��<Ԣ��r�1>�#C�fluzj�%�11�t�1_���7y4R����g�T/<���$V���Cq1u�d:�5�[a�{m��� C~R�Ƀ*���p@�uq%�Ss�bo��r�~Uc���[p���g;�Q���m3�3�2�I��u�n�a�mKêɊV����j��u;�0����ڜ�&����'�"�5�Az�];�2V�T|`�s�r�}Qy(N>>+!u�;��!��p�|�,�J�(�և�-s�˖���#�IHќ���YY�sw~-��墫�PD҂�C����z@�F�p/�'r�����;Q'���+3�=� ��rG�fmlh?@h�C�(ְ8C����?�⑞���t.��帠�2��ܺ�iY���^@�w8���`Yy��w�)�A��f�$*�s�bf�EC+�.�"D7��lB��7�M��v?�戔���m��!'���`!�jO�'=婝s������n��y.z�5�}!M����$J�i�]`H��~�	�&. ��:���F�)2^-���.Ip6�狿�$��)�]�Q����=�˓ <���L=��+/2�K�c�#Z��Bs�?�̾�'DG��س�A���<{q�˭�l���)Z�������3m|�ȁ
A͵����J ®���̯��m�]v�"�@�,#��(Ë�v�/��TH�E�oA�x=ܞ�c����y7	����@�(Ҿ��]r�S�x�O�Jg�^)�I��M���یF�xP,�H��V�B���x��lٟ��f�"���q�XC<�m��
��~�.�Qfe�qD�#��散O��F�n�L��|�}2B�SS�fM�
qU����Y�����H�R����3$?ṙ�:w��'L�u����앜'#A�ɱ�϶cJ!�Sga��:L(���69����{~)�|8����}X�H�6�̗s3N�uN1E56�����a7�A%�:"ԣ�S_3��+r����L��apV	�/
 @9��q���	���n=�3�t]l�%$���l�Լ�w�A�w����~c������&y2�{�"'� �|d��	���V�Ԑ8�D�_��d:�x�(�-�B0�Y�7����e�Y�_��4Q�A�x�o�ɱ�%�����C��)M��'�
Eٟ����<���i',ƻ~��Βz�/�n69O�r���"�t'7LD�k�Sg��2�X,/D���`�|��m�z�r����h ^Y�{�?���"��11\l��9�i0Z85���0$�T���E��\ԣ����*3�3��2'��o+�5�C���6��P���x�.0��l���:$�4�W�$&�(;�2��U��G_�|l�ͅW՗���x˒�K?qY�����*E7�\|ԱD_����j��̿�����c̬�>���װo��.g�v%)lv�jJ�;"��fa"��.��U1_��`	R�4�����q\V�$���M����r^/$>���t-Ƭ�jAa��?����$����<��^5;�s�׶��I�������NtqU�.�_�6a%�N����so����M�����	��[��:b�QN�f����O�nY9�	�4zS�ζ�0�o��SS�5i�"����r�p���ؔ��ضZ��[<����}�2
��dh���d#���b�ʖ+/u�W��͕^	��{#�jf�3��D,��(m��Z��Q�`��z��c��'zc�i0XS_�:�HJ0��b!V����9�>��+�sr`��
���V�U���Oei���'d����O�9F;�I�ؕ��#V��qU��fd7"l�c�|�޸U�Aը��C)�0��ȱ�e2)���N��
X�`�V���yѪ� ��=:����;�����[*��z̘��DT1ԬQ}�V,��y����BC"�� ��� ����e:)3��&�J��}J��b#��0�����>�"��{�!	-{����0#}6-��!��\p1�~tg��+�ӻd�G�~��,}��8vop���T��ߛ4��6& 4�^��)����f/�`z����k(x���?�J�aLș�����	���8�~,��N֫��t����ǃ쪶�T�ӳ*��HG}4@�ߗ!d١��Bj���Ӻ��IB�Y�*r�9k�Z�:%��w�	�RC:�o�3N���B�/���Y�M�m�OR����6���4{w4�\�v�V녭��[G�&n�y:��ʋg'8��̓�ޑ��%��<r��F�C��{�Q��C�ah����.p�F�sc��k�ucqE+"�8�샘6�n=���1h�-òy�4�3e�0�a#1�x	���q細��P
���n����e=ח&��`~Ь���@b�'	��?�:�7GGs�b1��|#)Cge-p���[e�< �$`�s�U.]%�5.��8T����a����D�)bB��&���{��0�I�F�?�l��[�0�|'�$�[۴c�#��S��XMD�Cޝ/;�X�8�����z��f]I�<��y�n��+�o�^嬳=Ƕ�(zx���c������7��&��D��9��ODiI�sȷ6�%�]�q�di��쯯�j?`&��x��c�Q|�IE�pV$o���H�9$KՀ�8Z�۾v7;��-��V��_.�:�Xi}�3�Qs1<)C���{`�ԝ�\z�L��w�f�W����1��bz!��Ϳ�E_#���<�v����
i���_��	��n��O7�뱋HeqA҅@2c�ҿ@��,�(��ɠ �1&��R�x���o�� }���t�O����C�����ȇ�����1�3�{H5�H��A��y�}��ֻ��Yl�ˀ���ގ��)x��"�!�ۖ��TFe��I6�=8Շ��v��A��Iױ���G��gp��� ��TX%H�jJwu��%�B-z$�X��A�Iʑ-�[��5�n#����(zD���.�m��q��ջx6�k�c]理 HnP�e���GṆ/��f�����I��gD���EA��4�/f�Q��ng���y�j�A�
��ؑ-�0T$�Bg8=�\�6[��$�ncUhs��5�+�8ˎ���~���!�5G���;3I���"ń����jw����ז����޼��~'��#�����xAkx��x����[|��Q7����X����[�p�UN��c���j0�U���!�X��D~���u��,|���=����皩&f�J�9��-�_ �
�������)[�<�ċ<aբ0��?չQMz���� ��	j�(yT/:q�.�rs�_��½���:��2s�/��P_�֌�D�m���$�y 叏�������rq�`陝��8L����K��:	����J�� �C�&�϶ws�/�L�I+Q��)��M����^��	8ԋ�`���T�����|+��fE�쪿2���f����Ľ���� ���C]�Ͳ0ц�S�k�`�y��B��K�mz�H�g��*�������r�D�靈�b�^������PPEȶ̷��ĄVSw��1#�/2|���0ں�i�}���V<��K�v�5I�{ĕ�89��wk���T}����y�e��N�Ҝޞ$QT���'P�Md�n���eS����S�����<ꃔ�,|˒.�Te/� �m��0�}I�@�j�9t��͔U���<��8;�TO�%�8�6K$#�Hgp]7�	�[�,#�S&5�"C�޹�0k��x+Ԉ���,��a�"A�����0u�y.@��k����Cx���� �Q�%�s˱(A
�����]��DfT�����$<��G��r�E��ּۮ�܊&��Mke���V	tBk��w�z���?��!H�9� d�H~��	��l��=]���1ͫ�ꌮ�|�1Y-L-O��wY�*�Ƣ�v|i�nQ� `�*�|��*�jr���j,�i���'OO��3���8,�q�͡_Sz|��M6�d�qH�����V����w1K8Ix���WkjΤ*� q*���%���//c9H=׾�.cL�E��$�L_����Օ!e8�ej�W���FsU�cs����J �n�`@��eC
]Ч����-B]�FY����l�M[T9��{��k!�ʷ`q�n1��;�R�!�q��ٰp�� ���L���ZșYUJ-���T_>��+��bb�q��Ȟ\5���,왚��R�\����޿X���j���t����ñ��129W#�@���׮K�����Z���a�;z[��~At/h��}%�t4%��0��=x�Ù{�I���E���gˤ<�\�� {�Ǔ��G{�a�����g&�[�U�"$���A2�w�  �DW�	��䣲������f�r�-���/��S�
��㛊�G�mdY�}��̅7��?����vİ���d��:��v���G ���Jr^PN�e�G*m"kR0�_���vϗ�N���S^%�֮��Κb�ν[ۆ�q|�����$��^t|�������Dl��jD�K���
��0��̡���s�"�k'񄅶3�]����B
�b*�J)�B6�R9g�����1�}���	E��'A:�� ��V*0�«2��H��:�����W����4�;�)��<�	kN؟[�����45x��ֽ�4��h�
���w
�sΦ�/0{�e��d��e�S^��<�&H�6�<ʒ~����"�w�4ז>T>@�i����b����n�'��`d�d��c���|Xy/Ѻ0顧ih�(k0�����,�@������ �ͥ�j�@��vK&TƜ.�F��i)�T�]s�k�k3UG<�`k%��Qޱ��.pEZ��DE���>n�6l7��X�IΈr�����R*'�dJ|��a,�����I��_�T��7i���nd�XgW�0��s̀��6:�3���i�U��g ��eA`p͆�ﱽZt�\��IL��ð��-���|�;�1yQ�Me�[�E�L73�4r�h��l)��&p��_F`�e�od�����H�cA���.�HXV݉$Iq�&V�ё���2��&&D��B�T���w�g+�_��N����%������hL=A88@Oz���K�S9��������W�I�F�ԍ`�����oñArϢ�K�.���=�,�&�пp�n8n��^Z�n7�O�Eͨ�.��ǣ�E��H��T���m�����(&�KK]SE��6s/��_�=��sݗQ���*r����퍸k�#���T� Zz ͳk~��n�T�
k-�;�.���a���l�g��|�=W�jD�4=Bײ��@�^Hx!}�婷$�;�iE�Y�r�I����x̗�J|l�2e�`jc��[��t�_��6�<��<�B�3�N)���S���g�������?�9���J��g�n����:d��;&
��mb���
-ȩ~\c��Y����� �
� j�C��xkS�c`�b�(�n����۫����w�
�������KȐ/a����v@Xc��v!qmo|F��EU�ai���|	�)���E���6�in�f�5Ps�Ќ�O@(���om���N4�,�{gx�`:�X4��ma��a��<��([�%Hi�^}���@5H屬�mtL������\4�)?M��lD��Y�W�w�2�������|�g9��x�3��4��W@>օ��/�Ȃ��I��	�嘸ag�F厮vl�G)���_;9~<=�k�N��z4�����v�Ü��)�RA�w+%Q+��z�lĬXڝ� a��H�-���Q��i2��`��많j�!ƛy��!�?�=��g1tN�D�98l�-��3J����U_����W�W�A�L��+�au���	�9��'�����+SK�������3��-��^��M8�V�'Ic�B�Uu��\�2��=�~�<�pH��WSw��-0	�g8�b�9��nUpšy����Gp&�r�R���옼�5��z��t�+U��j��I�� ���!b8�\ⲋ��2��w �&�z�	zm��{�8b�#������o��� �m��k�J#���[@�����X�R���Ʈ`Z��{Mi��`��?&���uZ�	�+w�����t�n��(ߐ�>�®���R�4҅�@/�n�a�0]��� h�/S�nD��qF��m�9A.����s��O�αE����j������y�#�G���-��*�B��_��@=[?�Mu�1��M�ܪ���1��죆q#����_�������7kOE�+�a��m��f�7�fPt$� XMJo�.�d��(���"�ڊܾx+~��d�j9�����3�!�o!mj�a��h���Y��c��`.�mmt������t����i�algL\�{5\l��Á�\��<�w0�{�n�ǡ@v��f44+�H��I�C���w oo��+��g�!���H����fZr�k��;{���.�jW���`��NG�mD�ୌ]�2�u���m;mc co���4��ɚ�*�-,1׭ݤ@Ig�hG]*=�_7�.G�ݦ%����Ov�z�j<��XfL�*?�����o�Q��
�TT@:�������U5a���Z6��7��I�q�R]m`+����t��z�ٵ��&2SSk��+�W�n@�
�x���Xeܽ�kpw��@Hrk��X#;14� ��=a}Q8��X���8�����uB��I��Cë,؝����|I�[�
��33�0�[j7u�������N�IGi��䈆;A�[g���̅�Xg:>���`���h��D�Q��8}���Tŏ�xDG��I���?�!-y�P�yC�К@�d������A��S��؛�ڍڄٍ��+p�y����e��G���x��E�P��a-EDŵ��W�茕=�C��{ZI� F�J�Y$�)QZ$T�\#d �������/\��  �3y+���i�@�7{����s�:�*V���f��	F-Ab[��(Is����}��@8�o$b�'շ~/�l�|�	FnT�˘��7���� ��%�Gʫ����H�+2�n���7وkCC_B(B�c1}'�({�k��6 ����L��;�y�]�_�)$��g�o�k��P^"���*8#���Y�����߂��.
�x�G����B.)H�)���*�Q�E�(����+}sl���@J߉��.�I�o?�:t��oO��^�ps��2��I�Xd�Ŀȯ�:5	��a-�Y��Rq�����W�r���pW�-l�lc��ƍ�1|8Sc�ݣ�6��8qv	�>� 4�Bhy(�l���z.�{�v�7|k+e\w���$W��������O�d�J�!Y6[����b��~h�^ބ���P�
\6�9���
0���}p��Qw�<���3��\<�^ �$~�2wa�c���FD\��C�k�D(���<�:?��5���Z�w[7�YQ��`�C�\c+�1k���챀��P~_Q�m���_ۢ�t<��ɋNVr�c���U�[{;��~�Z�w�E�嘜pmb�}�a�3��[�)xx8���؂�ҽ���~�S���(�I�b9���GIE�:��mf�DB,l�[�V�G�Cp��Z.�!l\�.�璤�h#l���.�ёkg(��>���8o7�k�;l+p�3�$�G�RD��I`#+�0�r����l�W�	���J<�����.A�
�AT���_�FoȓT+>���>>�\$6��V�a6��U�^�I�4�G�,��~ �3��>�qR����Ry'��v ����y$�2bm����Q-����9��Ъ��k�'n_1�Ⱥ�+�}c��#ʝ���1,�K%�����%� ���6�$q��������bSr�u��~I�������g����7��*���J��Y�m�;��>y+ߺ(�tzay����hI��o��4��)����/%�78���H Ga)�?P�,���
9�0RO�K��ղ�\�J�
 9�˚6:$~T4���bM/�3R��ޅdL*�b�e�n�<�%�zM�G��+K����^�෹w��SZNk�n�������q��'h%4�_���!��=,�OA��d�Μ���A���S����������?I0ۧ�7���P��%�wn�9(dt̩r������٧&�-��:7�!�0b���
��;1��$��G����������28��cD�O0���JM�iu�/�t��;�g��%��G�Ր��A�ǽ|FϬ�l��}��~G]ajn����c�9(ӈ�M+_���ƶY�s/��Z/_��[zզ�ٺ�К����{8�+v6�Dn}ם�x��J�>��5J�y>�Kz���툲�ŧo�!w�k��Dh4{ cl1�i�Amحj�m_<��e5.	��������@�RW��7�hf�+��/�:awScz�չ{-��
����3�IyZ�����6�FFv�	�L�̞�K���[�6!0�SV�V<�����;�H�>�샷B��UT�6�ޞ@a�dr�F+���E��1«D�w2�'r�Ď'`�`���[�L��NR;g����ܾuu��$�������g�>1���S�{�@hh��9�Z��Q$Α${��Es��#ޔL�ս����
�((��A��S�k#���̣|j'�|��	1y����Ef���^%_�u`��$;�BPK*��T���z0�h(���-�W\vpb�&����S��?\g�5��k�-��hCuH�?CC�۟�m)ܔԘs%C��T�m�n,�L�d��[��I˒~���.�-��<k�S���Ҵ�`*q�5ѵG]�h�rr��S*�!� ��7���"-�SF�9�v���������kǃ>v$��������L����,��W�x�H��=Q-�� kQ�CfC��ʙ����J$����W<�X�O��$Q��-: ��M/�n��X�}��p$0�#�5OI�ke�X�Y�e5Ф��?�?�se������Si	�S���5♳��W/��қe�_ ��R����.
a>t!o=��cf�@� �c5�A�]��ߨ���xI������V�v��UU(f���U��2_o�?*j"�vueY4!�L�
��sI��le�؇qI�dM�X������V�@8}Җe*�B�7��,Q!��;��2��+"V���"�	�#���>N�����rUJs;1�K���w�#ϓI�C�ÙԔ��1&���i����i+�~+��16)az{k���
��
��Dbɺq�T=).�Y,0%M{0�����8��/E'�ѿ��X��RB�.�j����8"�ce��H��=�O��`�QH���.b�C����â�Y��2 ��/s(1f����,�?V��:C�A��2��oi�@�g=�GhߚbJM���Š��i�u�"u�ҁ�X)���]Ļ�����WlM�?����3�N2&dyk�p�-�����}>*m��D�7T(�+[�	r;E\���U�oЎ��M=`�7'jf�ﺨ����d+k��g��V� ܐ�>��u��lnv&pj*�h�яU��Б�sQ���v�U�#H�s�
%��[ 1wx�ҏs�r~ň�4瑋Wb�rO��:�9�T>w�Lk}H,׈}�ը��R�;\��S6cj�S���E���s�.H.3�>����~�p%��F���k|�u}Fu�o��=�S��V�D"Ip�Q
�]�R5�vc��4|8-�V����V��<d���Ɋ�	�WU��NƷlC�KJ�1�h�g�n|�Y;�㐢�.v����U�I Q�86:���	� �N�
E�FN8��T�Bi�U ����L�ME�&��5]�~��r$���f��Gq�D�(W�އI�I�4�'l������t{�eXꍨhZM7,�/5Nъ�C5��J�ҭ8@[�;���eh(o�J���,��>+���W��V�=?L���;�An����)�� i�O��Dk���M��>������&܋�z|`^Q�	4�r@���T>XK�LAB�*�h�3�s�/
�C���_eA��% �Wz��.\z�@!��>s*��C:��S��Uw^g�?��+;���v1��ux4 P��-x�����!��$P9׵s�!x�$*����.b%�W~��Z�t�
���SYQ ��e�\i��!���MX��C�׎� ��}j�.`��o��4�WO��cE�L�Q�+�!@�j@�a�F���:��GuN�,��15�8�<���ep�Dex�ȹ=Dp��~u������e��d��*��@<!��lc5K�}�v��4�TZB@6W�3���
��Д����P��r������)�
�h��{��C-m����w3~]��:�f�A+��=�.�[��� G���ٮh�b�[ǝ{��tv��_�|�r��b���r��f��n�*ah�Ԃ����������<����m|M_����l�l�VPV����Y"o�M��f�b6���}�%<�����$�P4IJ��?hG�/d����c���<9��o�+t� ��:"*�y�����[���Y/EW�������%V�����珥.Ϳ=*K��ַ_���娚=Hq�3C��4�㘬�g�m[7�*�j9o�C֧yJS)��5����s?��_��m'Y�8<��Ѩ�]y�4d-O��I�()��r�~�Fob�����0lXL7�ﲭ�CJ�v��@_�̥lE�h��T����ҨQ�:�m�'��p>�ջ��/���*�ɽk��*)���;����m��)���`�,�$+~i�zSB��܀t�qd�*���::(*I<�ХÝ���BF9�_���Zo�Hz8O�K<���O�OS���	kGJ$���[9j�a���x)��TZ�­� ���
�v�^67گ����w\�����]-�/���Nr�px�(��US>ʠ�'B��{[�<؟y�J�����.�1О2��%0�/ݒ��/�3���LeC�=�~����k�A�D?KǷp���S��Ȗ�sBJ�Y�-��Mv|Z�>	���W��\NL��ǘ9�el��� 5:�e��㫍(+�h���́ i���0i��f���Z�=�m�E�m�k��~�cq"�*kIJ6�����_ �u�
�����AG����f=<���?�x�����U����Ct+{l�������8V4�� 'WJ��N��4m��ț � c�ޅ�9����B��M'9oRf��o#_,?Q�_����v'�=�pR�����|C�	G�_���!
V8U4s�5��:� �D>��pG���B���f̸���/]m��͙��].��)_�ҥ�-N�E�O=�_�"͇���LoӍ���Mc�;[����
��&��h��^|[�bU\������n�	�R��n1p��öz�ޒ2�)�&D��� ����&�Jw&�������>@����ڕiNɂ�va�?\j��z��mr\:�鴺 ��K@��^�U��j�z��Ӷ�ޅ�-������K�eݰ�R�;��~��2��эS�՞��3��hW����
ʃ���qu�_\��#�������.�ߩ�yK�n\��3ޕ�<�	�i�`����\���ʌk\v�rȌO����ais����\�f!k�z^�m��HI{�߲܍�X�O�:dj/�Y��'�/�OB��Ɍ%��)*}�H^�u��jz�&:xgĔ2�D��MS�];BZ�b>g���+��yT�G!�����=�;�bϊ52����k�#,�).0S�t�
��l�5f��,c_��5I��Y���J6�7�C5dQ{�":;^�s�C��Q�_7)��Ȗ�Ǎ\��\�2W�(���3��=�m]0��<	tT�;������Һ���P��rn u�h��g��:A9g��+��)+�-Р��;�<'�DWc,�j�r��tf�ê%#�f���W��R"S�e����o�ql�" �t�B�K����}~��f�2m�5fIy��Lp*�U{��K����0�]��W�`�0��(�[x�e�+.�_��P�����_0Y��';�����9Ռr��NZ��1��Y\�wm�"PXg	N��9?��	��UVxs��k�Z���"W�|R���r뵠��<k|��|�A�eB���Dv1�qL� �����q�a��R��jC�2fP�&�=sT&��}��%Iy��o����ޟ�{�n��W��Q�ߘ��;�_{�;UE>^���@�eТ��}�]b������S�������9�^�4�;4�t�{��^�O��;l?p�톂��4"��(���{D8���������=�Z�1��c4Ċ'��-��Tw�fM���%���u��t I?��L�Rw{jbz�U�G�R���.��� T���ou���R;���YG#�ô�Ř�)w��
{��N���4Dۨ�$FCSl�e�v;���ϐh�odUg�"�$W�����N�.���Dd�l~�Yl�'�#
�C����;ɺ�1�J:�U߈�Ra�<
�葺w�qǂ� G�c�2�ϫ��I��s�'>��+(X�0���|�f��e@?"-y�BO�������
�0� U+O:��("��5���M	�����nX��ymTĭޞ��[�8����[5fP�=�nΉp��I��o�Y=3��*���$�ͿEsp��:���]�Y/��X�L]B�� �W�&�g/WM����I�<�O��N���QI�흍�0%���d>�:t��1���>� �,\��ĜL,���3���Y������(Vg�W!��<1��h��U���[���1���D�(�>���*�n83��½���.v��ŏ�|a����6�.���R��8�Ol�hR�!C��	���:�cD~2׽r^�e�2Z�#�SN���]�ll��?�3��(����pO RlQ����KqBaA/v�+K�n���Iɺ�K�`��!S7Oa�����K�&2���y<�3��t;a�%wֺ��k��r�����qyK�\���Y�Ȍ�L�J���R��nH�)nA����j.��	���L(��D_UbI����b$���!9�8'��ߤl�S���8��a��h>�V��Wߊ��� <WE�g'�L�	��WC�|TŨk���͑�ī�[q-�qJn���S6:��Ǯ�D���>/�F�J�-�%9�湫�J�7Uk�qmKyA6�:[�P�ξ�Lma����V�V�&��Q���(�gX���e����3wE	)9�t�&�AZA�MU�!��@�[���R_*�;>�+�o�j�z��5��M�%�����y@�?�>�Dc�����Xק�o�pW�[^B?�+�O"Ę��&qy��c��٢V����������,j�)�;j=�����:�:�P�!H9���E��]�A�FuvxYW�':���c�Ǥ�2�  �;^ȕ���&��+(N�6�	��^�k�r�X�G>�ݔ���+�dMh�[�%��n�KYΕA5|n��!, �$'��|V֙?����*sC^"@�gq�o��I�0�h?������u�S0H�	+�ҵ��\�X����PD�w	p�@�Ym�m���Fh���Y��쭱�?s�Z˰�W+\S.�R���4��a��;<�u�˜Rn�Bf���X|vA�jЋ�K�5@ʫ�	�Wf_��E�pd!^ݦ��sU�W��w�3W��e�!����U�6W���C���!��ad�����%�<�;�<��WOE��]$�b����sRe�FL,t�\V�b'��+^��P�Z���d���|1#����栤�v���n��������CG��~U�K"�KK�-�����JgP1���D�/�C�`�����س�8��Q�'\�n��������]Gqu�ѣC?X����:Շ�z��^��w�>)�a�MY��r����X�7#Ϭ�6�w��y+�N�_�p�=<��d��*&w��)ۚ���L �����Z$:[�3�f\�0
�!�n��΀|ڿ��D�1T�F�9��pZ�6� �v�0�'>�=�V��~��.u5h��Wr�]���p��mA��o���n y�p����QTl��g��Q�/�3e�W�{�кau�a��w�ܞ�9�7#�
ԯ�3Do�{�P��xW؍�K�G�c�oi0�+�% ��AQ�0�����AL��G%����WuW��vd8�,O��yJ?�;�Z� �]b�,�z��^�pM���7İY���H��C�̨� �?K��l���L��
��Z7�CA�d���*�dq!~~)pc�[9���7=��Ì�@��53SY�a#���B�\���g=����k~�EC
-��d���S�������sF_�h�@ \ì�:}�;���=s��9L����K�i��C���6a;[N_�Ǧ��@4Zo=�u�80�(HnZ��`L*�I�����m0Е}��O�[��E�7����b���b��mqD"��i����rAbȝ�:i��-b���ژ�h�C��a9�+y�Wq�� 3>o�Eoͥ@� %��כ-��o�7Ny(���B��?�s���8iT�k)4d��)
��˻�����g$~�b���i��L��s�����w��?2ޞ�ׯ�g�>�֜T���N�ҽq�t�S�ݰzk>pt���9�8l�m	���b&H.����/t��G�r��L��V�.�^#i��R�w!��_Ӥ�_$�����hʮ�^Q�ِ�8��?����L���&Y5�0̔xψ�=��㧺(1�hL��mŘ�3�f����/�u!��<g7R��;���X$ s��]&���bT�������%��[��9�i��0��@Ǆ[���%Kwf���c�$���1eMᕐ�α�m\J�R@������`� 
�(��5~|��w��7f�]��1���;�f�����E?`��u��$z����I�j���+�lh޻����(7t�b�4��Sh`��'Nb�rSC��{�Y��P�6��Ф�8.޽/��6:k	I�/]�[׭j�X���2�1�4L�ѹ�6��ӟ�p�<���<�P�2��'u������-�)�"��� ~	�݃��*�l���@����X�5buج�^�lN4���b�����X�r����9!�*�(���O��S?��Q�����2���ND�J�,����6�N����xm$��rN�kM��B��O��bX��ȩ����0��3��)}��@��,S�:�[�'F@��i�^.����S�ϩ��SfH�����@���ķk��0	r\�g�ɔ���J��o5��N�����	Ӻc��ş������>�_x��v/����49�{���ى�L�9���
ψ˛\�B[�z EС�������R�;��<�7�������G���c�JĮ7M-�->p�N�Kh�N�21�I��L^'�w�\sF,����� ��v V.4Iy�F/��j3��ւ��vl7#���}�g���L5�'���4H��ߤfw�{�cܫ�+�}��f��z�������3��+������1in>��DZ2����xd����$gb���@��Z��FcHɰ;t7&�z=^�l6bk�(�\'\[�,��WKYcq�cm3[|�A�������%~�-j7�����n��,$Dj,������{�Y!�����������#�s8��JEW�h4T���Dy��J�9��-FZz�N(�bq�?N[`�	zԲ	��[�a����O0H��K�VgU��W8^���/��T�gЀr!wFq)<��ǜ,ꮄU2�G��^>��3Q��Wm����g�Bc5�x�Z��+�ф���������t{Ƿ"w�<����+�,���M�w=? ���@�}�xIm�]�z�WU�y�v��H�(�V����ֈ���e"'(�����vU���a[��mK�!/j�,���Os�E��Mŀh�;#�$5�����`+w����-� ؎�Q{�f��x��G(��$)-$��Vկ��đ7�7��������q���+$�p7��LљQ��K���*���	��Yͼ`�qS�K��t�~���f�)r��%R��TX��{t���� �Yc��a �b|P��q�����|�e*@���$uG���{ަH$v���C�8�y��zQ;��k�B&�� �D�B -�=�� N���xޯsJ9�E���y���ԼQ�&7��r{��DY07h�⑉�w�A��*ݳҷ˚d�<�a?;�G��gyX̸-1�ˏ������i�>�����j������{�g;0�p��/4u��؆��T�]h���G8�
�y+���HU�=\�/�4��E�I����=��c,�A���9�J]'c\�܉�|$����ES����� M][g��ndXY�<;:�����L�ޖ���@�Lh��]m�ܵ��a'9���ץ�i稒�4����t�߬U����b�ؙ�����W��[��A���z��m��͡l��!�P&� T�s�t	e�pb̷�����|+�b��$6���\!;/��Wv��,3T.���s��݊@�r�>I�z��b�Ц>{�H�N�@]�){sv;TT���e�����˓b3��ޔ50Dh�%J|��9z:p�R8l6�|���$�K��8���SW��������+J��*�	�D.�f"��kB)ґ�3�7KI�����P���Gd�iOT�4���&XK�ND�]�Wp|.I�p������ˁ��.*uK)2���M��Ү�OV`���*�ah�;)6R���2��2r�~�ze�};� ��.�6�\���=���Np*4;lL�P����@�j��D���W��\(����>�ǽ���`@��"�H����ȗ�� |oGPd@H� �+,r���ĉ:�p��d�M��x���`��Ұnwޡ �y H�d�ژ"걊�3J��I%A�P�I�.Q��\{����c������bu��R��U\�hR�sS��'�B��)l���n2?P^��o�b·��9�?��tWi��:�F��a���9��*�M��x��M�G�d�/����e�+����ˬ' ;�m5�,�jL��,zz2&��	�6���Jw賶�WL'���5r���p]��ʬd�i��v�r��Y3�(�l�����b��a�$��{�ȯ.��� �����ߣw��g��]��N���E���Y��V��"�~�> ?A��e'k[0hq��VV����J	�
ds��~:�*B�]s	&�D���Q�Cx�EۥLheF�sV�1v�[ ���tNuAa��o���"��q����i�(̫UK�*?-�Hh�T�ꏠ�-|�2�ld��%�A��}%� \H<V��~���AZ/�bCf쯠�����ܕ�`x�M6��>L��W ��'�͈}���4>��������4�)b���Y��(��ܢ�WW�+Bo��6�^Z��Z�D�uo_$�97\0JI��3`��Ƿ|<�sqot�������щPkh�H��h��-����y��y�{'�.\͑�$���;,-_6+�g��MN�*\�#Ma��wU��[R�ʚ.�b���27���&m�-����=���$EK�������	�>�j]�CC��q&4�Q��|ʎ-BL�Ip�˷�^���˸���%P�����<e���f\L��\�&��#���S�;
��T���^�y��v�S��x<�Ă���k����dǳG��sZ��ֿtȑ&9r�A�y��6�?Ʈ��d	4��}y�����T�M�I!�L����	���T�ω}tʫ0�xࡔ��ʺ�K~�n/�6у�ʷ��p�a�����|R�@Mͻi�����~9��t=(i���xW4T3r�l�8hhGZ�Z����m�8-\�f'.�$�\�+{��pT�,�yn����:��|t]�&k�}}c��H7I7ܴ:�#A�q�g���TvY1�VG��v)4��]�L����FX_��������Bc/�����p��hb01�^
�`��0�k��pl�L�R����IK�������*~�»�
r��t�*t��
8�T�h	Z�C�(�?Rd�K?�z����z!��i��+�D��@�\g���W#:��B[����X �����$s|��vج��Yٞ1
E��F���fء6�����j��9����~R�Ց�w���]����w����	L#TrvȕR�!����q#3�J=��(���������p�W*�ol��qrm
s�'�S̥Ǒֱ��c��>��L6ٮ�>on�AJKD-$���A����QA@��vg��ߜ���88m0S��~G.j1�Y3�	_/v�9D�@��LL�ڄ�|�x&�����Lg�1�<B1O?A�lٗ���G�-Oa��-�%qF�������x�/��ւ�=���3v��;9X��M�Ñ�݃!2�!�v[&�zSq�|˱C�xtr"��V8��UuT]dĀr+�i��&�Thc���b��%�J��1#�S�R����)t؋��N�@���z��ʮ�f�C6�E���P9�h8����9_w���#��sa?�h�e��HҊ�}F>�T�
u��Dd��H9��i�gq�6�V+(�U_���Hk9�G��*�q&�P+�pq��������R͒1S~���Zu��ɶ�B�Sl{yM
UvK�Wá�⬅���)�T(��S���\���P]6��X�x�֡S[�#�5Q XnQ��y�2�0����2���ᄍ6/`�k����x��	�����*�z���@�rfZ��gT���+[2Ӿ�m����j����ۤxQm������T��W���gy� ϯ�X'8J#;�.��)9���^��mj87����t<�8	%MS.��J��ZЃ�����v�����RHo����W�<��,�4�S�g(l�Fh�SD�_B���Q�>���Y�g�)G��1��4*<t^E���d�A�`C�SS����m��Ċk~.�,C�ཀྵ��Ҽ�ns�H�<$u%�,��y.7�2�w#������'+�2#���}�Y3٪{����G��N6Z�^� ��,���冯��k�f@xɄ>�s�GNj3��U�3e��:�S�|uQD[	�:��K�����M�����m3�1ݾ1�ɲ�#uҙp��C�5]�C)?��v���X=�;oHq�p K����6��X���[��[	4�i�O�p��/{��NOϛ 8\pN��یg�4>��[C�P�]+!�B���/Аگ�{z^1;�2�`a����xx[�g�q����Ak3�I�'U��o���3&�Ǯ�4��D�=Nͼ���C"U�����nW)�l�6��Xi�r �� d��ONE��P���eȌa̒*|���)�N8�ʈ7M�ל<omj��W�.'mi�*?�޸���Fڠ(IS��f�/���ֹ��#��왪r�7�>�Y�1s�y`��s{��Gy� ��Sف,z�Cj�EBΫ���i�_�Ȭ�u�p�ȣ+l�=h��C�a��]$���d� ���7.\k��{Λ`-�߼pq�a�K�\�C
�'���gN����<$�G3�-���`ʼ+���Ec�6���oW��+3�D+�{3vkt����$��|mezk���6���>;}�j�7~]��1�����H�x���^��E����[��L��_	���+�h�!8$+;��֖rA�:�dYl��#vֽP�w��2�y��Z�u�^�(�L��&�~Z_�a�82c����T��N��|�C�+���y���Ԙ<HM��;�Ed1�S|\��֑70d��/s�jf�.H19\]Q�}ԣ�]la鉓;Zs�.�:M3l�^�^�[ A���!��1�o+�-Z�V����� �#EvL�0�Ix����F_�,��,����E1�&E��[�^�����Dd��M�b��y�����.�<��)g>�N�f�oQ�7�v4P_��ڠ XF�F� �yY��6q���n��+w����RY�����ߕ�W9�?]���S����Č���_!Y�� )ZMFV��6t�XB�Pi�N߲6ب�߃��u$��*��u�"@�!>/�1�Z� 7��0�M;?}��@I���l�E��8�u� ��Z�m��z��)+�� ��Tw���'�W�#.[�<�Zb�����9do8~��ʹ��c�Vj�_a���w� ��ɨ�h>�إ�7�t��(?s x��t���o(�@�����uAX�2�cf^7�~Y'��G�Q�bV�Q���"+���w�9���U�e�S4�]�)�Ia�'E��z�����v��"n�_jRje%�B��W���q �8w�?���=��}|BӅ��$d�sa������4T���:�h��\Va�0�����k<'qTJ���2?�bP� $�� ���ͮ�iˊ�l�>
���^M��?�0�%�Z�6���6�� �O�,B��~)�F_�#���u�R�Ű����u�	���>$�!�z��S}�f�y.`����(+��+�i�Zi�+&��Ԃl�ĔH!�9%�.
Q���~یJ����ܩ?\�� Ȍ�sU"x�������]B0*TZK�x,�FT��v���j�g1aق̗���!�v���y*l�q����^5��7�,�5���V/���}0D���G\�e0o���N���#PߋLp�mL��I�"���Yw���I���:z�Vڠ�zy�qK�L|������ǰo���)ե�<
�V>�v�q)�Ю���5.�i��d���&�W��� 1[��qr��Ⱥ�{�w��Q�;��F|��Q��޳�����ܖ'��]��8�_vs~45:"~ʋ��}��u�"�KzCj��w1u r6��c	r�S�˻z?�S&��4jc�wHb�s��z��H>k�2��4�fz���SĲ��jI:�=x�4I�"�1��!˷hat:��_���(��S"�DcFc�������&�Op_�n��\3)���[K6�v���`b���`P�>��=v���T�	����T_]��r�\��,��@~����(����$B&��@r�֬���Fեw�ii���������-�;�8o��.A�]����%�]Z�[�Z,wӖ��������B�7�^8L��`s�$�j�5����Ig�J�2��h���,C���W`���Ԥ���0;+�崓ﰝ�he&�������8�swPP�J���gϟ��#mdue7i���G"��	ax��׈kj�̧6���w�-}]9#�m9��̶ˠ0�11�y�	����%�H/W��z���Č�.�~�
�`>)6o���N�����ǫ|�W	��?�-T��c���p^S�5��G��"�4���[�x܆�����q�?�ћ�J�<���4����(|�O;K$���[����O��R1̮'�f�w��s�����Zsߔt��o�� -�J�t'{�:���}j͐`[!c���_��g��O%�^�i����Rb8	}.�/޷�U�3��0���mp�<�pM�
�$�q��ó��L��q���ܬֽek2>��E�<�ˤ�t]\\��<Ey��s;"�1o噋�
7%}M9j�G!^�(��e����G�}|-����W�o{�x�����X~`�|HS\2j��Ьm�\qOJ�K00A��pR�s�s�a��xj�èp���4��g���>��l���,pj����m d���'~[|`Z)\ΗV��E�,��.豝 u }[�r�>����mP��P�ݨ& -Đ^G��m��o�xI�n�t��H`F@e���[I�w���Y;]p�xg\9��u��#���")č��mX0
~B�M2�d"����P���I�N�ԭ���R������:J�xd��J��M*Da�n4���n��;Zz[�<���` v��,�o�MR$�OO����9�p�&��ϋ)'��}N2���d:�$�j@�s;�yu�g[��+����b�ղB�	�\�,� ^���s`�d�xG�;�Ф��(T~��o������b�
g�Z��"ǿςe�S���b0Aw��B����{�":�7�/���߰m�u�+���q=v���>L�?G���)�<��N���D��$Y�,*Z�Z삥qñX�=r��`�!dW�X�������ꇱ#�c����vȯ(�*��/���^P'j<����8�#c�q�*q��>�G>̭U��G�ŀƊ��Zw#�,5j~�J�P�r��%2*��f�[����r̤�f�Ҋ�xd�`��>�kS����=�\�f%��C�ڤ����'��؂#�e ���7k9	���I�U�J�%����q�� �Y?1�q,̊`�x���ڗh����,�������jl���]���tW���t��g8THQ�5q \G\�Z�v��Wx	�4^\7�`���I{��d_��h�X�@�fA5�}��p�	k��*�jO�-�-.i�M�/����{��X��>�K�	��;T��(�tԴ!��[d�ӏ@��������,�G<�p�l���K��	��Ob�֔��d�ʳ��P!��F����0�C$w1��|Q����C�m�t�Ƞ�V�Ͽ[?@Ԛ������Ϧ�<�=9I�ҵ��s䧭��E?����F�j��o��"��0��U�l1җ���զr���b3xq���'����9� �����IHP�����5:��n�v�^���4���tg����Q}��گKț�b9���"a�b_.���B��-���x����b�{[E����gz>�H���,nq�	Gjyb���6��,᩹��ǘ�?�΃�xu�և�-���=j'���{XO�}ߠ%���Mic�R�%��9�����K#,�����7�M����h��c��YM�)���������X!��;il��>;���d�mf������у
PDV�l���~W�@���nP�p�X��� k�n& z��u���P*�i�.<`�-p�ݍ�Q�)�G-�Zd۬$c��()p��&{���
y���R�\]����K�9�#�c$"�c �&�^Ŧ@5x>!g��x臈�e�-����*��Y.���Ö-���f-=�T��*��qA�2Z&q��g�����A)��,
�U�Я?�S�ȠdE��R�ZH~�z���'p?NF\�c\l�`󡴧������8��N�u����rV��%�