��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&�O�}>Yo����i_�s�tu0�[%��#���E�&R���ԗq���)H�o����Lk���wk�1��0W�}]&!K4Ú��\Z1�9��F�"��&̯���=8��ڔW�9	,"#�otlA��^η�5ٰ�F�$���j��06ňF.�hF��4�@�R��H���QX��q����d" ���4|{�*ZvG��t�Ey	�n�=a��4sp�K�H���-�����v)>ش�4Eɫ��e�)� ��n��$::@]G����U���ҳ.�X	;F`���;ߑp
F�<���5�%ZI��d\r�DRʹ�-�C�2
�b{.'���2`�~LD�o$h���h�`eK�;���Je6`��\�t�>L�d��zq����l^@��{=���dd�҂&��h���ʼ-�Y�(_Bo�5+R�K'ҙ�,�΃m��t2�yC���)�?]q?I�ЃW�R0��T�O ��2�Z���g�+g�1'��`�<�A3�Gkiw�CGEw*:Myh�a���3����Q����!�cl>��r��~���j����w��cP�;�/�׀%Z��Ή^���=�q֭�=��FFvb���i�f��Z�� M�䩇�v$�-�.�!�{�_SU����ix�ɿ�	ޒ%+hB��)���D����@7n-��z���Yn3��E��������ˀBr�࡮��z�Q�3������07m/`2`����`Ԣ����	�J�ؐ�5'SX�mv�X+.�a�Q���*#��tY�ZMa��H���.L� Y���2S�$�q��Fm��\��n�ӏ�F���|y�5��!�]W����g�T�I��+�'|y�)�[R�)��M�$�����ΤD����������h�	x�$Q�õ��X4�l���p�]��f�X���;�_�c�8����c�H�6,�R �9h�Q�sI����}uk�;XA�j@�u��{A�/�H�B�Z\8s/���B
�4l�&�ifh���d�{kXą3j�3ƻm8��+�^��w�� �nyح���B3�Ex��GB�[n^�$9��h�.(�07ְ�!%��]3���)�-��]g�g�~)�����=tX���H�j6>��'R�7�δ{�lW��	��Ie@c�P�pM1lR�gvJ�E֔�q[�{g�L��%�
rb��t@.��r��ۤ�NP���n�����^MR1^ '�D��������+'!������\�����C�� ��@�v�wZ]�a�3�*,�S�N�<�Q��|?��)D�5X�A�B�=���Sa�a��N�O�����kԑ\�P6=#bQ&'1ewuV��^XP;*�S�^�4"O]�Σ��c����㒝e�W�y��ZQd��7��f�|���W��d��h�D ����Ҩ��
lfV�*gZ�#J�Wž��O�Klt�������o�]C:@���iP���C���$֔�k�Z}c����_$��Bn�X�aT��i�j1�F?y����3ʣ�Ge���+b�(F�@5��V��~�[6�Џ�j�`Sz��~ބ��2쏻HT,Q�L�U���yҊ����� J.�LaEK)����6U�B���=�/����Vٿqd�"��}d����9�'�s�)�ԃL2r_ڲ>Ro����]����-��B��AH��V���?&�QԮ� �P��͹���-�6JA��\��BA�b���"��B��M0�o�B�Ed9Ϩw˖���h�h�����w�ՙ���
i��"�ʣ���o����0[��8�S�G���n��l��~�EO�Ǐ�[��5��H�q��T�;�0�������㸻���<d	1����濊_:�|��d���VH�8��B|~�u��J��{��?��}����xG)8�ÁY��Ś���u6`:��@����4Б���b��w��ꄠ�a��!�a��"�<z������|>N�'�K����+3n�X���?��Wt<_]K��=���
�6��8�%�[����M#���fcN0OMt���r:O�}T�Ei@N��i�{Vչ������N �p7�JH�����g%��Sh�:�����0��V���e��gb�f��?#�VT}��qJT����{ p�#$cl3Tx�~&���o��Ws���Nd�P$�x@���a�y���站�r�ǽ���#z���Q	�O�s#@��d��[*��+���,6,M�K�����9Z&��7�2� z�a�Q�F��vMFK��G���uk'b�*tǺ���E�*�K����u�O�s�CT����e+�LtL����^���\���	��ᛝQqQ�rY���=�j��\,�ܠ&S?���I�E��%��6'� )��D��0,��~%�|������ng.1;5��u���g��w�I��F
���˙@�	�~g]�-y0���@
<-�#O'�|K�hH��\�Q6~s��S����LJ+\�|�-�F�C�2qf�p�{R��Q<*|�2������ �Q/s"=�B6ح�L��Ic�-��RR�,_�{.C<�:S�wsFs�3D~��Z������V,,�:��]����f������y�׈�C5]?|��\���1��sC4��;.�+�6��x���Z	�G�WZxU�\%XC{E3gd�����5�X�7�Fr1��
��kDn�gll@�8�cG&�Ok�  �-]4+�14e��������><�f�ҡ�^\�_%�x�q1-��4�!������#�,�����C̴���p���{b�SoW�E�+}J� ����Nk�p���-%�v��%�0�R���/�G��[j��ڄ+��<r)�l%�6܇�6��6B�y,/&E� �0�u���ji��A�0����3;�O)�%��_K�u��ij�ӭ/G\�sl��7\�t�Ku~��Iv�K2���=�[H�1P�ܘ�7�����"�nB�Ȅ�yH��!���t[��\%��O��h^�s,8�N��[���5ɖR)����~FT=7[�G=���U~��<a�I�K�.�	�,��b�8��rG�Mpv�4]P�pqg��8\0j���tqiJ��؄P��|4J=g.�u|+�u+B����O*)�*g1�yBh�M�>�O8�SB����4!���[��UӦR*{J��x+_>��9��|��P}�ݽB��0�=��uOgȿ��@���渐��N)�W�#2\3��^%'���J�ū�R��T�Pm��Yđ[x'���ΰJ���dR����
|u�-q�[��IC��c�W�[c���8"aS�.l`J�v�S9+.R�*\�az�}Nt�-��6]2E��l� ¨�2&�Cc�ᆠC�4�/I(P#��Qdwws�P<[#�n���c�ܪ@ľW��m���(y|�9�6���^�翤e�m����3?�12I���o;���r�������zԓ)Kj��j�h?����i��P]�mT�M�36�Y¢�!��T�;6���@�x��C��n�H�rnq�]zP �"��L��R7i+u�z���Z6�
�f3�>�6�b��@ Ft�WJ��6�Z��qDw��,�D�3M��%ǀ��""�Z�F]��(/��;	D��z�N0 N�`@�,@1�C$|le�vP�-�xOs�`����N�j��5R��8H�/5"��;��'�x��hR-�ҕe���Ap?�����5P� Qk���'K�g �����ġ9y�`"pX2U9�D��b�/��xg�
��<�C`�,)f�.	W@	11�g�q�4��4�]��Ň����L�:Z!�;U�Ꮄ��|��3����{��>K�a�0�ҩI^��?IS�DS)jvƁQ�:�U���Ȱ�;��>Cy+��xDFe.3�^���Pg�סn1-�b�!�Y-p�~	�a@�o0�Ix���'�ڔ����"�1�����5qX�9�g>~ga�hFR��
�P-Y��I�L��[h4p_�[п'�^nD�.�]�6����G�%�kl��y>��$��P�R���m�w���kD1�rEɥ&��{`��+漲?`S`�i��I�����W�t�صQ/rS�K�j��6�q5�h't��I��$ۓ�D� �� ϓ7�,�>�Z�h�#�F�g[.�0���� ���N'V�6��b�xg�% R�,���[�Q�c^��8n�o
���T��8��P�^M�"�V�R�;1�/ڔgL�	�,�)x%�?�������R�D������S|'����{�ǹ&�TQZ$6g=%����[
�g(���R����>ۃɦXWq�a9�	6�fM2�z���[!%�d܆��8��cY(ς_�Hc��B���K��BU^��������"G��R�<��<�|���[E&X˸Cv���1���E�$�ė`�"$9�5���_tٟ�G!(�>�a6���]�>�Q�;�m�����.����&n,�Q?J��Ý`�`	���|�q�((,s��M�}�P�9E��z��Ҩ��Įu/Ҽ�4�8��$]|�d��Z����4	~��p����ۊ��u=��s��+��D<��&�X5YfT���~ñ<u�1A��)��	���n%�����P�����g��-Q���C{"���ީ�����,� ��S��`�q�/{+-���u@�>
�f��r|�|g(�ã����`�ā�L��*yE�Ƅ���Oխ��%\�9hF����YrgI ����~����sh/�I��.����	B�g�
��Do�T��x�4�"�����n�����ߥ�[:x�8g�8K�4���jf>���0� �c�J%�	�]�e�a��܃�$,�g`�wE�i�:~2ũo����(ӜR��;���d(�L�t0z������ɬ$�s��������,�;49n���trͯYNՀ�?�/h=�w��X���������-F�y@�u8�~P����yyp���j~���[�H����f̱���*�h�nt �V-�	���9�ׄf)�6Y	νU����@�% ~/���K���1�R�{jF0DQz�]0�M9�k���9�����b�~J	_<}!<gz��^g�p͎��-0W&w)R(H���p�m�3-�g�����~~�~��cU1E�M���x��K�a��N*��^��zƙl>���Zx�o�R����|W�-U�Ο�<5���C���D|����ހ���&M�Q�Q����u��� ��^�6�/aW��R9+G=�����Z��*���e���!��@��M9�Y��&գ���$� ���˔��M#��2��)얩��[��H�yc����������6�W=yC)"�a��s�F��hsd�h�ZD{�LR��I��2� "B�]'������#X5+�����zk�[ݷ�-�	�� 
��x�]��TL�ױ�>�f�Ҧ���w]�aY0B���*� �j܂�p[�R�!x��kJ�7����H'�ꎜZ��O�܅��SY5�ʠ��j{�f�����;[1>����~#�u��Ӱ]����
E���4;]����9�!��[�x���h)ՃWrYp�!�S`�zF�$�=�,{E���
�v҄sa���Ļ�������a���ڟ!E�9\5�ɡq�;�����f��SƬ�Vs�Ld�E�V�N��x��$;�����up>��#i��S%	6Ȃ6W2�;VS��5�XkQ|�\~��_��eߟۿ8k%/ۿVڎ���_���S�x~d�b��x���E�YHSL
�7g�g����1+_�hoA�s��*�g����r��T��S�u�Tk���u�� G��d2�1��~�(�Q-7�Ӭ#wD�.��3)ըٖ84?�xm����o3�{��E�D�>p-��p�"���/C�)J4;�W�z'�>����!F�-EF��.l5��<�h�+j#�[��I%ou%;�a���j�T�I �c�[���O��s���-"�B�&"���P��ݷ�i#AIV"L�cX��N�]��򏮛1R,y7�"р����G���ܢJ��p�_�[qy,�E���a�CD3C�(J���f�B���tڰ	�X㺎1U�X���`�p1�N�r5"�j����tFr�Y�;F�|��,s9�&��~���z�5�ӡ�n�nPNߴRt�p�M-2�9��$Tph=еjB��9��^Yt�����Vz�Zzd6�����"�e�S�^�e!J�p�q1u���ԃS�LY��Ƞ��ݘ&�E�3��(͆4\����b*C�:Z�N�����A�I$l	�����L�����uۛ�nཏ����B0}�U3'NA�0�Ek�Ҫz9N�4��ҁѰ�g�`dEJ�p��F��=&:E_!�u	����י�
�L��gb1��I�j�=��R�U�6 4�u�|�>g4./�%�T����r�t�N��m���n��$�}Tɴe�?��,N����K� �N�/�tc=g'Ǌ��g�ߣ�VFp��U�w����驦C��0M;!w�kV��6*�2�N��ԡz�1,CHj�t�%��b;\���*y���~�(�"6$�����B��KH_��q�8�)B���
�@�+��^JQa�v:��T�u���;��e_,.��Ll�aK٨<Y7���'	�m��wL���=�MeB����l�'��4h��vܥ���D��͉J{�Y�q�f�}ރ;Ӓ��V�)ɋ"?�gS��(��X�\��l-��}�C��3�K����!�s�fsЕg��)��@��7�ex^��,K	�6ލt�nE����h!���[�L/�{�>�2�]�e�Q_��!!�B�WC��uqm��On����L��΁INDA��˫5?U!���L+�9֣����#i�iНgc�ql�ю�����K0�xM ��m��TR�T�1ݩ���۷��'W�25�'���B=�oB�5t�r6��@�/1c�8bJ*�V�h�� ��p����ƿ�0@X���i�Jҟ�k�S��Yx�§jrء�L�:q�>(�&�`����<��֣���ЍP���,�����x=�����q�g����%��In������诰�	�w��8��*a���]�a>�Kr��xz�Iz8�4Kٍ��1@s�	y�%��[I����!��Bh7o�\���7e���Z�[v���+RK�ր��c�,��j�h�w"�!�Ma�Y��l�� 	��K���P��O��6�S�u�
�N�6{�ǂ��B��R���!�I�f�~���V"��r�3�ͦU�?9d}
�/�C9m	Y�m���N����I�|gs��' ����$5W���M�� ��{_1�&�����v�,Ah��s�B�2X
���ag���Ni7�a8ai���Ùj}�[ݨ3}$KLs2B������ܦ���"���^�u��zՋQw"���?J����X���J��E��	a��7�q��A*��nC�I����s#��~d���UGQa��טc�Dd�j[x�N�NrR"�8��� ���^�9;bc��.���_�c�~�fa���8����8 j|�4&Ȍ����\��@��7����1m�W)�C}#�ЈꞖ,9�SP]�'��G�9ײ�B�}*"�5U/<�br]�l����ԁ�Ê5R�^[21T7���o�2����^��⧑X9����ih!�t��t	�z<���q#����"�)������u�h�n<Ǧ�gB�)�,Rӕ6J�����i�h� �Ӣ>�^țN@��C)������t���ɰs�y9�?�O�/[�%�s�f�yoI=��m(aM��Ay����i��S_���8;H���0�W������ۑΣf��4�C���Ɉ�d/����^ޚ��TYT�2/��%��a������#�x��,�w�#QL�`�ee�k-'�$��gRK���B��ؿ��=e��s�@�q'6�W�у��D��,���	mcC���IP̧B3�n�̪�TYԹ���,��a�IT	�9�UwY���l:&3��@�.�������������y&ƟN�%`�K�:��Cܖ�a��/����xk8������E�i�t|�룎�7����@D|6j�yȹ� �#�Lmә�QV���[l~�T���� �l�}9n#�#��m;�l�yw��6��� �����߯L�ܚs����4���һ~ދnR�v�╃�8����0��30�4�}7y>��a>�"�C�c:	���>O��H�{�&���
�[���hqBИ�p�J��]=�;�� @랸a%��R?%l��.(��D�pg�$����w�p2]��y �W@oE%G���s�ާ�JUB����A�N�����ia����x�ę��tc2`oXhl!��}5���L�,&W:odh �a#������X�u��T�*x;�!6���X�QH�l�<Ԯ���{f?�5u�<7QsQ'Ź#rh<�gX�(�+0���&��U����n�T�TO�l��M��\����b���&�[�GHoĭ��.��������s�܅��h^���sh >�q�a��m�j���b�>)Fwh}>�
:�wNn^���DQ��5e���}�C��J?�'�3����vv��ڑf�@���چ=�Y�Nc�_��w�����ıw���6��(�,{� ɳf�UrkZph�`_���?>�A!W��¡��Ry�R)�>� $�gm�����z��ս�r.=k���M�?����V󡨃�>c(Wꎜ֗*\bf�%�goU�{�nY�J�S����s#���<������]�TQE|�
�����d���	��Һ	%�#�y7��R�R���"�a�N�����'��S�="1P�Iw)����m��6��A���3��P�Cg� �O���6PAs�V�,��4�J���k�M��HC|��$Ɉ�_�r22HQ��䧇?�O/�o����d�(��]7[B���f��M�������2�Vȳoq�wUX�b��藭��GU�r�@����0
��#+�%n���y���9ߏ�'����	ĵ�+drGmZ@���<�Ϊ'jjx�OT�����W]J)7w)�Vb��jU�~$שqjC �=Xj�59:G�T���/�N�[��H�U�v3w�N�'Y�3&wj6�<3U6�����ؿ����v"�b�<]�)y�`	YW�5;�����R������$b_��Q�FI}�F��Ue�<��T��< է~H�����5�B����ٺ���i���G�D'k)�Rr�,��魇������"��(����G�o���l�'0�������z�aKO��>�7�����ׁP>����S�z�,zs[���AgMj��q������b2��cj�?-�Mq��T��o���AB]���dG��z�^^����bޖS�nk�8>�`5���()S�@�ʆ�]L�}2�'�n�9��2����Qe��8�墈g������_^Q�n���