��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2ȼ�W��z�V=����d�]�x򑉘�{�	1���ڢӕ��CT�v[��c��0z���X�6b�BJ�+M��1�6Z�:n[����ɿg��Ԑ�U��b(,O���z�Ii��@�9���	j��䯧D���%E�	q��jh���{���g0>j�^��$�|r��uL��r���E����9�й���g?�M�k�$��u1\�[��g)e� �����3�v���d1t���NW�n��Sʦ�ǟ(	�� �[R�h	��y(6�:I�_7ˏ_H���L�*|��4�~�Q�D��Ϝ
��X�Ǒ��"�d�<�k�7C���mє|��*�u(Y^�`ȧ�)z/��j���9:��Ѩ�n�Ѧ�0]���Q�v�x��K0k�E ��N���.��vh���Z�:���;1k��#�DU���z �]>�>4\ȰV��xȏ�&���2񲶳=�*�w(�@u���I���R$9�Rm��­H����3��V�u��ҶY��؅K��%�kc���_�g5,���5�%wuK��6�^�cu�Z!�1�^�,e75Xv�D$N6I���?c
^{�w��u�YH43�5��Z�ll���n�4�>��p�o���[7L��^�����gX�֚���`�E m�5�Јv��܌�ۺ��5��@����X�w�j�h���
���s��/<	>��Tۃ޸���)eKٱb`�X�}��P���qj.O�s*}N e�q��}`"��CG��<c����&l�Br�U6��LP9;�{��	yN�q�h�?�2�tA�LAL�\�+W�,�ܠL�%��Y*�W��HG-�����U�-��׿!��	��V;�M�����5��_J�F3 PV�PF��G����kX����o��t�7y����2 ��@=q����􉭝�N%��#P���T����9C{��f%8P�#�N�K�����g��{@���O�^^�l�	��Xn6K�AK���\��&ڀK����L2�>4�U�����"����Ͼ܌�~h�}I<f�7U=�=3��L:*�0|�U.��u�w�6M�?�������97Ep��-����T� G�OٟgW����mti�Mp9B���)?:Y�m;���5�/{4�݁�.z.����i���c���12"�=~�`��斂�Z�_�D����&�� ���/X������Tsky+�a@�Ѷz��w	�
E#�?�	�@�4���"̡0����P�P���j�t��z�N��q��"��D*���]�-~�8��"�3��Df�W��L��F)�f�O/�1�M4h8����!�Y����Ȧ�t����7"�S"�x�L�NĤ>��A!�\�Ε7dƩs��S��*��?���}�G���9���0SgҚ��8��Sw�&_f׬��k�bt�t{��@�!�i_@f�"aPݸ���D�7�J%����:͠>y�oF�<���Jkm������Q�xY M3w���o��ܗ��q�-*֛9a�?=r����`A �:�Z���<
>F��k��a��YG�}Tq�d73�#�ǜ]����d����6��x{$��Xa�!��< ^������:"��8������+�x̉-���Cgـ��������$|�i �2nƝ�?n����H��j2���}G�]mS�ѹ)��p:��o�5T��|"r� ���P�`�����\�B�T�����T�u�; +����JX�;%�Xn3/�T�J�-`�^I:�V��\)�r����	��>�澴�E�0�)�|����E�Υ}��2�t��T<en@�ĕهT���V�og�>ۈ ��!�`u��V��9�=��e��B�'��S��"j�����w�wR����q�g! �~9v���������s�ޭ�C6���+�k3>�j'Z�u,�0h)��K ��·욪K@r)��^�fJ���4D9�������M�\~Q;�Qg�����k�i@�WzV*��ɦ,���.�f��k�C��~���/J�E���C��im�����ee}� R��D�d�;�c�`̶õ�oN���Ȭ�c<ք�I��w�$�����]]\J��(��~cy�E��"͜b-�;�1�:����YV9���I�mDd�!&��������!������\��c\�g&�s�.r>�m�v��W�P���@���_�>���$C�Q�S#��☛qm�4\�{���̺�'�]��F� ��ڱ�Յ5cG!vN��b3 A��&�|J'�s���W � ��w!|#�p�R����.�HodT^��_��ޕ~)�eϠ,A�� �;�۽�U�D��K�KW��9�֗%��Jދ�iԅEA�'�0㋯U��L~X�i���܀O�	BxF���cߌ�S=��OUL<F�>8��bi�̈́���Y�����.��R�vJݡ���K@�eL ��]ټ�t0ߠ�L8�e�
~F��l���^~��w@0��N�I>v�8и��Ju�8�)��X/�v��DW����
 �N��kmOn����ӽ~�-`^��@B�K.���`�}�d�l.�L��e�k�\��L;�F�H�J�W�:�N�KvD�����O������XnKo�qF.�:B��PF� ���۞!�n.ӈh��]�H�Fw�L���e���p�.�&�W5�4����y&8�(�ՙv�ZI+�����ÄNP���g'&���i�{>��i!6�5�Z��iQ���X��I@�"X6{��J�7�S��?2���c"����m
O �4�@v��$�[y�vIs�y��mH�f[� ��(�ݚX"膻P#��ir���:mo!H%%^Z�Q�F��a͚8ҹM_�/j��F��/����q��0!���O�����y� U�R�K>1�ajz�a��� ̪(?�gk|ƭ�N�{����� NJ�3e�o����9����QE���p)��xSd\����§���G��Zp��˨�H��g��!EF��B֮�Ssv��ͦ8OsС��6o�#�4�",�|����z�jY����b����76��M}��m
��@?#��f6��6����e�iw��r󉙵S6����.цy������Y�S�^[�b��=T�GD��#�u(�� <�糋(��@gfJ��x@V�XDe�
}�'Q5�9X�$��x���y1�ؾ|瑵P}�YP�V��R9��6e\�vCH�m7Τ
��s{��s����5���' p�0)t�9dǰ�rCp�Y����F8��*"�PJv�a�.��$��Xp&��bY��jY����'lt�7�x��jt��	�à�<A��k�8-�;�b�A�"�Lsjؽ�KX��� 6���=!�s-HE9�$f�:�7���8ō?0o��ۀRf���8���:��0�/��2l��栖�4�(�[�E�յ���8a��Q��M���n����W�N�L��V�c���2.�?ޝə�B_�&��E&ɍ�#}�C��r�m2�p���B*"���D���s:�S|s��O53�9���@���/'��U;h����J��|+�y�{�H���?��1_ӽ�K��F�x"Q�nG�o� 2�7�\��D�![k��V��J�¹CCT� ����0��h�����m¯9���k�|o�O���2��Z�3aV) ��pN6�WUԈe�Q�^ϳ,�F�Q96�bu-G��s��i�eZB����Ce�b������f�5�G�.���E-���qU�3�m�{�dFAX$9�tTylO*k�Ah�t����n�x�
���#���-�аy,����׎R���*�5s�z�a��a�=%��mf�vLe�AJS�r�Ʌ�LMs�z��gx�@�0\��aVwn{rC��ǰ2��.�G�MHD��U���-IKZ%�֎��[�et\k�f?����񵲩(�q�ht�����/�ՉW��Q`��g� 0�3�w�ÌF�Oh�!�&���_�ac����CC��\�>:��!�p��@�p�i��;=t�Mt�"�gyI憧�?+b��۩� ���5`h��B Np��ԗ�l���Ι�3�B/�9���>��[i0�!\�����kEǩXi�4}�����QQ�AEx��ߧ�Q�%7��Wb`��l�w�h�}xk�]�&����kS����I� !�@cQ @(#n~��n[Y�D�m�
�J�����p�t]�Uۧ�:��T{tA�&�ߊJ��8��a9�
p��ϩ�Y�.,�_,��+�7����?����~�Z�3.��`�0�:O(M���=ͳ��F����Y��P}���P)��퓝��úw�o�U{]jux '�C�G�?��A(�B9�T�Maoz|�X�8�S��AG��~3�=���~����`���Ќշm�*���=ds$0r����De�@T�!?Y3P�R�X���f��_�����:�B�z����ڐ#W�XZ��>(��}�WP�%bm�95:�S���M�c*��͕x�`q�wFX��|�L�C�V:���s�R7�Xr�4%;(U0�3Ѧ�u�G$��U�	>"�)�`�+k��ʟT�3!{ѽ��1�Օ�F)��@86��bZT�L�aQ^m1��<��:�,��+<�����?Uxo�6���<
�u$�`8<J�N�	&�2�Vs����W�ζ������ţ�]�Ŕ#��g�v�d�lM�N2w:��T��rS͕'����1FͶ6�R���46/>��k_��l�
��."!˓��$��/��iJ�u: �����gW�"�cS�Ҷ�ޫ��N�w�{u�+҇��H<���F��&�пC�[n����wO6p�m��/GG;�dK�h������~��I/f���)�G�5��\�ˏ)�����e���ʝ+��/$IR����fʃ��<G�������j��U�P<���AeG�D����<>�N|Wq^��V�@Z�"L�R
8��\c��g���or׭/�ڸM�x������gU��j��Tl�Щ�]G�.3�;�f�ž/F�����0�Cݎ�r_oyT��@��\aW@��6��N��q:��o�y� &q6;��}�j������H�����(S�0Y��;j|�p�u@]9�����
�Y9�խ�aA�gP_ۦ�]��T�X�L�Lr(���L���jI�0EO)���"i*����8R���J�B�}b�cв("�9V��Y��ө�f�}�f�4��NѱI& $�Z^��ų��m��nx�+�_�����H�'���m����m��M��C���#� *�6}Q��+Vv&Q�X�$]�D��m��f�|�*�^7s/O$�aO�^�P?r�W���V�+Gż&�I*���#M�M�X&	U�8�� 
!�����5�� ��;m�e�ܟ�������Ȃ��h���,��s��=FM4����f&�:i�}A��I�ga��>j��P%|��Yi�&tml.R4%�R���h��A�I��Ն}��^� \��a��p���X�VV�ٍ�!�����hC�\�"��v2�]sa���\[����gs�]�E�?���H��/>Tlӄ\��Q��1d�o|���9�<�eL����;�����=���Е���m?�V�8|D�Wp޳J�z��k�5��I�;^!��ZE��#��� �l��G	9iZ���[�g�j�V��=��ԯB^���}�gx�>���<��._>�§�#�Re�����]�0gS����q���<E�Wˋv-�y�D���l�����x��ids:�6��b�z�a��l��J�Z����!i�/����Yk��.�Nz��4���������kX��e/�!���:z�ު�@
ž}ς���ے�9�U_CO�vq��|��G��}����I�N҈�֌���	��w9:�����ID�Kh���t��������gp��k�"�fy�Ϊ;ݓ��9�����lɩ�<x_9�/&HTY����L5٨/h��͹�A�1o�,���T-m�׉�!���*rf�4n�x�	������M�p�e��af2\�$�ky|����ǂ��Df�o.�����/I�7{�
[;�#c��;������pC�xq:��o�U3�,��k!����Eǅ�3d��aK�
{��m�crE�1���g�����GCH�������d>�@�}�QZ&�G���#�t�Nx��L��%К��O�մ�7������0è��Q��^?�6�A���Ok�;�G�kؕl8e���b�Ǆ��xw �/��C�Ъ�R�0�Ě\袙&�F�����Ҡ�W�R��xG��7�!1��	�$*�n��^���jf���cr]�
5�a�z�*��V�t���n�=�Ï}/��nhtZe��e+�u�pߧ��L���KL��5 �?�^��v�ɥ��	��lg�ʙI2�t8�a�3�����tMb�yG�|y%o�v�p_r�P&�{��D��ۢ9P��Ӊ��o��.�2���C2X���T��ʦr��q��e��M54��%�v��mn�E�d�����z�R#+��'�'\�#C���A�-�4��F�'�P���)Q[��f��rxZk,˚�p-�#l�k�UU��,�_��B����4�JSG@"��o�_7f9ϊ�Qnk��)�	 J��'���{�W:\��v�2Xb;�f~y1z�����M�[W�G�wuh�)/e���Y�����~��֎*���(���:hB�
��j�b�eV֒u(vaǽP�����ݟB�D {��8�y����s���z`�I���.�@�|�rG�D,j;�j��!Ջ�<w��(?l�Q]aB�BuR��4�hmEUd�r��p<���!��d�n���I	��l��0�*"�%�b�΄qW>���+Q�sW�Z��{�H{xA�V�����	�͔�WT�sp�/OΓݭD�z��u�h�Ww]� �<� �I�AL�k��A,�r��i�8�����1�:X�Y��G2�x�.S ���-�!Y�U�{���$#��#R͚T��f��lw�AZ�F���Lo�k�U���'r�L:�yW���I�������F�h��f���l-*Ў���xrЫX���j)4��ڣ;�����J��������&��;�{�b�E�HY��;���XJ�+��O���y6�g�P��Ը\`�lou��6,�t�2k������eO/�(�Ҳ�v!*����p�u4b:�< "D�D�@l�uT�,m�4t<��G�an���휛!��Rh��}A5e�V�D(��h�a�M�m,Mj1��C�����)�{��*�
�!�{Z˽K�۬���:���סEe� @�"�(6?d*-�Y
���j��c2i��/ U̢3Tv�~�ɣi���Q�^�l�!�ruFbnE��ȈE��f{D������0�*��7ˮS��o�f%s@)ȵ�zx�&��_�����S(�����ۛ9c�$-���I��.x�J �C�e_�ɛ�WrJ#ͬ��kksUOg�8z'����=��Si/�8A�� t��Y�܎���kzn<I��s�y��Lt�1��r�I�,#��<5Z�]>$��t�f�.u�QTt)S]-j�:1[�]�c����;���]c�D٬�"��-��өb�e��x�gg/�&��XcǇ��X'���i��(��	��J`_�~�P�d��Zč4���y^Ee����}Ἒ&��y�6�N���Hz��f,�1&0%F�����ǽ;�G�P�#�4cΥi�����iS�:�7���J_6p��i����F��8�}q�4. ���E��UUն8GH#�xũ{�c҄���^�l����Wг;�eID������|�P�Ԁ;3�^�R�|!3�ԣ_/��a�.�{���W8�7�\����;U	c���K�%� ���k�-��A(�ۃ*��B��}%��e!+��ӽ��jP#��a�zb�H�v<9.�b����+�Xo\���L�>P�d��Z�i�����vO��J{����̐�N(��[�����5�dʓ�H�p-�����[�X@̸]�Y�ҋ�W���o�U�X&ф���I'K[�Я�߯&Qj��VNJ�2zb�TKA�G���.|����im'�!�&��T�ϡw�4�儮�!!�A��)��W������T�l؊������ܵ��^l�����M�Σ|��k���U=�Y�uw'0��$Bǿ����_��*]^���>��*�C���]cG�^J���a�̂FUE�ˮ�:Rת�����g� ��V���j#^��"_9O�}��^aw*-�!��[!f�5�ۥ�T�U5Fy|�8&�o�g�n�L�B�����V6T����!�uȟ7��6 ��%_ʩ_�)��#��F�j�kx�
-������&N1r��a� {�N�u5+o�n����0!�Q���މ2!�7�]�D�H��(�TE��X�]^GM�_L�&��r c�j���W�ɫ�����=�6	V�Z���ΐnl����4[�cNr�Qђ��%�m����]�ѬXQ��i����N��x+�Ve���q�h#��Q';з�U57�����/��0�Z,l&�g��0��g�uֿB{����X��<����w'��$�����#�{�2wZ+J���f�24�x��ڍ��',M1��_��<9�}�1ĩ*�
�;���}C���̦����=�'"�׆`I�N@dn�L��rY$$Ć.���q'�K:�j/8抑t�Ǿ�d6i��y4c�i-݆6�4������X�0�_��0���1C�q��]��^�8Y�	K�п����9�f��ǵ�T���=��?u�����-.JH�v>0�ʵ�X�<���8��(>Ts_ŉ�b�56AŨ'T����i���!q��E��$��6��87���cO����tt�I�Mcv�w?^�c�20A�U��Q|4�X|�
6Qvf^"?Z ��@�U.��9�슥$�(	y�X�t�R�}�~�x4��~�^+�<���Kx#����
B�3����P�EN?�%v4|�����jqB+cB9_��jVZ��S���T�d&��.�$�Q.};!�#��4���{���6�<����#^ R�_5�mOE�{������<Y��%�[!eQ$��$���]adC����<i��p��u�i �ih��JZ�]S���d_���@�����	#k0��$�`e����\�VhfZ�f�dh���N�Ne�m�S���XU��������Y�p"��z�9����́|w�k����}�&I�s@��� ��d�:=�_�o�i�`��iz.���*�NA@*�&!��Ҽ�1��*I�[�\V�b����:"w�m�~	���`�h�O��C��j�o����Zu�Dug�:4�g*P?��g�*JM�u���HR�t�rfm{��qֈ�5��ڛ����qN׭�J:H�^��B�Ԩ��w|��?6�[,� ��X\z(1;-���Ϫ
�0 �ׁ�\ĝ��j> �	Ep�/~ܼ����ROU�.a� ͂��m�b�
��愖�O��(��i<<;m�[�ޮs��_�-c}bi�Jl�O�زdH�C�d��?W��/��D	���ͮ�& $��T4cmRN��"�F���loU��V��RQ.USS5 
�,t	��KN�j.���q��Gst�V#W�+�E���=���۞*Yν���8�&�L'�����(5��={⽎
[��ɟ ��G��Ϛ&����ͲG�!�Ugj�Ƒ��������R�Rܾ8�2Fb�K��o��Nv9�2�	�k?,��c�
��vn'��HQA��L��{ܑ�p�B"���^�!}�}٢�P<�����/�i�y����򨃖5:�0�^ӭ����!�9�I}�R̮��SRی!|4�����։v�Ci���%,fy��U���<�f�S�0 R��7"k���e�]���|ˢډ�[���=������8����mI$2��(B\b����z����HW�1�-De$�V�0����s��<�R����W[��v�)u5���N�o<������3f���ޅS���@'��+�h�ړ�E�E2���D��k_�ο律x�H��e�� i�si��Tـ"������(���C�*Ǒy�Q!NQB�x�ro��C�i��Zc��J(�!o�n�-MT	���EI�`��xns�J��xF��>7l�������@�g�Yjhݭ|���x��4S*�	�M+��8q�JdM�$�gT��.���X��)��T�O>��qn��ցzWЌNw��{�\w�7n��:[|drH��i.��;�Q��s�/�3�ʙ6얍<����/J���,3���^ �OD�ZV]Ńe�M�4��º� ź$M���΀f�z�@�J�F�o��9��{2vsn$�S����yn$8g���^3�y�yֲXH�`��4�2�2$%x�f ���C�r�򬍅�Y�N���%�ĕ�?�>]r�d�]ucǻ6�T^�Y�9�q��D����D���:�p10P���сz��\�������6RV6���q ����ېe<���a����U/0}#0�kDU��Z��[ī����F	a���5�g�G�p{�O��T��[ߑ��<L��ܛ,��б�ˀ<���� ��	����6�+��
1�\m�N�����ZxV+A$������y�<M�{�f%t�&qlF�*P3��GT���\�p�g�Y�NQ�tN��d+�Fd�Hk�������C�k�8�����p�u��ՠ�����[�d�������١��#�0��2�yVb�ȋ}���Q��ў�^LGY$�������ɽ�������Yb�vU������bI��G�(aٷ���y8�Q�J��߇5Z���7~}�$��. �̈́n��C0s���	�G���G����`5;��!aU
TV&���F|�AX�k4RHdQ�NP����-�����If�j{+��{�2��
+2����/�i]N�I�5���)���������`(R�dޘH�Ԕ��^�P��r]���Ss� ��������N]��EŞu�aP k�ت6H�����,������ʦ��^K�A�ȣ�lf�K�r�c����v"�ɳ�o�A���8�o#��s��˰�-�Lͽ����a+y����-K����h�3�a���ȣ�<[~v���m#_!
ȕ9�G��	.�S�0xd�pl5�@T��1rA-y����[��Y�[��=w!� �ÜI�T1/L�&�i�<�
_��&$(��_�����%dn�Pd��P(o��>L�=~���{�줙.%�R��"����O�i�A��,Ԝ0��tW���	D��ծX9�Ƙ'�|�⩱�+���o�����`�Xifn���Q��WGlC��7ڦ�@���!��)�N��y<��Rw#:��R�)e(-ꔉ�γ�Ug^x�@UzX!���k2z�N�r�M��"���2cP�a��q��*�����6����E�|m��&2�D��W hӼA�=^�n����S�]��r�[T�a=�������|��U�R����x6���u�W���%�.CI4�|�?lP���Ɛ��N�_��ة��;��5��d5�F@-$��B��) j��R�&Yɭ�^����R�(9�;�N���O$"wB5ǫ��۰7(h����n�X�8���G��WQ��7��o���oo���-�K�5���ib"�$;��v�?��@ڵ��o�-��	;��z_��9pZ3�^���M���S�2W�w�����)c���-*p�h<�$��jQd�ha�W�2��W:$��͵�����}�aW?�f����j�[%���WSȻK���ozu���ժ����R�5�>�yµ�*w�vY�O�����✝�&���:EXQ�7X�Pj`�h�8ǳT���2�2�z�X���D*
����_=�E):��(;ַ_/6/ �ӆҺ0E8����sW!f�&M�2�E����&|+3�Մ�2�b*mZLk_S�=�&�)����|��H���*d�-BO���>����ET�_�o�����j�GC���Dc���Y���l8j�dokX(q �����B`��޷$��a^��.��I���R�u_�DNt�経�~��C3^�� �d��X�h�n`UG��X��~4�-g8�α�a괇
�nb�J�.۳��a4���IS���I����(�hG�̝����e�(�7TJ̩�tH�vZ�BV��ݡ�Ё��[7�k�H�5F�%��ڼZm.a�{���8&��j���o$'!G�ɱvnw�q8M˧N�ğ�/ ���j�L�0��>������T����c/��1l�vd[�m�V5ǷXث�2|�rJx2cH8�������~۶��1���){PU�v�A���p�Ҏ���`;�>�0N�,�����C� 3O�ܔ'F�ʴ �8|0I�8�3	�T�Թ闽m�"�H8�?~�]^�b�K�	y�&q@�
S`*�^u��^�}������k�=�dﲕ�x���&�C/;����?�1r`��@�x�h�R��1��R�p�������(������"Y�e��'{a�K-|������30���#X\)�K��)ʺ�W��;S�'�6=R���;AG�����3�������iQ����إ%��~b�{�$�k��(K�UƉK��}����aR��ӏ�5ؖ��,���j\`.�(�m�R	FEz��C^IVμ�ȓ�<S?��L�c��1��y��4�
Z�ȃM�i~S0�ي�;��d�/�[����=���*�b �n�k>'�c���Voq_��7+u`��@u�����g:���<Lb���?z��I��X����x�i�X֎��G����.����&��BNL��0���K�D��3/�f����`_�{5���:%c�'Ak����-�!�n��0�np/%�5����ڏ]Z߻�m�}�Ӭ(Mw�x��b�x�q����H���U�LV�K2���G3�t���g��GLB�vM ���Ĺ_'to�4��=r�hX�qC�!��Á�kк�^F*��?3������|ܫ!}E�H�G�e��'�E�~�:R����0
2����ur���@�����z��A&��Ue�Q�
�C�$p�q>_W�����AB�g�(3��ڌ��<�AS�Ɖ�6-����ROf] Iߞ�+}v<6�j��/�zB����=˛�����أD0��G���z8�(ְ�
DڡJ��s�����XZ����E=W�K���47��]3 Q�]s�SsK��֟+w��:@��i�d�?��JO�o����p�h��v�4�g`�ԝ��8�h�����(�H0�9� �m�U�
�k��4���7��-��S�f�R;��wF�a>�=�6{�p�:Ҩ�3w���(䄗�)��@jeX�P��NUq;�es�U���r��W��T$p\�Ӛ*w�WW��Κ�q�.�#�"�y��"tu`��t�R��?NZI=�W�.D����	�J����i�4�p��!O��>a�&��e��$�znN�	
�b�3�w˭�I!;���tOr�݉!��mDc]&�c��s�