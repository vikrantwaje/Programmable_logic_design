��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2c=�Q�	�l=����t@�����C�g
2��� � o~��R��Բ�.�)"L�A�L�TJ<�R�qԬ*��\ia�d;1~�
+i�Ax�����k�O!�4I|R��Në��{��������3�x���;B�E)� ��8�j�}D���ݺz�ї��q�ØM��a��%��J<�f��i�:?0Q/^����lw�$P���GƋ�u�����B+������8 �h�|d]H�P�Q���^S@��wڛ���v�Ѝ��P+e�z>�څj��������]�a#�1K�3�g�87��-A���/̄x�	>����.�X��JWWԚ�fج��LOx`�ϫBkq�_��L�ϫ��<*έ0�d���E�Ξ�|b&��K��fS�L����
۱r|;h�2�4X���r��Mw�KD�R+w�ݱB`(��_��i�;Ӎ���L���t&���>�ׂ�{��G ��wY�(_�����[��
h�����,)���N��·S����y��U6j�P���'�����d<���h4�. d���#��]Y�m,�B\���Ҹ�qǺ㰺��%�:�����^<B�	��<��]�
�)�r Wd�>����n�"�����+�2&'�%�_ai�	���t�yԡ@_�k!�imS9"�}�N�)����R��Ԁ�����9�c��n�-4����o>\]d�+檊�-N"�I��4*�!����#(tJvM7�&rm�I6H!vN��AA��@��T��f�m�&�=�V�)��j~9"wҜK+�����#xǟlvƛ�p��^P�0�Ʃa����I��CVS�h���Vt�vؖo\!�.�B���a��.xiݷb7��I� �9����i��-Ů�]7�v8�Fq{�
� 4��(v)��.�ё��׀v�����ьR�),e��?���ܓb�56���(� Ֆ�A�X\���A��PȀ�Il� ���|�_�?c*#5}�,oD)lS5���Cg���{E�F�}��B��Z7�:#��&��y
:��/M��q%�?I��O'�d��R���{��-� ��e�cGE��!'bSC�$�ܪ�ݤ�*@�F�A��W
���KV&�� 4�V!}�bD�"���S�l>�s�"���%:C1K5�����6<��-|ϬC��^�t��:�m��*?D���l	�c����8@j&�T�
������t*��S��` vz.sY��r�v'("�-�/?�4���)&����DhyV��d<��MF���݉'�/��s��tX����S:$~]&ڮ�P¢\Y��V},(p�gO��q���G@y��0�B
�f�}�W���5v�u�Fݢ�"���ei�<y�&:]�P^�����f|�
�������{%ۈ�;���|y��
�KN��Kh�}iVt�y����8�0P��Z$ԭ2��w��ʀ� |���O�ek���?ܓ0�Mw���d^Ot@{mg�k���ꙿ��>#4gޟ\�+
p>�8�%E��7j.B��?3��ӌ���z"/UM�8r�,:�7��RN�N�8�����<dH;��lWc����" 9�g�@il�����|ت|��N(Q�Eh�{��J�}�>6\�N	��^	��突�ݤK�O���6:K_��/�R㪎��9��<��;�|`ض�.�ѯ��ǟT���ҽ�ms�E�����>�����2�ka�$�8��o�
��uP�b(�� I��!4�cc�>��:��q� �
W
!`�5>Y�#�G;�+|��Mi��cƌ^�C���nV,_�@��yi^J��+<?]����h�Jr4Nv,TvmǕD� Z.�1�LJ���.G�)7��}h������e���(YB� �5��6kã�,ur���j�Ʈ	�������x��M:-�:ƿ���+�Y�$b�zOO7�k�g���k�t�l��Iv��H�l��K���3�5�T��/-n6�W|��П��>�8L7dVQ|�:�yw0p-�1h�j,���|��SWʨ��}
�ú��XWv2��~����㒟�b����t�b,�b8����H[V��7ي�� yu�x�����KD��`x ��v�>���k��Q6�O�X5�X��]�CL������>��ĩ�b�Q�T�~	�*s���p5�-�����'p��$�:����~nn�
6J�ږ��X[��ɉH�d@�B͉6����`<I/«AǘRyP3��0:�"��v<:r<�*�j�4��U��۽ K��l�^�d�`H2L�[��۪j��b[xź}	a>V�^D6�&�D|�&�0U�Lp2�ݻGv�[�����z�7#�
�Q���B������1H�;�s`�o!�m�F򋲅?*�AcHc�������%�Gd�JV�F�R~�q9�=�J�C
���x�9�X�������S/ ���i�8�^�q�X�辊����i�1M)��;��]�(��g0��^rn鷍)Z�_�~,�d��j�5Les�=P5/�-e�u�m��L>�X@�H����I���6��.��E;��������|;l0=I<��ˠO�k��X� ����<�/@��a��9��CG����?4^3����ܒ`+P졘n��C��d'
�������,T�]�,�*KG+����k�H�,��=}��i4uw�z�>��S���lU����"��j�Ŕjf�3d'n�P	N���<���^iQ��D~ 6��5K,���jX���� ��X�ka��Z���(ť��:]v$�y^�
�V�>��	�MV��)��;�pg��E_V��.�z�ۧ�9�4��V�%��>Oݤ(C:�]=[2GY���h�F1�Z�U��4�HL7�
jS�+r³m_�"ԍ� 
��s�핧����U������?TWх�"F�y�[�&��p�~yS���%H����KȄ^�zD�!hLOpo�l����ps�g�/�=U��s]�p�M�i�om�V|t����Gh#�+�^3�M	z�gk�ŗ��tl=�E	y}[@���-�[㨲�0��F�^F�o�蜰yh�A�<���u
1O���WGq������	MҢkU0��	
�1�[�j���P��<Fi���P)C������[�k;ҬLkW�_������=}�׶.{�^�(���5v��u�8ռH�^��e��Q�5񞄏Ƹ��m:�����b9��5��n,�D��B����ޖ���%�+�(���N(x�8���<W��d����~�����a�'�y
�^x\zO��"4�f�RY{#4La�����ku��L��x�oN�,7�;��`e9:Y��<����M��G<�K]ʍ�۵��Xtv(�q�&>tR�s.��W�a&f��|�i�
�_�h�����ܵ��-͔ ͨ�䓬�G����Ba$����x7(��!�8bKe&dx�����m�Z�>�{�R���t�Oţ_��[����'�[��t��/8_�Au)�W`����cb-2���6h¨���۠kZ�w��/��Z ��:�r��~�O^�����hb��� \!�/h�~~� ��C>�T�}�F�EE���$j	�8p}�b����}G�l���B��q��'���3�x�����:�H�6�����a4mR���%��q%��M<�=/�3X3��A�>�.l ��p
����h�p�QZ<Y���_hR��g6WO������*��B/˪����`naɦ[w��m��$��6[iT)�����h ߽�Lٴ���M�@ˣ /�n�yy����Pi�ir T]L �~�M�d�Y�����5!�;�M����;���0��eq~Bh
�r��U5��=�L�5�"3㹃M����|͍��M�D�e�i0��l�1��G�,dcS�>����+��r���m��( ���aEڌ�,�+4����$�!�=�B�ό�}o����˄�����	<S�Z��41Lڭ�K��S��1쓢����$�z`�\�EZS�CM�����	�������?r�QM��8�P6v	�7;��3�G�^��T���/!zB�#��gca�c���n1�������P&�SRm1� ���b�[��dC�i^Ɂ�,X-��i*��=t�/-l5��hug| ]�l1�8�x��Vz�*&6�0�d����ф0�J�]_J\�`��y����d�vOڠ�$2ք�=����і�Bl�����-C]���k����08٨��ў^X�xbH�F,ʕ��F��)��
d�y_�wXϙ��DҚ�J�b-���'�Z5�[T��W��/c�h���U`Qюg�uɹKw~ z�����u��i��©���pH+S�K�Xo>�	�uX���#=���E&C�2�5 )ќ{Wtn;��V���\�nQ�y[R��� ��;mĦ�׵��]�R�O71��|M/{�� RW�1YI�����y�c��r���CYt&����#[�^a�{�?���3�i���=��̳v�;3Q���z���+A<��:(n���(�n",r��/s㾓*Pu����vg\����I�k�$���� ���g�� 123����VO3^��tf�wn�h%���=�i�{<����׎O�g���x�3ݕ+wM�\���v�q0��E
�����t��h4��-��3&4��6���Y��^h>؋[�f 7�r8T��y9`t�|����bht8��s�y�ۧ��̣W����G�Vw�j�:b�������w?�8�cϥRXӏ�ې����6�������;���,�m�	�@�APċ:V��� ��^]����,�K�2��5j�-��	gAf`P6G*6Κp���bK��J�ΐ4�7mY��?�F�ݎ߱�V �tF|Ƣk0������8���Пs�����̵|�,�%��m5���%��G�b֩"�O��6�����/1a�1>GLO�>sߧL�*z�5�����2����x�m[V��OY�ŒYJ��69B�X"وl����X@̡x���p8��E�Uz:��3vXjZ�6T�2����;��ݻ5�H߼0��5G D��*� ���ٸv�����q�s�3i�G)��!�w���x�JR�<`V��h���S[���#�9/����=������"n$C��E~����,��s
 n[,��b'�v�,۴%˷���������>8��;c�JڑoB�K��^A�5�Pm>y��Jn]U���GX�OQ9a�%$�d�hf�ܣ��E��CvQL����&�V�sKB��U�r(?#��u���Ǡ���k����M�=�7�k���w%n����O����U�c�#���x#f{b�)%d�f����3��G$��Hr78�/kI���e���܋��
�����t��$M�����O��k�3~8��[�5:D�Q�?WW�I�gU��5����׃�2����=]&+���^ Kh�xbP@����?)���kLGpM�:�Q(�܅&�#{���nΜ_\�>7�$ϙa�(Q���7�*O%w��D�8�GX��{��[$���,�Â� m�3E���dS�/[Bp-�����_W>�*��}0�!g���«�mK4����L,co����u�aQ���t�����q�I����U���ό���D�_ߜ�A���K�3�C�s�mE�
�:�t�ZPbF�ـ��� )��+��@��ؙ3����j�M�ؗ����**�g��R�C�9�d>i�]`zlY.F_t��nD�9W|�|m�^;���x����of����a�~מo Cm1Wℨ�-K�g:��yJd�'}�Vժv\�?������ο��]G��<�~�ZW�I�)���vVr�@�q?��h���;�����������zdx`����>M���$��WX6O7�CD�-�ѩQ�J\���@�׵ή>�����_:��,�#m���z��ӯ�%��q�S9�-���X��s����S��xD �zZ��H�������\F����
��WG��qVy���L�ytK�֮ك;�_��x�ʎ��o/mX������S���o�<�Zq�,?H�gL�rxM�AZ�]%\�J6�e:�j��u	x&�qT�m�C�Ȃ���a��mw�$�H~r�Q`�R:x6#�E��?������ %�䰗��DD�қ���Iǈ����� }�E)�ɓ��j���1�z��{�M��1���f",�u	������(�Ɔ�
j�E�����:�$������nC ��=5��UD`5ITU��$�o�J ��ӆ���l���)��ٗ�d�ʷ7��5���4!���H��=A
'���,��Is房����S�vBbj�<� hd��������~qUO��Af�;�Z�'X����	I�)G"	�H���t���]8Y�����0��?��Da����RE/�&x��֞�6�eH�p>�K�-Rx��'s��R;�~$���ʠ�����'
��_*�6�0��yP�b��i�Z�]�Jx��W3�x���z���m��(�%2~��˧��B��L��lv��>z3Cz���OV^U�8� ��^�Z�����js�V��2ۄ?%R !���|Hn����� �����^o=ok��{*;��9W'ئ�Q`^W��-����3�]�����S*бё�"�u���7�U����FK�ey��4�jhO�q�V�<���/ ���ָD�MS}�]���D�6~����|4Ujp��Pk��M� ���HF$Ê��W[�%c��>-���n�*8��;&���B}|~)�t�!F3b5�/��~�V��Ǚ\]�_��gށ䫝񊡰Rl���|w`_�6@�R�"���N��T�E��ժTqs�:_[�}�v�An'po�G��*��Ⱥ�B旯J{��@�qМ�x�g�Y鱽�$n1XW�u�%��9ޑB�������p&�����h	�c��6i}"�8w�쓁�V�]!.�H�#)���̲�vF��.;���Ɲ��ezٷeI���H;Hì��:Y/��ᮡ���qf@�:Oꭑm^���:ZR��Ț{�o�U�.�C�ː#b��8��Jg���yh�4���u�R>-��<�<�D+��>��Z��]+x�{z���u7�׋N�d��_��r;��dJ�G�����!P���;�.qd5�>&˔
�)�����%����-$ߢg��!���zz(��7E��rhJ7����K��K�=��Y�$SCB�rK-���L�9q/�ҙ� ��hO��"~���M�Rm�C��Ӓ4¼f��~�����q�|�dM�޳��j:�P��(;��\��c���{:�G��?i\]KC�%��+�LN��t�fib����f��pSЍ!�xDW�Zt���x@)����	m-f��~a��w�{V���&�dJ3�j�l4�vb�g�u˝�q��b���W�ag�T10�0>�{�'�y)�ըZ���U��y������A����R�$���˪�Yį�\�c|�Ry�_�]Sh��F��B��
9(�W�A� c~�?{
�LtU��/�5�~�kQ&/},_ኁppq�2�
b?l�pF�6�����#�Wp��Q�$��۪Mj�65>͋��5�Owt7K9��=Z��r�~��&��Q����-���B�"q	S;/�X��;�+���a���Z)���N�o.�W��9��H��;�Z�`J�rZ&HD�ҹ ����8B� ���Y�h����sCg���b�v'�|x�"��l�/a>�S*4;���H�HX��=W��V_~�ƤB��W1E�B�mԟY����?㵡ƽ*��ΧO¸�_�aR� ������f-y�r��In!�0�4��7��$75��ӵϴX��np"Yͼ@o	�W��P׭�D̏�'��@d��@�ƶ2�~�-�4˕��-_��l�V�j�<���bt�jK�*A4H�MyJY�������f��qL���W�� �1 f�����Y�N���'B�C�p{2S�-�s��TW8�&0���������@[���Gn�k�u�PJc���B'BJ\�[!r��Z/IGi���	�F���"Cn�[R���1%߰�ϧ�.�UE�]���}&4E�
���-�-�Yi�Հ(n��ьi=l+ц=�5՞�6��P2��s�ߖ���&��[�XxB�g^1���iƀg3*�t3�k��Y������/�%�B�BD`EU�]��n`5(�����8A���'V��X��0�WGw�����;	֏��$ 9��F�Ls�|U�汏��� hJ}vd�K��i�6�Dh7k��8�|�&]eXQ}��WK��ǡ��R�t��w�O�)�G7V���� ��=��Aɣ6�ۈֻNem����$�����|�h䙀ַ���\@U�$.ef��kOR!�q-U����Y�!�����~X�@��+�u�˱�^;|���W�z�,dy�H�AZ���%Hv����u�/Yk'�"M��6�#�t��6��ͅ"�*I�AX�^�OH4"��[S]H����tB�[�k�尴j�2�$��ײ���2I�A3�W�u��%�m�V-״\�$A��A_@cr,t_\�fHU�s��X�
h�������!"d�c��z�]�Hz��U3��m0Q"ڙ�5bk��( bu�������vCd�4�&�U>
w�h�F����-�.	}P��=N��(���vu�0,��aua�4R(�=[U�M�M���V��ܯ�&�k���Aj��!��BV�^/>�6|�[��b��!N5B(ů+���y����ɠ>y/�b��g* �<���N�� ��6�x�b�������ذE�X*}�i�2�9' �Z�bğ�/ձ�y	u`%��@p�-��w ��ڝM�"�MV��������(�
�0	Όz����xq��4�ޔ�>��/��u_9MyN�fi�6��-�|%r1č�|�a�vMYn�w�l��Smk�4z-�_�L���ِFs�߳3? �� ���0�
���K�nc�P���p��_�Ta_�V�@�@�+AO݉�`U~CyT��Uf?�3�!��m��ƢCJ���A���p��s�8��+"��#ee�v �N�� 
������`1��5�L���1k�Y�SZÐ͚.�^Q͜i��2��[����~��-�^���'� �r���d^�#ו$�!�z9�,`(�^@�J����GzaE�c��Wjv_�05�*0�!=����W�R|��ςf��	`���0��<��΢�7+q��ZP��s��\�V��+�s��J�1�2�6{j����W�8ֈ0���*X�)*�k
���qŔ�h�ۀM�"N:MiHJ����~�w�����c����4iĻ@����c'#�YI�r;Q��Gk��~*V�����*x���'����,N�D����8ǋ��∹�� ��@�߽�<rX	��$J����H��>�̈�)���{p"��0�R��W����1��!"њ)`�NY霴�7�F�fXD�(@��.��	~K��T�@B��'rӟғ�}^ZjJ�6b �w�5�.A�l���2�Ub��#�.��,9S�ĝ��*CjOo����19���n�M=����sRޖ�S�hF�B7*&�Zd�n-����Oqia0�:
�tu�D�@
Os�ƥ&�k	gS�o�z�n.�t!c��,��D5���7#i�����:���ϼ|&P7 Ƃڳ����}-N�C���0����Y|�˱[�8�JǠ����B���� �J��<\�g�z����We���f{�$z�?�[�I��?R���P�f�0�<���d!No�
�&|X�z���4W�ʪWF/#i�^����mx����C����$�[����l����	4�J3
h-p3R$�J�.���̸0@�1����m���8����>�q�������vM)��ZjL��ϸ.}]�c9�� �
dr�TO�EW�H��UJH�cUA�5��(,��]{�v��)���%�6D$��r�덄%�aD��Eh(JW�fݮ��������o��ә�@�>�Ƌ��������/9�����>������B����9i�Y6 h�ԇDC�o���b��*[�c:چ����c�tdZ�i7Vv��5�3�8���m,�(�EY���+�:E�Z�x��$����؃._3��J�*�g��4� �/�8������`2���N��V6$fO��@���7ظ`�UE�-����0Ua�	z��5��B1��2���ǯ9�5�V]cH�.@����3�'�r���-L�\.�����ك?��Eo��X�6v��cV0j5������a��5���}�ǽ0�2z	���$��x5���ׂ�{�zh*5�t�rY-����g�����[��?�/:���$�3
Yخ�o�<��Z�o�p=��_4Q=�-�����%�(ʍ�ؓ{�	���0�W�r�}t��e#��ؙ��k
�Gĥ�f �U�CC��΁��n�cG�*�W~Y�����O���2Dv��'Q�����D,�i��<K⑼��q���`��oV���'�ñ�&��c��]h�m)�A0�
UB�^�rg��nL�\-\�8�^�m�L�T�O�RC͡�Y�Q萋U��(��a�.��X��m����z�����/c���6'�C��[�=T���i��9�m����_�T̲�6���2���1��U���j��Tm�Si��Ҵ��o�;�����Y�3b|��;�G�M91���}��N�F�ܿ�qRBz(*�^G���ouj)dM�T����x(���� O�[^9�����V�}�%����/e�\6�����r�~@:��<B�
�t� 2-'GBUÖ�S;󄦂-81���+�����>��t!N^�5/b�y����[��R��Wu�����i+��y��o|��V3о��DΒU�
�+n����u;:����.�%D7��	[�i��+����;~��{&v�ő�� 2��CY�\(�]zK�]����Cqؑ!hb
�{c$�ي�`�Ӽ���<��T�j��#ЬF�aQ~�����\��3�Z��Ƹe+1Ѐ�`č<&���s��5�@���b�vM��k�"�!` �lW(z�Ɲ�����x�%]z�Zصl�C��i���؃�pK3��OI�'����||�K^Ֆ��j�+�C�BP������~dG*���M���#�|Z�Qym�/��'�����_�U���5�t�'Ѿ;�؏-���x��7�|�3v{�s7