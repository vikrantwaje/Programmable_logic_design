��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d้�^��r-�>��s �8������h�Tw#���#/�x%������N+*z�ăZ�4;L�
�:��"p�Xa��(�����g�))����<)��	K�>|�	����� ��"�ߵʄ�7t�>sђq���Y��Z7g��^��M*ϐ�G�飋��69!�xb	 ���5��G��r>��T�CF>�br�Dtݷ�ǰCD�=����7����Bq�%�(_q�mJYT��U�4R�/��~�/�?��Z~���1"l��X�o��vb��/"������Q</m	����W��
�~�d���O*{�3�HS7�0�$��oܯ�@�fөLh��֊���X�ȃ*�בGWy�%a�]�G�^2vV ����O������OE@��4��W֠��~>0��g�3t"���q��#�6�����jW���ۗU����Q���H�9ӯ���Kw.����oO9K�Y>�f���˱���5�'��lb���;Π2���ۯ��D�_>/ƽ�>Ak��P�[�Зc��y�+�~˒x"(��;�F_�"�KHR��C�ub`(�Uᾎ�;7x�-sS�"����e�p��s������q��
$ڀ�Չ�ŵ!�;����%@ә�jo��#��(��X���/�˂'3�ܛ���]�q�/225���1w�:�[k���㕊����%ń�t��fH�v���N*|)�°� ��!v�i"H�a��͖�����~�|'/n��: �EK#�PZ�a��?�S�l8��x�� ���3w��w��do������6G;�J�	�{��K:LD�y}l��� �����;�7U�;C��a_"u=巍��+��j2I.)��{�c�D�8C����KvTLuL�[\����2�dĢyP�ê�lyY[��8�s&����J��A����d%HJo�HW"������K?�s��+��+Ǥ�ߤd^	Z5-��H˙�[�x��s�PVa�`_͎N`mM$�0�?�����Xr|�>j��h�+���L8(�R%���׼���V���=�߹����H�9h9��R$�w_r��G��|31絈���~�s� 
i��,�*_�+w��8.��b������+�3�������X�%yI��F�f�`]�����(�9������ojQ��R�ы e���!J\���o��7`�4�W�״.8��b@���-���θ+ �8Oɚe�3�[�.�2܍�E�e�3_�]��r�{�H	��;-��dq�Ҫ�k�u��u�c�5s�^�,vcCZ�F:��^/E�$9�Īo�Dt������n��)^�Z���������iKp��~�%��-�O?��sS���B2���P�(���>��k�����4�]�D��-%xD&��&�#�0�4΢�c�p:����V���'㽺dow��
g�1N_����6`����2y�P������i$� ���� ��+��cc��ꦰ���c��U��'��b�ؘ��|K��G�n Y�o�q�5'�$���C@���x�!�E��dJ`K�&��3�MK��{���G�x��Rf� ���H�2H���&i�K^��/@O�p��F�uB�Y�9���׉3��rni�?���L�-y�q3����=$�.��F���5�Y��䴻���0�`z��+a�պ$�x�pq}ȷ���7
�`����Q���q���SoLتeb��-��8W��`&��&x��p[�hnV͆�&P$T2�'�{b�b�ޣ�5�a�  ��GZɉ������\�L}�WЏ�#�m�"Q�w��� �F�C����'�"�������B-���K��y[�Lчq:Q�@�)}h��r�M�)_CWg������IR���N�B^��A��8��
�}�"�f)�(�a}"�H�P����h�Z�O��:�kQy�Ъ�v�y_�{�j�S����|���m��n\!U�4>�޻e漿�U~�HG+��@@�ֺnw�>_���պ���ki�X�[) V<X�}7@�8�x�w_��M�w�w61�R����`)ɊCu�:��KI��Qr�op�*��tE��>׸V$���i?��� ���w�e���z��׸`�m�@�{!a�e�,��uS�N��Zh��;3�r>f�"�g-e����$�?fN�w�ʗ!*P��+Z���d�X#���W8G���=O/Me�FI�rA)n��Pgn����1��)���l&}���
xqy)��2��-�����p�,�	7�h���|.i��n	�Êr�k�I�
/ͬ�51��_��zIl7ٍ���҃?�Gx�q��Y�� ��lb2�= |�''�c�C/�f-ب�Z7\��J��X57]�$,��ŏ�o�����ֹ}x��.��r� r1�C��(c|ic�]Q�1GD�U�1�)����N�bXQ��5*W�ے/w�
����yPB��������6\{ntg����J$n�;�fKoa爴��N�/k�v�?Hb;��'�wl��p�͍���c,�����9���l�7jY�12z&�ү��[&r/% l<3�q@�.;S��%�C�kb$▁ j x����]�rv(JY�}��݂�O��uށhO�M�%��Y֋����%4u���ZLO���ה��qघE�M��x-�/�`�ʤ�Kȼm�t��d�fRv���>~��+�HTS�&���T$prK����#�uoC;��Rߙ �z��y!�R@�u�h�B�[5�n��1�w��bF$��u$G�"�(�+�ky�r��-��0��K�ۺ	UCvs[6�0���~�&�ϭ�:ɐ����m����>����p��g���;�-�.���� }f`,z����e��7�,:��.� ����N���j��#w�K���!�S��cv���no�Rs�ί1�Ä�*6_ʻ.g�`�)�m	��W'DU��Y��׈8��6.,��{�UΗC�A�N�����+���� r�Q����#�цH�6�[�{侗�-�QL��1�;��Tn3�EX�JF�ͼ;���nxt ���J�A���w�;�n���pt�>�t��0ǄMUy���|Gl�ٲ����C��f�.]+s}�?Jݜ�j��z�>��M|+�����$�,7�E�@���~������
J�79�&���$7��t�� ��Iu�ζ��6�%=���A6�l Λ��
%�v7�sNݸߗ�0��UD�P����7��Ό8#o����bz�����?/N�	�5�hc?m����4�:���"��a�S<C~6�I����fҨ�FO}^,��-{�OS���l������Ydmu��O)��lN:���׀�Kbݚg���ѳ8i�uc9�W����$;���ږ9�C�@t�Y{���;��t�c�i1�"6�H�|�2m*$��5�P��G'�U*��������a��ݤ�>7QA�B��1I�3ɲ���?5+9�������f�II�@H�t�%1�ܓ�s������a������� ��X\ñ���n�s{yB�7I�g�V��B�h��G�� ɐ�=�mT,�.^����C��E�EI����� �l��?���J��?�k�N7h�<�*=adnV�k�ک	�Ǟ@���z(eD7ד�A��{��9�����v+��4N����0�A�}�!C�����w�ӟRX�e��}	2�/��}�S��V����:��ZV1p)D���D�T�s��ŗFV��Na05gB���0+#I���͢�)(k���і��y+^	��G8S}�^�s���*���F��a��k�152�-�#��/ؠ+Y���;Lc�7ڙ��ADZ�TDJS���=�Y�}>�.�V�*��~$�beKܲ��f�g:=?ac̭��� ]��|\�o�,���8���}���T(~���N�.O8�ſ9��gs@T�I�Ӵ��h���◠��㎏� ��=�����2�"KE��Rż�xV�`W�ۮ�c���S�4U�1!��}Ӑ)��9��o�Bb�}ҭ������A��LAws%5����6�^HN'z��+�+�[@�\_N9���S�vP|�	]�OVQ�fBM�?X�&�����㴛t7��O�3�GhW����%K��yg0������eJG`�#min����c��	|�S�M�K��L�M�g,`�R.��{�5J�����SL.���;F�~���6��&1�2�=>R�:��Hf>T�s�-��k<�$+�ݨ�u��j��x�:Xl���	��zd͞?��nK��k��T^Aogm��	�cfRYJ�ƍ;����b�uym���k;��=�4"=+a�IG�P�E��k+��Λ�P�]��r�RX9M�n]X���!�=:�����|!̈́0۶,� �����K�Ͳ���'⌝1�w<�����Zz-�i��(��C<b����@$l7�l���[�_Ml,8�\��,�Jh|�D���-��y�u˼�Bz��!����P��?�"2U&%DI�vN���@����K���7�s�������� �� �F��劤"���В$Z`R�>��I�Hu˃��w��k���|XOd�� �`���͜S�`O|_�cy2�g���ɔ�|�:/B�;m�����l���cI��Ơ�o���Je_�*���/���C�ȻՄ�P?���Ju�Lj�wI�)�F��?��n8kcC��x$���AaR�a��\Z$�@�X_��6j�ތy��6u��ʤ]�vw�?�;�*�e@�d���v�pl�8q�����U5n�
�_s(\o�
�X}|om�2�iE)���+m��jH�� c���]K��O���#�߃|g�v��,�e�E~=[����ѷV��r�Z_���u��7�-A��>��� #y�%�G2�3T|Z��hۉ1*_N^`3�*�`��7�!�x�� Qii䣕a*�Y)�^;Ŷ7"n�/�����:}�*"?� Y`1�B[̎"�[+z���S��J�a�z�,�(�{9�������GA���Y3��֯�[��c�����FǷ6�a�Oh͒16��8�pZ+; ó�#ڜ�(A�k�����$���F9s�@E#��T��Ңr��E"cw��f���n�`Rf��7��t�2AVw-�2�_[��q�ɔ���9��0v�J��@u&�8�R�Ha�{#��|� X�]Bf,��3��/lH(��1�1�V� ��ؔm�E����!bB|-����(ei�kTѺ=Ƌ�"-�{Pq��J�C�z���Z��!ޘ�Tl�]g�+B����m �lq��_yC+�����N��_�D��c΍�
O�LboHUx��Y�2�(8w]�S��4�A����8�s��V}��һ��B��cd�+B�gMV�,��2G�^�]>������4���x�C�D�u�7�>�N��q��rgƀ��2̫(V�&���<��Og)�Ɲ�a�Z�b�H��NL�����RʽA���=��Y�Ӡ��L6��|�O���(3[�D���|���=j��M�=2�1�v����qWOK�g'� �`
�U�2H��(uz�t�����盶��I��3��mE��.���j,�f-�D*�|�����peS���?*��t��d�0�Y2ez|�c�5��Y��~W���������{[w��e������ñ����m���ـ���s͇|����=f�"���0�G�4>_\���ب�O�ȡ$��^��8��:
�`HH7m�Q�l�	��n�peo�WJ��h%A\�<��ݴ���,8_��`�kQ�y��u���E'�S�z*�U��p�v h�(r�#���3�Pq�L݁4���Vy�F��j�����I�ѕ��mRr�W��/�͜e`џ�2��� �ͳ[q�$����𳠱��,h/��O��.��'���t62���HEy:c�� p��/#5r�X_B߿�-j�>�]]�h�4�۸�t�^�0>#����k['���s�8(��2���b#$� ���n�O
q�V��~���;�I����Sld:Y㑬� ��m���_����t�p���*,���e�,�/��U�5U�G�`<-��G�im��z�?�}خ�G��j2pUGs�h
IN/NfN�k�.d�)#����'}{����d`	;P=L����<ĭ@	��� ��!aw7ʛ�)�w���w�'&����(w�HP���)D��f���n3���?� 硼�H���5-���]��^��$�ئ��_�DC�e��ѿm�q.��5�IR�Q�sD�AZ�A"Ʒ����y<.i3��לi�T,!�3�Y�p���+�C�磘Z6#>�؅����]\4�(}^��f���;iǟ	����ʝ�%�x_�X�z�O��2�\%�������.�g����Z��i�+��e�b�����k��k|���^"}h�ڔ���!�#h�V�I��@�ѫ��`4[]�V.���c���Pp�3��6��s��D6��NZ��*�d����KU��TyS^��GB�>��v^�ϖ�����N^:j6�7�`�wǟ�H1��?]��<�k����A[�uBd�M��"��,?��"��AL���_>������f�X`I���r�x4�\Y+���"�Br��B��d͚�9\׍�"�/;�O'�@.�²۱�E���S�:@�ωV���O��>�/ט�Ox��}��ƟcAa9]��F�3�h�^d/b�G�j�}�0�%�����)=��$��d�X깠�\Z��c�=��<���}Fܭ�b��k�:s�s���6�N��s�ı�gW���C�j��H�!�E�}������� �Bg��mF�3�`x�;R�o�ˈ&��ۏ��+ ���A��e�a��� �Oe,��X�"�����a�LY�	���If%x�\5�?�������z���ň$�UjߤF �w^�51��(���H�0�;�#���h"�&}�H75'�*��Y"�O��lx̯��$N���H�c4?Hd�|�F�_��i�ß�p_��[CB�������#�'��V��O���ԉ��&���ÊK�£wye��1\�������J���Q���k��@G�$}��^�Io��$"9(�9=�h (d#ٶ%9e�N��~,S�G�J��'3A���fR6��PɎ[I��!�-hQmf�`h%~`�]�-؃Ƥ{�����87(y�L�ưkC�~y�}����l䥂��%�	B9W�����P���V��G/��~Y�U�9�e��wQ��B"bֳ��qA��ݐJ4��L��s����JoP��gŀ�����ݟ�!�I��D����f�OQ��Jl��_�~�+-F��t� �����E]���ב���h!�c*=	�!vI+r#´�-e\#�Ia!���A�����+��8��QMa�,�volB��RW�U5�k�j����vu���%��5�@�z;�>[J�4�wX����֕��]�آiQ�\y14�H�MC��p��Tr��D���*r����՝��P3��:�Mqh���к�ɐu���F.Fb?�Mq(�<BGuz�0V�I5² ��v_Ǻ��h��J����_X��v�|� C��Bw=�o¬@I��W��\2tl�6���X�|Y���i�V)���Լ������G��Uxc�g���Q�B+\@���5�3>�9�"E��ۮ����.�u/��
�����	������;���E��mr�j+4%N���	�%������04Q&�LC�洅�%zo!&�\�3�F�U�%��j0Ҕ��i�wh`$�W@;�=���e�(���e��鸬W���v�"����2cC��7�Jk+V�۷�hm��Kɍ�����AJA)��s�Y3��IV��E�]�Э�Y��L��{�q���D�
n{?�q��L�����h�z[��L�&��3(۶���$Q�.J�/;��0x#$�8�m54�d���H�uHooN;�[H����U�� �T��������e@�����R�r\��n�n�����e!�a�i.9�)mr+=9����hܰW��ꢶ)î+�5@3EMో-:���*N�����>��M���aE6�Ҹc����3z�׻��Q���`ۺ��#?�\�مg
�P�G��2V���4�����X1��K��������/���e,��1�&(jI'�PL����c�$Z�a���4F�]��/��`�Y�MqP����b��	|d��t
ܿ��zDV�k�_)�B�5��a;g�b���~����-DN��2�]zD�\^*�6O�����5�1�ƀ��Q���}G,J�ZnN�+@?�"��@�UP��mՔ ��Ip|.t:O�r
x-��swJ�@���9*�$wC;�J���榱��6M�̤WFuj�	��$�H)�(�b��zd(\m	��ERY��1cS��A9���"�m��n^��_����N���;g��)�Ly��[ޭ�e��t�J�ˤ�N�0;̶.�>���PJr���[�nvY��d��Ɓ��e���$;퐋'I�*�ma)E��z���!}l��}�ll�k��{� I� 
�Nh�_�������6�:�J�j.���b�oA��i��1�]>����E�Ч�����3��/�"���G������
}�P�lQ���Z���Eո6>u�O�����M�m�� �9�*�����ɗE�n�d��-�VM�v�����k����>�L_��b�*��u��z��K��n�ν۹?`�Ε����.�4;�0�L����SB�^x�0ma�55h�6y�N�i��gqTҖ����lKef��z��a͟/-�{��gB�M乞�P�^s��q�d�P��i�L�:3ϻ���V�nk&���l�ۘ�����B>gR}?��/&X��f�;�����B%�ce�>)	� ������sQ̧�{�c2�m�jUR6�ռ�7�WO�kFp�O�1�ַ�~q9�6&s�p���� &l�C|©������U�U\������0�Z�
� ���|`��-Ok�z�Q-�A<)̣�kM�b�g'%�%��|�7�\�Z9��L�3`�f��l��H��[ۯ�k��'l`N�Jw�8��	����Ӈ&sL�I��\�l�b��s�~�1D���L�.��5q�u��'�)�69)X˃oPN{��4L��epu h��M����+�w �S ����"�">���D�U�A��lĬ��Ȏ�I���qיuz�=��,-,PL*H�w���*�����v�U@߯�P�X�[xW�4��Y��1�L����@�Ԋ���HMNk�� tj� v�|�J�[�E��po���_���o*���KJH'�e�,��$�ݡ���Q3G'u��~�s��\,k��Y���$��;����r~й���c6�O����qSh�l0eӈI�S�����ț��=�_X��!?����Vbk\��p��|��,�d���,,��vҠ�^-�?%��@gը�Z���u��"�/1$�q��pOZ.ٌ�%Ɉ8��7��]��5hC��S�uO�@}^h�Q�:	���w��v�EaW�.\F(H�"2�Lb����aI!�K��
@�~Z�|�ɾ�4��}��e�/O>����]I��;(Df
"9��	��ʄ�F����h�M�Ok�ֻ��_��Z	ɻ`s'���9�TOU��������ݒ���O{p����@��䢌e��o�����'�=�`���&*n��?���1�`䜼��N���|�m����^�y@%��+�?k����	�oQ@���ɷŎ�rj0��| .?�W����h�cx�Qi�!�rf��wSM>��=T��������l��{(���\ŊpU"(�����}M�AD����C���a5���a�(����r�C.
��i����27����}R�3(�
�ĩ_tM����V���a�(��(w� I�D7��F
�h�ٺg�'�|��F��t��%^C�9�4���k@˔
��5�rI��
>��w����ˏ���jqc8���B�84pC)�f�/��m0�I
���/_$�����o;=�d�',Ζ:p�J���AV��g_��0�N��6�:~?_�К��l ��´Ygd�T��h��5�� �I��d�#�f �
)ۖ��=�1w�U��l��qq�>�IN���(d��k3�~��*��,��IUR:;��z.��ϥ���͎@1��3����;�x)y��p�Ȯ�����E���'R��o P��@�	�)q5]zW�|r�w���/!��=jj�c7o~FA�Ā0��G�TU�0�<ɏ5���4�T-�l304Q�x���mǨ������|_u��j���ay����ݻԚ*��;�~�nK�2	�v����W�ęE�7��]�'w?�q�3�m�-�;I�'��%K�,yAT�϶	�~������%sӍ�LJ*
��x�b�tz�1D.�Y��x�%�"�Jo�mvr.�3C2��ۋw�z����"ڷ&���$F�Ӊ�U-�~�[�ڮ��sO�Y2 [Y h�4����Ž�s��bc�fd�MD�l/����L����σ�;� _S��?�~��]�su���Tb��V4�kKO89�������M�����\�����_�T��� n��WKVM�A�t���/��}$}Af}�Ns�pT��.�G���a_@�>����;�ژ�����
̫���S.�f�/_�88��>V�;��b�݄8�'�6Q��>���=0Zzɖ/ ��}�;��r^5[1D)k�� ?m�sw�(�?�~�u��Ź��$^�a���_�uц��N��� ��FJj#ݍ޳S�_�m3�l�2�Hȣz�@��P�B�ƌH�%y�����q?�"�iщ@����|-�qȔ�ElҊ��K-���E^�}������g�l�]&����1E��lL�(��ɚ}p��JB���m>%��T�c�����K����9zj����ˬ@�S���T�}����>�m4̪?�aNN�Ո�a�{�����q��z��p9��ù��R>R��kc}��p��|K�ٟNuV���fʾ0� �0�A��W&�Rf>���	:G��=��s3���	��$�`��DKb�2Nt�t�K{�[b<�S��� ����Ĝ�$����
�^rݬ_��P��֠���f��cJ��XN��u�_�yH{X	쾨<(��0�||Z�r��/^.؆#�~�DW��e]����"����mL>׮s��K��de�V{��=����ϡU���C��>[&`�� <�(�C����������6פ���/5��P:��ɒ{����l�vT*ΤK�oTy5��g��YXyS�%�\�굳�2�ttF���я��9x�v����_�b���Y"q��w/�D�Z҇j�K�<�3�	`ӊ������V�N�f������q)��<5�Y��k�}�|�Րtu��	$�%�'>�Z0L:�f\���dҭPHi��|i�_�sp�8&�>p�Y2e�u+���G�*���'���M�k��{��o��)�q��Vh����V�Ə�[8�t��f����G7Bc�g��0�hY>��푹�l|3����<�&��H�, �=�=y�I��.#`Q�'Eo����4P�ŋ�k�m�����>����m]�.e/#�r�a` ���Qv�wm�ݦ�p2��Csb?�v�Xm��{R/����hx�:,�.J����qо������4��K�YP�
_g�&��� ���3��D��.��|-�� ���3@}]���R�6u6ڬ����U���m���əh�lh:tP�Hj.X����窵-�# ��߯Qz��u#j��ŗ�B���g,�)�)�c*��Z��7���0�b�c?�0����y>8��� &��̈Q\p�<]��_����������ډh��D�h<tl5�̄FXǸf0��Jx���%��nġ��`�b	`8�0~��^$P�Y'�]C�~�
ߊm^{c�����I-��03���Є�Z��p���.
�a���DZT$r�7���9�?��n�gc6Τӭ|�--}�Vj�ߴ��t�u����@���>ݙk@i�M>��r�$h��K�Bzg��ڦ� xظ�G��-��2��w���e��1.$��tg���/u�u����6���tW�W�$(�ʎ��������-�si��rK�:̡��Ni��Y�Z�\���]B�0��GJ����oN=呶ê��x32�quK��O(u�O�ߘ
\�#�EY�>��n*�e����^�N+�<y��?��4!�"*�*���:����{�h�_@��!�̓[�bqGfX`׳H<�?3Q?��x�N���1O��S��6
<ʀo���,m�c��Hֵy̄��*�)��T��R2�����ɚ2#sӼ�M�ǲ^>�w +�uTZ�>�~$Uz�{���!*�� K�L �@���)�:�_T�,�]a%���j@P����G�Bk1?p������A����C�d$9�Ş�HF�N�4���K�/�u���7Q�s���Pe�������[J�A�i,����@**�22Ym-�,q:�M���u�vP��u�C�^,���%�<�OW��|2�����3��X�f�M��Y����S��jFw�G�'�ΜXECAe��,��Q�ر�,������9y��ute��3�5�!�y���([ܝ����m	C_��� � �i��6�H��qAN���N�����s�Y��?h��ʫ�%�߲Q�X@��#[���O�6�0��W|����,�u�u���>]u�=F�]�J�QhL�\4%�=?� ���{#��A.�Z4ӓ�bN��XPq"�Uэ3���aA3�~��76V�>F���FX���)e� �UE�o@2�C�U�0?o�&t�A|7շh83,���s��*��N=7÷�/l{��ҫ]���M�73:9��*����0˵��Ge��^ݮ]~H�����\���}���YaZ���S�a�z�B=1�)>�H�8�0R�zw�d��\�@�hqTh�I&
[���w��:�mF�'����3�b�倊�0k;��db���y&*`�� B2��:ƲFA[�u���f '��f�@�� }� Z���;S�s
����7"Am_N�M�kq�Ii��"ַ�������Ʊ�r����$�*��
��$Ӟ+Bn�~�_�G��}� �����C����|TMI�@A�up��]��*�o\��1#�):��淗z �JG-U܀��H��m�~?,,0�cM�N_`f�r �Z��T���	g�-��2hD�g�����j��[,�N�i�L��Tq�S�n�C�H��\��+;Q�A;�	~T���҆��1���D�{J�b�����M� �R��s����. a�jXG鰟C�&���-1�n���/�+;�s����bЌ�ȱ�bS��AdΉ���[� ��h���nĹa�J�] 3qϕ��td{�����D2���M$����֟���Ĭq���*�2&f\�N�F"tV����b�l4�AOCz7���2�Xk�9	�;!%�<�e�ڌv6���z��K���ڽ�(~^
��#�I?�R��2�>|�؋�t���� �塾\-�w��/���V�5Ww��a_U?C�&��Ly~;=D���3i�4�����C����8���#���S�`�v~4=@��� ۮF���UHe�Yjw�]S��|n�ݽ� �dF���<v#���m.��]n�5�zfǇۼ,��#��:���1���Bh&7y�K#6�NoRO,�hRϓn��Xd��P�{Z�j3i��k$����d~0��N�mƎ.$T��C(�X���<p�[�4/p�v)�C2���S-구È=Y����)LDŨ�Gp|)�0n	���r�d+�K�p���L(:�j{��Xz3x���e&��	e"�^��@��
�;�%V�H�Ɛ�2�r�t�4�5�!;H'�:)��61���S'N��s��ZAp��c�v��1��@������.���r��K�����~>��d���_�^�5T��p���<
��ǟFd��T�
n:*�2Q_�5�DkED��{N{�]��ˏz��f�,|~��%mDGH��|x�*��{�Q'��2�c�a��wCE�樓��o���`Ū!��S�!��e�)k�f��ǵL:>�G���<v��r�@�qPD�o-�
gEdEMB
��fl�(1b�n�y���	�Ma�iO�1�F�ܥ���V ����#���)�_��TvI6��:�8��g�>�%S�������^F6�-sC�'�F����-4;����V2*�)�]���b����:ͨm�]&�5-�T�)Zbd�4�=,���	�P<8�@.�=�.�! ��A�:5����ð��Z��ߛ�`f������k\���k����v�	ʿ��di
EȬ��F3�k�>�'���؟�D��w���G�:�#��f��������<��ud��X4�+ԂY�&�[�����W�e)�a8�y@�j$4!�R\YGt�p��7�I�V��$��p��F2��a�7�!�#^K\�f���� �Cm\���*2��W�<���%x��*�D��D�3�!��a �����ҿP��{B��g�sNHq��O�k��/*�V��������]�b�7���î�}��:�w����|u�q�;t��}�&�9M�D�;�*}��n&/��=>�)	��@֥���p�c8�ni��j$�<��pձ�o0����NŬZE,���Ag �UR���2e"�}.���JF{V�7�G����(w��[]�QK}�죀�
3Y�����w&���g�o	c#m���>�_��V7�sO�6#ܘ�C�R��,ڤKI9�f ��:(��z:��E�LP���r({Zy|�5�d;�0�6��0=�\Jo���U����rֳ��*h���	�$+��X��$�j�z)��Z��?�m�����Y���&
M�uD�������\	{-JB,%(`���x��%
�@����?���p��H\O?UI&�gO����]I�cs�$�D}t�Q^��<cց��׻�}�M[@v���d&z&5bٝ���-����T�S�� ��H�me�����JR�c�]#(w��KQ�q�2�z8
3�� ��@��LrU8�����T�'���!Z�n���4.�W��}�რ#3���߅:��s�cO���5S���>�i��D�Eh�G�O�0������� ����2����%E��V׽9X��nL�j�ެP�I'��^9��l5�M(?��ܖ���F�������h����s!������*��"�`U��6)o2c'��������u{�'%�A�_f�_�=��|�!��1\b�g�Zw��qǞR�71V|-�7�܋��7y�B�lo�AH�*@1E�����/@��T}"�"/��'��4/͋O9�a��=A���c������_����z�ŒUp�6N��s��ψ=�_�����dҳ&gi_��X�����ŧ��x6�IW�Y��	��A��ә���W�ȕӿ��Y<��BP�;T�kj�秎��K��ϋ���K���i�T�=u��2#�V�f�)[b��l�Ͳ����}
��1���fس��kA��?NMa��_�4��}ѐ��}>)ʞ�80�c�BwZ��GW#���RGC���t�=J�	������!��;�!4M��Gr����Q𢁶iy��^j��]�%�dOD.
�ie/mq�e�˘�D$�pߖB�"�%w�j�׏��ς
�M�����l���� ����Iw��W�k9���!܅e��R���h3Ym©�3�0�ސ֫�b]z���1	��弿������=E��坦9��[�g�~ڲ3L|'� t}(@���7X�r/b�Q���a�P�"�6�j�B�Q�1�3��q��i-����>�l����2���n7��Kn�?��r;�v�����F(�qu�t���y��;�07��/��)̯��s��.4a�jw]#�T������L�����yZ����'|9�qR�|i��C�ћ}�tb��!�)ӰX�:��G09�}����vq�!Op�4���<�,/���\��P�Q�%B' �#ZZ����몋���J������&qi3��K��|		���?�wP�*��b�B�%I.�+�a�o�I�S��@�ќ���������9ު�V�TS Ġd:�Ѕ�VN{w9��ŬE���b�c[\�M�ƭ]!��q�l6P)�Eӏ�o��&%�Ƹ�q��%������_�
�:�T��Ԟ���O����mMmO��m-|"����9��#mX����[��	�C�P�����:J3 �6�g�#G�5�e�T����n���%�=��,1�(�`���FJ[W~��6z6�I�����Ne�|nR��^�=J��F��p
� ô��9����Hˎ��@Pg|r�
%Է[n����P�A@���Z:�(w���]eW�v`��W��F�:����@�����Um,H�!R��%��c[�����GKv���S�4�Rg q���:<���?*��|��p����"Ҹ0���M�oM�M�$|0l˜��%��U��qA������gݵ3�Og:�3EZ���x��q�I�ME���/TH :8̺m�^��3�a��[d����L ��Nb�KM��$�V�l���G����8�
50��Z�' A��U�e�JG�A�"-�ʋd���ś�=���5�V��.����%TD�[:��7pf� )GSh�z�h��\l�[w�^.R��\e>R�@��>N�5!�{���
Dd�D6�qblw08����L:�Ѭr,M��E�h�ivE_}�g�mᐥ9�33��w��M@V.7�kڅs8��S�n�f�Q��	��>{3AJGE � �B����]u�/�UU���ݩ�)Ԯ(���-w>sweX����ki��	��j��o����ب�}�x��Y��>��9qL]��W�bQ����Jk5f�w�z~�e��k%��T�=�3(���CrU��p�Hs�P�H+��!�1�<���0E�S7�v���8�e��N�ّ)=Ua���Ng<'�H�0��C��U<�8t�������Wn����҅|F���t��|Fxi �����ԭѿ�V̽�zL�
��Y�`X���3	(�Q3�i�<^�G⡃�Y�|y�O=��ky/F�)ԧ���pcV����5g��T��v������ی�҉;����*RA`��6<2͌F_��%rB ;�
t<�Ѫ��P����
/
�'��:�Rm�H?��H�^������x��X
vPa�Z�޿��KŤ�D��_/�~��.�����Zc�]�1��^Gi�>���1�@"��O#D��	{�ܛ6:/-sQ�I6A=]e�*C	8��\h�tї!����H���j-��N��J�^��)����t"�_A�b��X�sL٢)��'�H ��9�
�R� �ι�@~%��A9ϧOVu|b�S�=-H��g&7;�<_$i~i^|Ѱњ���s��2�~���^���g�����*(A�I�hy��?®��{u��$�NX��çD:h��r���k*�[���k�$�7U��zoSZK_�Jw����+�"�c�?Y�7}��0��@ǌ��E���������*��@���_��ӏ�r��<aq���Nu���L����g'�i留6�,�EԹ�̾����Ft�(���j�/���۲�_��A�X�N%şjL(�/3<X+�љ�Ώ ��G/���n�@������=]xK�R~�������0�wƮ�S�ܕP	V���+��oB��,��ւҳ�n/QO�.$Se�M�5���s�e�.̢DpM�����1����Ҏ�k[+ZA�������Ag��?�n�6$f4��R�'�nt&�,�m������V�@vپ�K�!)|$���p @v����Du��6U 4����e|�b��YL �:"ڦۏ���L ���gW����7�m���q?�J��Dcb^��7���Z(�E^'I���З����b�����qM|<��'N
��-JB�a���C��~jY>uM9N���W��?���T�%����w�1�w���~nǾS!����uE�F��c����Q̓��}�����*��M�¾:�~I�g�4���P�Eo������ȏV%����<kRk��S�b�kɮ�!(�W�-�d済�WeC4�?��J(��4uD�r�N�����Z_�B�@����u]cD|�x�q�A�����8
��݄8��M�ߕ~jsӤ�>��(Zz���a&r8��������o����ԎE�P����.�o�/qh�z���t1�<-��'s�n�(0����l~_��X��f��.�VVk��j͢�j���b@T�
��I��<���W�u��R���osСW��Xʽ�hfBnZd���5]���<��j+�{��w��w�����E����^'ag��K"�mA���R����W- K���6,X�)�!���1�"��o$նZ�pp�t��(��x�l������.�+w�C9����Ҥo�
29�8,������ř|��4��<J��	l6 l��UŃ����TVF��U�ެ��֏�\M$����F�n�������.�D,�z%�.�↭_�\�%ik��%'�{�$����[�wL-@J߄�|�QJ�eb��m���c����$�w�n�Pu����F���a��[�-Iv8��(��Z��$�+����։2�<d ,�J-�0�Ԟ���D��9L6�F�nM*�Q��ܤ���`���v�4w�"w�Uh�X:^'L�[K�Y6�=��ZwI�,�ð�o'zd��G��Z�Z;����b��(r����)&��e�)f��r���R��u�향tJ�n��������,�;��.56�d���ٓ?�0���H�R%��-���� {�Y|Uj[ ���'%��O:ơùcy}�*���w����?N���[<�M ��@L�fL��/b��+����.����a|�?`�,�s̊pF����� =��Iyf�<I�H���^�Oɵ�uǞ¦�[*�Þ��R��[�r�1�<����g]l�P�M�����8?Le8�ml�S��c:t�ʈr*u�S
�^�?��97�}�֌��"Q�����drK����ra֡�}�tT�oK���o��&�K�^ݑ�h)H����!���[@U0�mM4�f���L�H��Ρ�{���dº��ּ��B�&��oRjJl�~��S~�p�0�`��[X�V1��탉9i
�J>��/�[�e��L�ԁҹ��3{�/��H��I����P���/<?���>�-w��"�cG�����Wqm��T�xpC�aH�C����8���\`���J5�J��'89�X:�Bܗ���C�5�nAOހ��8�b��l���Ƕ�;"��w��In}zW�G�k��N����Q�h�gѱ ���(3��%��	u���'yU�6�S�Pw�A��L��� �1��*dC���%|���!a^�Z��`b, ����N��>JD�y��l? ��p�p���aCIhm���o�%���9F��Sv!�흦��Ӕ�?�U���P\O������!��B�(�L��!ԓ>�����}p�g���L���m���?aK��ˋ�@�>s�bLW�[_
�1<Uݗ@@�e��p�L���{D����M�ȅc�a���K�>�F�p��j��6a^֝��ᚰ�9[�"��+�5��&ɇ�̃y���͈o��;
@)n���f�7�m�f�f.�L0����V������V4-~ ��u߁�E<4�ת����l�E�l��?k	�R�w�F	��C����s���z��@5m	�ry�l�j�b�K�]�u������f�"Fm 4�h�k�(���@��!c�C
p�h��yS	z��Lo�\�2q��GK(��:�A��lT�5���u=��7�'��Z�����z3�h7��nA�LH�t����x��H�j�Nۉ�]��/�{x:f�VI9�։���KI����Ήj���	U&����{�YK��J��j�eI�H��#�Z8�n m�'���C�e�1U-u2F/����S��
3���2�{��YO@���u�^�[���Z�E}�/��̼�삎�4�YX��GYj[B�pWU����-N����mo�ځD^�49[�NkX@��ۘ	{��P��������jpL���v�< ����b��2�t�L�)�G�|'"�±D��/��i���*"-S�*D�F�,�a�������S�f� ��P٤+���%�(���o2ly���5 �����ԃe����b=�4����ѫ C�7�Yn�$u�Od��Y��K]F��8!t�(���Z�E�H#`՛��_��B4rP,���5�"j[��?J硑z9Z��:r5� �;]$�L�L8�����3�W4>B�i���_�O�A�	J��+�/���CN��;F��-�꽈Q�����]ﾸ�&˶�!��h���g�wD�9V2Bn�=:+R�J�4k?����>���yM��κ;S�o�Y.]������]Ѻ/λ��0E����=���Xh����5ʃ����efp���N�X���E6z3�b���G��9rrH%-R�Q�B��g��s�+p#`�Zl��i���雘
���_`�x�m�;^4i�Ϊ���V��]���cW��P�C�ٲ�}
K��@o��)El	2�@2�ƪa/�d��k-/11Ʊ�δ(rC5��[�[�6�o-��)�t�W:6:�4�X�����A��3w)�:��Du�p�t�V �jG(D��-{䟚�3�Ɍ���C5��ǥx����P=z�>��wdi˳@^1�|f�K��:Ka�uw�$q\�o航�"�ό�g��{wjS^ų��
x0�ە��'a���ٶO+M�iﻇ��)��Er�/��3q��)t\ 	iw�K�}�Vr1ֈy�����em%{J���8k��H�j/��NV���iG4���	��}#A&pF�{?,�l ��:Ľ��f<i���tf+�!��}��4��"v��P�3��)�(4 
��}���x:����E]z�F��ţ5p<�i�9�MG�#,�Y�Җ��]���I	����8������T/3)r��.ر���I�2F���!ri�ђD�E�J�U��`iqy~���w���e2x'���qe���;�'r;P�|�!���f�G��Y��?��*+���
�Q,� ���Q�4n�©��D��!��<^��O����]��:
�/]l�+Ǆ�o$�����S
�X�����mF��i�@V!qM�R`�-?�$l����歕�C.Ɍ�pq����DN-(ς����泋AZ�Z�g�|���z B{;`ƣ(��x��M/��,��m �<@ek��eX*�����Ɠ�E��ꎯ^vt�����L���j���s����.3�z[�A�&�{#�z|���1�z
����f%�֜��}>D�DT����)�������GQ�ω���L-gA������-�d2����u�j#���Ϝ�ӆ��ik^���HtNxEۑrngU|��߀��YV�|�yb6�]�����'�+ozÝ�d!�W��'W��G|˧����Ai�Y{�0��������^�:�ը⒟UpH�hyEb�4�|�T�y��9�-g��d}�����h0Rpߍ�ן��{$qy0⼹�3���'j @;��Ͷ�#nfv����������vn��Mv�Y�u��"��j�MW�̝��-���DN�ko�lR^e/��K�H��5�#�}P|���
lD �v ��R��b�cK��g�+ϚM��bSs�[���)����lG r�0����W�J>���ax��&kx�?���TG�2�!ZJh|���a���s:����L!i�z�V�8����(J��Pfc����(jT��I�;�XѬF�w�tƺ��������c��I�Yh�)y��e���I�c�����w@��N�w]��r��}�����C=ꈫMDm	TOh�iٸA92{�#D�uR���6X��Lh���ȪR�㰴�~`טT@�6?2�*���Jֺ3{�r�ۅD��Pc����F̻tӰ�O���9@l�DP;F��:����.��e���\n�Ns<!��� 3s�[���*.�����0�9����p{��4p*('x��gt���#�� �������&�»?��;�JizKb,yA&xch㽑��A�A?�Ns��z���p�y�}:��>��Ha���:��w�ZZ�M0��γb�(����=�6)N� !;hL�<�OP��^|�6L')��Z�!��~j�7sw�fX�x��Pb�-����Ie�#k�FiL�.��B�D����k$�`�U��a�����?�B�˨�C
�r�=��"���#��Y
	�����0v����E�z�~	KeW-0�*?�4��x����\b����B{}0���5�)��/{t W�ݪ�-�z<l&\�dtjص��	��ȟ���gPLt�=��^�����P�/Tֹ��py���S/J�ͭ\X��#N�^x$�K�d��z�����$Ad$ c�>0��+�D�DI��x�qP=q��q����x�KW\��z���Ot�^����igޅW=�H{�>~�6M��T��B8������|��B'�5�k���>&ڄ�Yu���H"���?��v̇Z�C��#�x���v�ٯ@��8��{& +���r���n��i6�c�����hp�s�����c�#� [�,L�4��c��9�iܰ�6����Z{��׶d�����nE^_����-ՀvK�:Q�&�T�[ٷP럈�)��q���.A9��DRuu�DDӜ��H���_��ĕa5�t���`�����^I�/��Q�T��1~�.K�'�i�|z�KV�Z��4�"��Kne��	����$\����ne���E� z:C��c�f+
OX��"��Q�e�;�d4<p8��_�I{jp����J�~�-��m9l�,-y�W=���KJ���.4a��`$�w��8�[������u4��Pz�@_]у���R��i+�{RD��p����T����P,�48�8����8����\f�$|��M�����?��ϣ�@(=M ���,���/�}�Ї9������i��ػ��h#�v+�f����M�~�5;/W���ҭG��rی���!�r��8�l���佨E���$�������Í���Q7���0ȏ�R w�Z��շ�h*���bqj�x!B/�7u���U�]���bdp�#$��B�>פ����P(~�M*��� JV#�2�ٳ��g���<��y7��JVv���˾qy�gP��+oW_�U|&}�(�G����8���f�߼�b.�+j�O	�t.37�J^�pEZo��<9�BH��MK_���&d=�.��m�����̱q��ѡ��T)��/��^%�W#B_����8P|��%[$�+�d�~䜩'�m�<��.*�~��{_�g�C�LF4���_z�V���<6ξ�]�@������r�g�ဦ9#��SM�^|��eIr����I|$�8H�u��F�2�����;�C�zg�����Ndn7���,���ځ���,�c>$>6Ť�2�ݒ��iO�܄������%A�m���by�G�&G=6�����bmƭ�u.Ҍ���P��m{mz���gN��Wr~|[:��0�&��&Y@l��f��O�yaIw���uc\ �c�F"r�d�2ɰ���X�I����̀���:�H�� ��N�)����6�����CѲͧ~�����<�q1�^���?W�w%	��}�$gB�xc�c����:*�TV����J" G�Xm�ܚv}^�Vfu�!$��C�>B6ŷIs��"��S/�9{[��*1�%s�,\Sĺ�yS�t�M;E���	(�ERnT��=�;�ݰ���T��`�0�+FO�]�(�,jzѬ�
��P6���CԜ�Y�y�+���N�׺kc0�$��I�rn�͈+��\_� a<D4�r_�`�xVW*�������ݵ���RR��ѧ��Vč��IևP�;ߪ�JT��/^�p�E��m�v�	\O���n	����X��_���?�K���ڱ�s��߸�������B�[̆B��7��T1�`����@�y��q5 4ٚ�Q�x/y4IsPWA�@�u�1��YWp�)�K���7ѷ�߫:43J>z| Jû�#�%�؏\���v�Z󔊺X x���i���@�
�Z2�n6���uԾ"~�J�+FT@�L�"��R>�ch��Ƣ�Î��q<H�5:1�4�p1�y�i����0��2R�CV��5<�3�����i2Y�">��^p��2� �o	Mu�f�L�{�3��֌�ɣDy��OA0��L��|�!�Z�@.��*&�y)��2�2��~��kEԿK�ż��<��t{pԂI�8�fu`j��"0��;�i|��5RX�A����|s�sL�����;=�r�2>c�c�%q�=	�r%3�-�2�u�#t�ie4�W��q�߮R���͛�Lz[�hs��n+���x�]P�bm���Dԗ�v�h���Q�`�UGe�S��2���S�_�A���AyS3j���Fe ��s-T+y�muJPɋ�b�p��ЬPY�}��gRݿ]��K�۾��o�˥�F@�e�p�����h��>:�Ykl۸Aҹ[k`�O|�K���[��g�U��[9!_����5^�v�>ؠgK�%��r�X�~.�|�!<,�T�"�����#M��FT�*P6����c;{��4��I�a����bR�k�h��L	�Z��OqΩ��% Y�\,����q���(�߉�4g7�ٰ�ׇI@ޜ�Te2�FԜ_�w^�r1�r���*bO77�X&h��l�,`�r��LO��A��Go��^肊�c���Y��Z���1�9��r��C}�%��ȇ���b��w��8��b4f>a��{�{��K���0'��KDdBl��	�bi���o�n����:~�� �g�_�U�)-���J%RI�^D"�k�d��|/�u3��O���
����D%eW�ԓp7m���,q�v��؎R�}X%�)�oE0�Cl6��d�1+��J�|?
t-�:�p�s������ygQɞK\j[������U������p��<$9�t����֪�+�?�:���?$��.�}9���L򊆟i`4�����D�^O״�a���6T�O��fqL�9����>�	���pY��v��fp��F�w?�=�Wn3���%��B"�e�mÿ=��}�n��0��ȋF�Pe�:g����W��i������������;���FI����4ٕ���I�_�P�C�J#IN�;����������Vr��S6���3>�L�\���J�_a�.��L8q	dk�
���c��C�`#��I!���ȃi+!��h���"�b�p
"�|��s�g��h�}��&���m5}"��	�?���W����>��~�����T[u�ZZ����@h�;�/8Ccg�Aj����Á��eH��!VC(rcR[u��@f�6�Gd�fO|m(ćPY8��ǰk(���R&�eo����N-��L-���> 1�%@2F���){W��hת��/�U���S��T�J~b������o=��#-?%��ߜR'�Q�<�K���S�v���w-�̥�?�mx�3��3q4�[@��L���ۻ=��S��쨕�K�E	�*�7-�W�h��ہ�R��"��K�e�3���+�A�N��b?�A�S�:�ܚ=\V:�����g�9�ȗ2�̶�Zr�������%�#�N[r��y���372�5]���DS�`z��L"D�����Fy��y�]�:}�f�	ފ�U���A�&-��@�H�-.,�ݬ/c=�_�zB� �]?���y��w�����o�@J����ٺ*�#�~ই\1��"^�*���c�mdP�c�K��T�Yw��d9n%\���U gu�>�*@��H��2�D�L���gǁ���
H\�jT FQ����[�x�E�.�5��
�Q�8���#=�X������+�F[tv�-��3��i�C�ac����%�X �eGo�j|?�G�(�y�	{}w�_��0ON�J|�]ZM�"�0���^��iE���"��sp~?���J�}$t˽WZ�2x���z������{��rS��;x+���$���[�v�#42�b�cn�.Z��6^4�i+��>�4.��j��&Wd�Q��>6��������8�̨n@� RN/ca��u����x��U٥�gr9ڹe"���P��+s8�ό� �@������d;�[4��1�Ʀs9M���C��d넎�b[��.���P7݊p�l{��u
0DS�������*���ㇱM߈���!������D-b>���A&]��A�R�Ƽ�+6��cD�X��/�q�,K���#��l@��m���,�e�h�N ��'���{n���շ��M�>��_l�&�E��j\D����}/$_����"Y�mC�Ի�u���/����R�ҕ�����AT��q��7r_�#?����q�v����Ϳ��e��Z�[**�Q�!$'�#M�R�gT	o3�e����ox�Em���y��-�H���x"�?�B4����s���ح�1M���8οj���U_�+�\�3���a_[�s�V��5i䭴]H`S
�E�3^�����&a\hC��k�+!��\fyr�ƄB�s������mU�;��\7̂AW�}��2�s7a<Ȥ�
b���;q��]1"5��U���|G�b;�}�*+�2:���z��W�&><7�y���2P%i��"�����5�s47�:�W�KY�J?I���{�3���5% ����x���lO�_�v��@��9�+j �����49Jh���]���e���*
] �^w�渝&8-�g��i��x�+pqZ��}Iؾ�'	����w,�\/݁ԉ��Yt5�-��8J�f�D�z=#Pp[W����H $v�խ�Հ�E�2@�������O
Y�[br�ڼ��k�����m
��G3�p�>�sE9Z�̮���{�0��8�+6Ig*͊{�U�ޛt���I��F6</]j����A0��{��1G�߮��h�f<���r��z��ƥ����C����k��T��j���@cN��q��]� 6�KR4c�D����W�hZq�D��_uhLJ��Mp�-~�A�"�P[S77���%�Yn��{r@E�Q��=�؈��������ԟ'A�k�/��_��0r�!ڔsk@��'�G�+�0#�e鼕��6vW�)� ��}ܴa����O����0!�!����C�tuD�!���Uf�}���t
^1��ݹ�����5��@z�1�A�e�Qp�Oqp	�����v|��,�"�4]WH�Y���-�C���Π�Go:�MM�@� v>:����r�2�LC?�r#��O��N����&%��3��mCF���oXg���٪�>)�`4u~UFr�l��@��FF�y�)�h<`;�&�ҟ��=��/�"Q� ���A�hbE��&�b}z�����^��Lg�p��>&ȃ�Z&�],��n�8/�詵�B�����|�N��N��~���@aD���P+�dn��3+���G53��~�U&2Kt����H��Q+�4��+'H^K,)��:M�B���>tƉ �[���[��g^�+�e�C02 �M�}�x�&ӧ��k~
"{�,_i�;��@��|soL��e0.�N{�\�I�����h�t�P\��s�օ�0�F�� ˀỤ��J}��}K�M2Q&����-�e�A�jh�ظ��fȺ���7'������X'`|�&��[)?u'��v:��~}��.~c��6e��ry8	���*�ENL�|Gh�u��*�&����|�Mb����{���vߥ��X�?�Sp�#���Zvɦ��^Ǽ��,���7��d���[���{&B�71���^��7��*���p6�tf����8��QC�Fd��`��-5_"�q<"k|�H�@�P��o�e�7U�5���n�����!!GvP`�j>��l�A%�K�i��6c簠Cf6*�nf����^"�Tus��j��&����̬m�p�����֭[x5o���]�~���T�
d�����аm�Љ5Xˮy���������~��C+n�����m�]�~R���a>SE��Y�0j�3�gטר?.ቀeP lQ�H|�a���f�&�;��̂�v'�陚��4�p�n��
],N�;�MzFx�ϣ��qPyL�`���˹�ͫ�}2��p��ۿ��F[׈����_C|Cg�-Hc�E�����G������
�APfX�Y8E\��2�+�Ʀ��^t|�T��*����]�a�MψX'?�5�f�LZ�Ж.�����9�>Jǁf�-G�\.��M{��,����)(���P�ő����o��\����D�msE)�7�0�$�~d��!��"����B9�34+p�~�*�����_�k�D�v]?Q��_^4 ����0|]UU��k8Sz�[c���j�n�HG7!��r�];�}�)J�@f�+F&U�����k�7��s=w偔icB�ĵN�Ԋ\Ic���Z��a�fIL���"t�����F�\�5+��A���K�7zC�P>����ީ�����_\[@R�	\����^+�(l�Mp���ҷ�~��=Nՙ+,j��ϓ[0�|N���d��,����/U�	�S�q�m���o�a��E��a%��[r���৭х\��*I�N��)0����U�]Jѝ�b�����'p�m�.���d���� �2�ۜ7e����,�/�س�����ֲ�t$ڂ&8	�:�
��v;S�@ij����Kh7q�<�P�ED-&��Q?�^x1e�j��X"��j�Po=t��^[P�H)��gm�a,2	��	[>��2N.�>���X�	|���<��B@x��D%�A�Ź0)�}��~mlV���O"�ln9�qQ&��'==Mm��S����A���T�v�kg~��%^9�1�>��י�)��3cRDͨ����-{�y��65o:�q� ���&����,��i
�*<2{|����m��V���u:�⹠)��+GŸj�����I��V`㱵�Y�3H����ih؅���*�/����)։g��E$xB�0N�_H8�R��5�m6\Z��o�ڈ��,8�߹`u�zvO�t�a�����_���_��Ww
�P�\��oX��4��e.T��/�2BK��!�1*Eh�x6�w�!�y<��4�Ml�G���&�w*�9�?��n[a�_���s���\F��Id{�P�e�2o�w(�m*#HPm̜��1dA`^�s���ax��/�1�@�����;��e����Hm��i- �	4<t���k+
/��ŏ�c���~F�ͺ8t���:)8����i�h�����^�[��[�3���:,�8�v�$TVƽ�_kXK��m.Ù�e���x�V��8��r���r\K�n���aS�WE�:v�67ghY];�sZ�
���@V@�C��K�hC���u�od�k����躔�a�����B��vy%�5\�)ƈѝ|�	�k�Y^�Q���X��^�Q��*:x�h��z��z4��$Fn����e���&����]�h�Q���c�ŪNwS2G��,�{�a�a�K�e�&y"�]R�&��:��|����s�`��B�Ȑi�]e*u��ng�V�o�����#2D}Ԍ?�I��Z��ɐZ��Fm�ڜ��0+ρB&���j�e]�����Vc�G����U2�ĉ�+nz��,ÖQ=?�h���"�~���l7����<z�LO��Y؋��%�CU���;JƮE���B.��s��v^J��T� �h�t[�*}u�E5Ԯ��������t#��k��s�g�B�x�Yמ��wG�J��Q���!s�5�-Nn�e"ǆo]�SW���>e�ĵ��室Z���#Ozb_��J�P����d�*h3��&�d��X}�E���82��z�6K@m��r Ҩ���5���N�RXټ��F�E�f˂P�jS4]ö��B�?�� �56�ϫ��6� 8J�&���De�f��7�F��=�v�jMl�d&�3���r�� �5�3W����9.�}~�J�^J�������f��b���(0AWB�c����LҴ9�/c�6P�}�����	�c�c�����B�k� �5Vtŷ����Eyw�?	�xr���������HQޫQ��2&&�3(��pA���.Q�؞?�5�x��	�f�b�d��(;^�:]�m`�b�������!�J��);�-E!��#��E�ϡ��<�Eס���b�mTߑ`����͖J�[��K�|6�=�͖�!2��p���yy���ˉ��W	���hݒe���k;�$̆�s݁�����L� �o���~Z�t�P����8�Ow�>Q��sU�Ae����dR��2P?ې�n���)fN[]���B�n ����;\�B��O�W��]�϶���i��՛(��&�l;�w_�11`\�P?U��]��}�皵b�Y��\�.���E4~�Q2)sE��n%i��Q���7T���W�.�z1�����s�5,F)��J=/ď6�T���⺠���z��JeN�Q�H��b6ٓ���9�~0�yK/ٰ����o
:��o�̻�ɝ*����ڊ'�-�i�:���tLI��6�>�A��>��V�Wy%2\��0wK�h�j��R���v�Tt�V`�4���0F�@�:���MRNqoң���(�w<��XeZ�V����<�%�0TtXN�Xl�W%BJ �fv��wE�tp��� �$�V�S�9�E���)ǀ �͒5��!�S�� �'|en���M�I��Q>G�
��ɦV�tU��#-��܌��'>�+���wo�.p�i��h�=��A����p�B�4�W���¿&�wz�Ԧ`�f�W�;� .��G�(���"�i|������]A��A�!��@��f:@�&֘a�Ȓ�9suqrׄ$��\Ƴ%��m�$5 ���qпZV#!���ݯ/&�����s���C�\6��J紕�-��9�`����U.�[Ub�;��k�Vo_%SWu����-�Ҫcg�Q���@��IG��NV�<ĵ�zj�1��t��c�Hx/��O;�
��X8���!`Q��p�wte��F�ʬ�d�P|}�װ>���W��~�ۃ,�oe���6$���*Ճ��SR��{.���4�"�i	Id����(��MQ���A�ɿz��f�Ѓ76�����H����[`�yWtk�YQe�o��^��=n��ޅ�90\��O|���ʴ_t�WJ�.�4�!Yqo)�)y<C�o>=���/���=��^j��å�s�C�C���Cӹu$t�8$Ȭ��N�-��imFT�� ����g
�����)K�;܍�����^�58�*Dc�\>a�\������މ��4ANk����_�R��f��/D��b������7�,�xԼ�l���4�kp�ٰ����|�x�ow�?�NW6�i&�Q�:6'�u�������DL*�c9�ɳ!�s�;�"E�m'�x�_�&z�b\1ԺdE�^���L��1ا��
�G�e7�P�q�E���^ �̩⅔��H	�㵡�6�<�~`U`W-��6�ˇK�_����&�y�?�`��� h�h�:/4�Q �"UQ���+��ŷ��dj8���JP����v%�⽊��]�{�7g?�O�1H�e�ͫ����#�s��y��f�v�IO^#A�������u^x�!p��0�[lio�4���E�r;b���� ^�h�"����q��)���,f*��,�,B8Ty��O�@z�`�����5��S�0\s�P���F�����C�Ah���gGr?n�1ʕ�X2�v#��x���z��E�vĶ���	Η'�Q���a�epQ����+��Z�d���0w����Hɥ,�,[�RG��6%b
EV.td�	ǥ{{� �����2��H�e0�>�8�"�>�I]tU&�K�~;D�Tlӣ��ӷ��[������<l��habB;T2����e���d?B�I��#��O��b�ƚ�I`<�@������
��Ñ[����k$!�r,�����K�v�9T� 7^��β9�����x�	a;
���V�U��*J	Ѵ��m�٪K^T#�����0z�m�������I��R��F�a��K~:y�~z狊��$lȋ���T���苪��ms�(�}����}"�m���� �@iq�b7Dq��'FI��̠%DD{��2�s.�s�l6�c��a��ݲ^
&D����4������k2���	j���>���L�U#�z�uC���MC����{i}�t��ME}�ʲ�,��'m5�U�0';
��e߆�IL����rkgqд��O$��a]o��iJ���
8�o�����`%��`�؞a�$$q"�h����3�B|tc�ɨZ���" uc*�ԭm1<�i�����t���t>1��Oh>���UX�a�R�ܕ$����IyW��D%u�3�ܮ�Q�
�����H��ݍM�W��qN\��8I�\!��aY��`cmY�۾v��W^�a#�e+���k���Q��|�5� 9�^���
ڒ���������Kbg0���ˑ>�Ba��ʑ�>�堎DZ����4��B��N���`�6aϱ;�XC��(DՁ�~H�epﯽX��]��H���+dSt��1Χ��J����U�Fݩcܣ.�ݏ�u�t�g�\޳�uZ���-��.��^��R.l⚢;~d�ǩ�&#�E��,��;}cn�4�;��y�잁��1���U$I�I�/Me�ȅ;%��b^�>߉�9C�|N���kꭐ��K�m�z�s;+t��-�� �u~�1� �t .��שx3����(<N�BZ2�ez�Yh�.��|� �m"�n�	���H���8����� (��T�X�����a�/�#Kl� �u�h�ӗ�0�8)tǞx�m{��k_�n��x�'GL��� �=z�����Z�L^�Ԑc
�_;�_�ꗍ���@�a�u���8C���q�	ŏ���xik;�5��T� -�D"��E�U��Қ"�G�/P��5�t ���7��=\Z=��͆&���	�$�G_��LI�D��9�8<@4����AQ��,Nj�>z���C�r�֭EW�\�����H����4.}�����1��0|�L�mǛ���ѿT�h߆%�)&�%E�P����6Æ/\�(�C��s<<٥�@�2��Or�Oڼ�B��ϳS���<�&�\zd���8�$)a��9 �ss0���i���8�_����^UÇD"h�D �_>��i+*����Z�T%(�f��j�#J_؍�*�Ԣ���~7(�䁹�^&R���&w��p����'1�2�O/r?��L؂�$(c�j+�_��=�w���t��o�L����W��6��iU	�%���ޘ�
��n�Ƃ��X?�u����e�4�V��rO�k��Xc#�f)n��%1.���02cy�Z�%7���u7�\y�LC�h�N��ݷ��%�����R�ڔ���;&{���^�:�f�7Y��`�#�h[�t�fE�j1Y�Ah5�*J%S��u$���EU��lZ�3�G\���e��q�T����\�ETl����G��w:��Z�J;���އ�e�������y�8�Т�ģ=P�݌;̭�(|���DƍP:��o�<+��3�A9����K�EôN��h&|��s�L���u;��ڤ�󐬁�����2�4�aw��B��<�nF�J8������DYxo�=�T�9�Ҟ���	�f���)#O�
�x���V�ا-������^<i�>n�pY�T�y֙��/�A_|����� ��v��� �]+��̲�.�y���ނ�G�R�p����X�g�d؊�G$p���g�k}���c���LK��=��7��!�I�V%*S��nQ��uv���\�l$;�It��=9g�~ۤ�F>�j-|�2�o2Xf9��ydP7�v��'Ιo�͕�����d��b�3�
D�jQ-H|�v��=���/��}�QT��.ah�{ٞO
����;�ޝŽ�O�Ly���ʅ��W�I��
��מ�"+Ξ3��Ahg�Q_����mz�@���Bǀql6#�;�b��Y��CC���Ͷ�"W�8kbeZr<>��+
{F������7��`����OЋV�>��~8��d �J��ֻ����k�n��ш��z��ђ�0m�,�e����nϸ�/�;1~�|+t����e�2kH�����nŮ���iґ�Au
��5zፂ1�>%����\D��`y6�D:Kml�9,��C�#��I@�S)���sf��YD��{=]�u��w)��ɰ�2>�cL�m�c}f�j��&b��Q)8�(����v��$<�S����M��Ǯ���~q-o����Q"���ph/?�J��n�׀���x���CjD{r�����l�h"�DҖ����I�[�or��e��Z^'����n�w��56.�+����K�op���´A����4��
�SI�B��o��T#����lR�<��гl�I������4�2�u�g�"8�/>����B;��ևf:�� �F���>Y�F�W�,:U��ϵ�6k"�8�H4��+rFa�WFha�h��8��mE����t�u&���\�Ӗ�ok�h��R�C]��t��t�-Oھ(��eLh^[KS�i���ťO������&~ֺ�F��m!���S�t���W�� "&������a⟲z���5;{�8zT	�)�jO���b�;�·���"��� ��G(������3��/��H�\�1��fs[��2��`��!�h��Ƥc��r7�Ԡ��ts �*�o(2�Cl9�R��x� �?�vVD_�zd~i�Š�.��uqn�F����+l�~R΃'���]��B �z�J��P	�4��*�|q3L:p}(v���������5��/@���csU��(�ϝ��˂�������^Z41O��yJ=Psw¢A������'�\��s���'pHD �:5g�;[�l����K?��w�ZM2#�ꘗ�za���0�5��/q k[���_�S�ܨ��u \T�N���\ �;��$�B:���L8������ViK7�y����dI�8�d[>�b�.x���cH�q ��k�4h@�^��W^Ah}�Bۛ�R�½%R"�7H��J��W��Hpo�%Bl��S�wl;�,��-���E�.ߒ���D��j��
���Ŷ�:"v�x�N-tTPUc
���3eE=�H9�%,�CfO
������s�B`��I����>?V�@��>��eן��<�_�j[��c}�Ox��^���&�+aBƕꭺ~8!�M�B�شMlN�gX���[�n��cR' ����ܙ���TŹ���vᦛoE��'0�\�}����F�j�g��y	a��(vzf '����ñS���C/�Gy�<�����="�3�|� �f��tT1t:�i�;ff��E���U�It���ߪ?�C}gbe1��4��Lt"I$��*�)�~c��s~�Y3�8�/}+�2͉��D ��)�]��*�r�������e{63[j�Xu��� B}L�ke{%��X�>��$�I3�=�|�ݳ����)�3���(�6c�mŦ�v�&�k��oyʌ��~��ɲ�ec vK1/���2�p�� :;�
���Q�XN�����)h/�i
�E(*O ໯�F7�qv��'S�ࠇBKc�����WgEk��iŠ��m�4!	|a��E���?�N�4������XUCaj�����yY#����=7
pv�'c��q��C��r���E���}�:�	ٖ�3	h]~Fqo3ΰ�.�ܾ ���b ww-��}��.����[m�!�e
hQ��?a����a�ql�����E^X�Ik���R<m�V�����t���98l�,ˡ}�ѫB]fu��(Ԃ2�5q^/8v�ݳܡ�ՏY/�V��8Y�6vE8�����N�1B�km�*��� +e"â��&_2FB���Yc(��Z��:��4z�{�M���qb�@a�-̰F!���9����`w��?���oj/�be5�ϗo�F�����6�ǳ4,�eV�	��Y�?!ҥ9|L9;�P���Lr���T�K�'�k�:חd����㼆���X��Tv-��6����>�dYo��f��L�b0��P[����'�[�:��?����y�&�Z���|��ω��rjH�w�ټ��/7s��Q
#<��a��3�-}��@"���pZ��N�*�@w��)�&���v���(�h:�o����W���T3O�f��n�-��T��j��]��ĉd��*�r��S�� G����։�V���SA�~c��
�O���e�̅��m!Q���2e}2nk�F�2X[ͺ٩F�egHc�KfK��}�/��5|T���^���B<�X�`���������̔���d��Z�,m��c�43˞�ڴ6ؠw�J9 ʈ,��b)؞GT,�l�8)F^���1��[(��B!Z��!��ߑ����c�g��l���\G�����J�1)O�,8]�Z�.�M�趋�����'�n�Ww��~��kQ�д�,��_��t��߹�I�"�Yq��qx��J��{�CC~ u�X��Oc9�B���h�$p�������(��u|��A�c�%�>���%Y,��W��kY^�N�*��q�d���3�8K�i�܄�c����SQ7��eC#Ŗ����V��F �8m-"�#h�6bIN�
�<�0r	�a`��u��,.�B�L���\�g\���b�:��D'�H����m@N/R�/��8����aaɝw�'u�a4|Եj�l��@����eF.�݉ T�T�7+yĂ�;o,����m���P�G���5jA����k�+4RR���Mw1��1lLx�'��Mo}L������峁i[�����o�kF��I�t����,��s�/0�a�K�y���	�8b��`����W��)�	1�si�n�#�Ҹ��i�q����I�r��R�*����y�L��0%7ٻ8��6ka�8І�Ҧฺ�w8m?�"_���7I���[m*��V�� �pD�����V�R���m�c�p`��d�2������V�Y���(J�# E������{�����Y��`�q����e���/���dL��Ab�X��T��s��Y�w:�K���G�5QP��0��R�?����!*���sR<�Ckg�!��Oj��$�_��!�4�-�W��o�0:z�`��x��m59�w2פ��捒O�w�wAƯ�r�I��p�bU&��0�Xt�����3K�h1�ъ�[�f�[��K���`���p�)���j@�Ԁv�0�����h�UIf�`ԡ�pIh����Y^y=�[Xe��� �0!��<�#/��f�g2�W2��^�Y`�Ub[U�4�ܗ'Or��fέH�D��"��󴁜��;�
�������P7q)�7@W����\�27��}y��ْ��<�f��l�`���h�z��e	��-
@�_zS��ԋB�j"R�E��r��ӸGM2�[�k�v��Y潜c��L&$`���/�׀o����p\5#�7���9Y.�7�Hx��s[j�Q8.�`GK���C��vi�b�A�l�K�n�ÊiE�EU�]U�
�x���<�Eȷ��1��G�4��q�����C��w�N�Lҵ{��r4�~��b6�d���?��yV����]q�u���.$'���\顧Jzٸ�K��{S��z�h+SǋHd����Oxs��.O/o����L��ޠW��NWgb+�q�<��`��i��2�^�R�O�#u�y)��7�oƸ�ތfd+p��o�����:��Sϐگ�h�T�R��i��aT[�4�DL\lŮ����{n@J��Z�V���(XJ$;����?)�A������S�/ª��Rʢ�dnY�"�m�+��QJD���F̣�Sj,fGDv������7�17~��俶��U�l��s�0��%�(#9���iѷ�N�m�z,��nE/�#��A��<nm�&� ����M���բ�ulTZ�9�
Se�����/��L���oq������	8Bm=��ԮZV*�K/��U��a������	�7m��Kt��-���޴s������E[�-�b��iM����T+D.)4Tz���ը-��;Vh$Ȳ����z>�������;��S��}|1�����6��"��1�d��^k���!v(�.�z)��=�'��Q�E��]�C�OW����ZM�`"b�倗��`檹N��ɵ�r=��Y�*E�{X�[
j�FBY���0)�$�9.��̆��x�5e�j)�F�6;�� �1��gZN$� ����̙��蠋����2� �ǟ��;cI?� WP#\�B�9ݷ��_��U叇�XК��`n�APQS��	���O�;��/�;�iR�o����M�AAMN���"�o6����z�(ǛJ�hu���s��P�7�o�Ag��^u�K\�߾���<�����+ˁ9R�H�����Iz�%qQ�+x�[�=G�=�|�&喰*��qy�,�:���ʚ&h����9���W����5�D�j��$a���@<��ۆ��[�)x��y�i&�ɝ�.����OJT��8,�]t&��V�u��3�A�����::w=�*���+ڡ���J��<�+NK�Ȯ�:�Ј�{(��#ĵ?�T#��Zi��=�Y��=�����J�f����Ӑ��@��잕'�����hI������'i�R�^�]�\��i�0ilG�3�����%�z)�ƾXaP}��K3#�Z
C���..�e�d�<�g/ع��j<��7|?�B)��]�)�y�G�0�u�6�?.�/��m�⸍qS��l*��p*q�*ڂLdL?��le�H}q5G���;A���f$�w�R�	8�5k{�x����B]���wa� !������ӯ>�xW�k�7�޸�6���2�ơ������%H�a�+����\�s����>����-�p{��$uW�~��qR���v�9$v�<RW`��a
G�}I�4�;��^�ű���b�,~H��ca�s)��/%�����Av_|E������y��켫����,V䅈�)U˘	�4��2@��׽�Q�T��~MX�DܦF��'���<��M���u�J�r��#�Å�&W�D�Z�'͊�R�i��-[��B���̦
����G�\�Ye1��BF2��
��d?�m<s����E�ȬEj�m�<vh�V�'��rZ��N�jVꈡ����Egz�3�1�>�����"�A�<6�c<oJs�^�¼����R�j��F�\v��)�<�s�G��ZҘ�}��+�z�Z���:Q��A����I!����0�DO-Skn+�Jd�xK�<����[����BX3Ԟd�	��6c�0*֊{g�\a�WQ��<��l��m7��V� ��0�~Eݶ^DQ��MZ�Է<�ܧ�J��Lݕ�p�����!IRlL��&�b&����@�u��'�?����c�8��lP�'視��d�5:�*Mľxӻ2���'Z7h.%i&��B��������eà*�j]B�s��ݩsĸ��oƝ�QG��J�'%�֞����[l�+�}�"�x;�4����x�+`C�1c���V|)�G�48}��r���ﬥ����X�ff���a�D��i��f�����Chp�%I��2�ASҤ����/�1p�
�O٣Ô��Mxs��Ŋ�u�<��B���a�Eb,Y�r����cS,�t$�䇘�h*=o�U8d�Jf������.I"8����r����T�A�j�&� �σ@ ��M<��.o����E�'j���P�D�x�x�R�-���O�^��T-�[�](�D��	�r�@�qT�{��?�>�:����[����^q�ڒ���6�����*K>���͂Vm?P�w��jj�8	�;�nZ�� ��BxK���M\G�M�im9�Jt#2"�hr�"e)�������@+1���J��ԁ�
xHsx�@�ǣ�I`e�f��C[������o�_aA��VA���JF�i� [s�����o�Ħ��f�t��6�U�\��3��֡JQ��4n$��1�%�W��@ 'X'5��c2Kf��� q.�r�|�By��D^50�24ɱ��T@��:+�{A3(sͅWv�,�ꕎ)4��
����g�YmX�Տy ������7E1	1b�F��i'��	ޚ{,|h��7cM��w����2�R��A����ZT;�8��-��?��h
��NՋ�3� ��o"��5_�pз?�Ԝ��=K�����$�o�p8��7z�v��~F�(0���\�ԓ��bH����/��.�����[���@C�,>2lLQ� �
���Њ�������f]��u�Eů��>/�`��/�+���=�U��\�U��ng5���r�Ͳ��Sm��{���軔!��N �0�
��y[5�XqL�I���U�9�R�TK��ŇN��f]É���Ry,֭��Xa��Ɍ�3hؠ�dS_�Fΰ"��[���Q�=x�G��F~ ��.��Ĉe8H��(�M�\��EѪX�H��%��W����K<X�Iی��p�D��%�4'���Y(��?�&||�1�;Mx
�?!��f�e;	�rg��i����NFd�lA�AL��N361h������nUhu?�����g�0.�d�C�'�-��M���c,�5�������-`=��-u�G �U���D�3���u�+�{G����)Æw�c��#"2�������34C�:Mj�1���)�o���P	����o�.��K��Aho?��[�ko�1���[�A���
7��9 �H,P.^�T��w`ʔ�e�&}�N�� 䤕@���N��8�|��y  �Ma�8�}8Cn�l-�<�[F��9W9I����"R�Ы�v��\���|-�C����V�Zf<�p�`9t�a�o@�&<�4sD�TbJ������DO���S���p�S�Yʚ�=�KI�EOV/�l�7&A�L�j��D��X��z�Y�a���������cBh&���|@�
I�=�qwTF��]w�z��b�`�ٶuKF>���)�z@7�\S�)�罖��c�����SS����K�o��q�s�e�p�œ��k��~V����h��(.�i�K=�i�aj��Ce�@���*�Ƀ^�-J���Ш���ګ�G�9�ԫ������8/!�L�y	
V1�	�"o�Y��jg��F�l��I ��5��1�:QA�n�ķ��+�����M��Yp\��>{9��Z��q�l�)��t��a�]��-�jP�d��Ι.���̣]b�D��|�������)���>(4�C9��Ͻ�}gJ�	��]�XQJ��Y_1�7�m9���`���4��K?��>3M| (	y�B�;C1������bm`��>��!�M�)Ur�\�Jy����*q�j�"ѿh�g;~�=(��7CX-�SBA$�d��=�<�ս��)u�%��ٳ]j����A�93�P��c�6�ʰ?���Ɋ �6��}J�����ܝo�J��"�?=���◥�қw�6>�`_��7v�|�?�^QUb����Y��~8t�� �<C0N:���G����Gw���r��o�{_��;�K�������/����5��	2����h��+#�>0��bP���	�IC��-���1�m�v�����K#����3�����8 ���N��O��悝�"�0x_�o�;A�"��+��χ�^�m@�����Q.ȿ�"~Q�Ǉ,CKo��;��x\Ox��ऋ��I��Ńȅ����$rpy�;ͭ��ގ䂁3��e�l����I�iM��N�����A#��(��圹�ډ���g�u���?�v�5?,����D��,���{)�3��|v�T�	/A �������%i�[n�;�'��j `Y҄B�f�o)o'�����ۺ��K��tԪ�4��X2�k�VN=�e�e��r4z�:ԉe�xY���(����wJ��+�[$�(����{`q���a��\03�2d�ِ ��K�~qnR�R�~�~���8�X�t�عF��ҩ_� +����k��j�ku�����6�3�;񫡁�0$7M��K#'�Y�L|��4���r����at7����D���c�X��orNU������B�
.Ưm9���[�f=	����WX�][B�4�J�O���Y��^��m�'2 !Gzyw��=Հ\��.(@��~�[�q_��l���H���	{����e�����n����	�p����G��~�i��y�<i�_�صF�f�K�-��
Rb��uP�9v#��d���QP���TKp`-6Q����1h���*��� ��m�Q���;��]�Q���f	�&�i;n�kH���6q���`���&u<}�&��u#�}m��Br��(D�7ld��7^aFE�b���e!!(�h�_��*жb${kP4(�;�yנb�<|P}u���m�����K��Rig�M`�u����rY�� }���
�	�@<,��m������gc:��t�G�`�5����������п�'k6�A	
�Q<R�^;ad�2�9�UI/�_i���P���.���(b�Jz�zq���5X(���[�Zh��#T��?��0�k��Ӈ�DB ՍDVR�1Y�����ml����2���7z�Zt_h�MA�H~v�ʦ%|�){\��ϵ����Tuܧ����K��X���Re��0���6�����u	��"A���I=�찮�lu�|3*h�~�%�ޝ��c��+�ց_Q�ug�xi�5��>zm�Y��@*9�BZJ_�>�p��)~n���wD�K*����8C����c��;�p�k,��ʳ����kΑ����h���g��h�F�ɴ�|=�G�$�Y�3����g��3e�M1T%�UjVT���(����?k��EuX�i:����ℸF ���>�����yR��!\x�ƺ\��/���ˌ��bXq�"�IX�E���;�Yɚ���.�ZƝ�q��n�s��X�_MߚC͚���e�x۫pɍ���ֹ�����Orp̂��ε�a��,I`����^�o���0�a&GZ��ce���(��"�~V�z6���1���nf������s��hXt����?8*3� ��g�a�4w�Y@����6�*:�Q*'j�nEtΡ�kb��V`·�%�m��Rܞ�X����	�5W0M��Oc��牫�I��I�`o�)%r��8Ka��<���"��x��)�2�w�j��[ձm�k����^0�&�5��5�c����� ��0�ras�bb�f5C��86��o���ѩ-@ca��dj�^tA}M*�Ǐ�/F�W�P�U�Q��u��l(`l��;���w�K����l6�M{��$r�
��dH�g �����˞����K_����2���7�M`Rh変��Jo���~o��������^��{�N��v�!�39�A��mhjQokwFFֲz��3���&�o��a��W�}�5ﾲy�g^0IG�~7�Xa�[�)��7(d��M�н�-��~�|ه���CW�EK�s8���XGb頞�D��Z��\��V%�4#6b!��,���Zؒ_$��.7��ƭ=`p�D�hiE�����E��eW)\�]*
r�ˋ�ru��MS+�:���(���iKv}U\˶�vp��Q�Pd���܂�ok�I��D����1_�y���D&S�b�w#�X{����Cw�w�4A:@SX$J�&Q�vh,]ʮ�y�$qx�k��q�f�"���Z�k��̼��l��͊�xulA�0�����K�}��s�X�=��/�>Ao�k��[��2�D���K �iX�����'�{a`���T�l|����eVrӮ�ݼ`��W��<�q�|����'��}o��4��x>�z���%�1��Z�@x!䐾ͱ�}����Is�ҳv4��$��s�|��v�cq�aF�b�a���^i��'y�N݂ׅ�Q��Y.IG��Spc6���z�г��Is�P���g��5̬���������n��0|���u�_�=��~����,?WT�����zTD���	R��g�+�x�m��o0��T6��Ҿ�����놋K�F��7��=��S��ZA�8T�f{�Ģn�t�ǃ��k�w�fƱ��R��<s�n�"�1׹�f(w�ׯ�N�m����%�݃��ZNGnI`�� �+����bV��8�ʨ=���B@rK���$%�t215#Z�8Ƿ���M�bԽ2��q~2r��+���Nh�
Hh7j�k/4�*�j-�a&����y3c_e�}۩}G��̮�go�O��P@Z��&��A�
�+.�i�2�%Ż��e�Gq��
���Q��Ư�� xIڍ좢S�d�ZE	~���y���$��\kL�yGq~�x�F�ʨ��N$}� =+H����{�y8�C>�F[���Ɋ�"R��n"�֯
čΕ�c��o8���]���Dv�SM���>:=����K;	7���p�@|��[ɪLaoy?���\�k����w��$�FtW\z�3�&hH�Ȗrp��Ϗ��Kt�6:}x"(�C��9P�����!@� w,��S)B׭:�����k��R^�$S��?��g����F�=,�q ���%f��ɰ��d+k����cS���#��b����5���i788>TG?��A��v\Drh��p� �1N�������_�@��zl�q/� '?FJ�n8�G_q��:������v�h��Q�7G3�'qTV�Ā���}�=#��cd	P�'A�-.[Ӓɉ�P�i�HW�԰Z�� >N���"����G���)�CiI���_��d���E�8�ꢲw_��c�<s��R��:k�L�z0h:fQ��4.�,�B�O/6|�O'���|��0��@2C��U�1$���kr�Usq#-�F!@ 7{�����S�	M[Zڟa������
����!�;��m�8遛�h�*�F�,M�-���{M5�9GH`��ZMad��>�[�#���*
��΃�y�G��b���nt��^B��#Q����7��P�,8\�?�/�?���L����Src�\����T����&	�Ԙ�>N�ަ�_*6��~/,�LllFap����	�o	�h��v"�/�6���� 9������_�b���{�>��y�����U��_�t�PZ���{l�^p�T�NSe���ǩ{��G<�M]f2�$��rÈ�r�W-V�sk�c�s&��AN�E�F��.��S�� �a�$�l���z8	�@�%5�D7�z���פ�b�r@��"�ݢ4'�hf����W�B1�cM��#�%����`/.�rR~�Ԛ���g0���%�d��kV/p���<�{�CUSh�Q��@��B��ض����Խ�����$�q���R)h�=5O�m�M�;��x������/�� |z$l�{`����p'�ŗ�Z 'p���/׺NI6*���q2��d�ť�N��D�H��΍�`(��d�U�y�ʭ���힜���weO&��V���v
r�PE%�f�DG*�m���pG���gp�^Y:���-��?na<Z^��D�NK#���	�,�L$��*duL=y��ʰ�t�	�܏T�ƍ��>�y��V0d��q�8��%�iv�U?�罬I��N��V�ca�~���61���he>��F�/B"O�^̺g�dv�k��S��}�H���q@���W� ��R!��;�ԃ$Q���{�m�U��e��a[-uM#���d��p�27*4�g�iQJF'���)q��hC�T�^}�<�Ы�Z�W��<����˶�~������������t���~�.+�v�qN*���T�F��'G�t�3��q��髈U�����-��8����KG�:q����_�\9g�B)LK^�.����O��.��9�Yj�-]�������b�|��F6�Ώ�ta��M�i��a��u4���x�����zJu�m.����.]���W�ö���Ms���Ί�8t��r�~����|F�b�����_��p~OIE�Mz����ݧ�J\�s�^�
z�
שc=9�|��T�6+��n�%$��z������P��q�t|@2Vg���72��M���R������VO�!/6��}�lUn-0"�[�D���N�c�m�[�,̈́D�w�Â��u���e�栃]n���B��a��X��.�k2-�$}U4��� 7k�0�*΢��%�y_g�CA��?�l��x�4���b��� ��\�Je�v�r�Y{Z�2
��!n��p��tt&V�nӸ���&� g��P��d�z���\g�ZvtA�|��m ct�`v�  �A�P\���v(�׻��*`�@eZ�X����ظ�ʡ���h���5r��\k�����
9���]�G�{�%�L���vd��y�C���|��V��A����ȳ3G|3� r�"#}o�6�%�C�G�1��\����;�B��yX���	�-��0Y\�OVg���V��I͞�H�.���u��掠Y�{��p<�l�W�cz"%�8��f�	�񾰄j0�+gw���k�rD�}g��7%��1B��]�T�������	�#0��\�؎	�U:,%�?�n�Q��[J�c��b�+�@&; x�����|�B�I�,q`��S*l�v���L������ɤE�$^�[�1��e6u�(�b�v����	����3�2��2�Ȃ�*}<z�:kFM����Y��h��Z�)�,Pt�vF*�����
��8�(�f���T65Ռ���y�G�=C\��6�=���H�ۈI�N��<>�4_����!k��$(��=�5P盈��	i��۲��s�EQD·�ޕ�rvyIMZ~����Y�����cx�V�o��r��D�a��U�E�{L���e��[�o��4�f]v��f߱�2�o=8b��@��@�72�E��3�\ou��{��&��uA���#�a�t&�8O��	�$���s���%�v�I{�
3D��d�^��p�l�y�ߜN����X��z��4|l�(��$�Ty�4��h2�5�lE��֩!T�Y���a|u(���G�=�/R�5{a�̷2��!x��/d�뽗;l�I�������[<�C�@�.2��Tȣ�/$Ip�`��Q�h�q;�@2���t�P��B�0��߼G����8n�(8�Ǧx��^����#�޲bNΖ$h�FnY���������������ij�HuP��l-[V�=�O��15޷N/��섎���N���D��9��� ><& �O�S�-���/H��ۓÐ��2�ht9]X<�m���/703`�b�,��{��{�y�J��[�Bk��UZ�cE;HM��7�R�V�a脯Z�U���9e;��.Gd.7��M��0�Hno��Ǜg����H�<W�"�3�N��ܪ$������L��$��Sq��O��"O��L���WDq��|�y����c���`gn'��k��v�='�l��Y�ˌ�IK�%@��*��Ͻ�É�)�C�#���dÒ�U��I�vu:����5��~��9|�BC���ٜ{=$r�Gt	�j��I����]T6:�k�"����ۙ���.�I��+!!�o♬|�����s[^�
R!!�Q��c���W�M�kim����F<�$b�������[�����(?�����ң�c�����Q���st�cK�� ��`E��A��$x��B�̘#}�l?|�2lZ�����pP����h�7�W#AZ�Lv����&>Lk��r��p��rH�=Lv�#�H�F��=k#��U�_�o>w�(z��{(vy3
��-�˷�|Z U���(=�a�O��1O�IЦ}7��!�U����x�S�L�/v,����KY����(]+ȣg#A�OUU"=��>+^ �����W�gJn��I^ �4 x�%�RR��)��An�oԇ�H��A�=�"���i����2��߰I����@�.���ߒ'[�W�:����UlG�b��Y�&Q{�_Z�|��!�K[�>�Xєb��S���×n��m�m�����;�=�Jqg�ĺ�a�/E�R��:����)�
��,ppۋ.k�Z �V`,Q� ���2��?"�i�nOg�*M���ל�t9���,r�*�*��\�a�}���%�Q�.�(MIp��4hbA�� >],5i2����������n�i�9��6��F��^g����T�\�}N�^��VrVr�F��m���]����1R�It����d{�L��I�cɺ;#���~�1�g���w_��}>�����Qz�6S�Ē:��Mq�}�V�V>�+0N��[�i��N/Rt��Vy�AN�A�k�%��E}�$����6�P���bۙLr��m�`5h~�}b!���;h��!�tRx��G)r�Ӟ
��r��G�
�!�
�<Y٢��) *� '�.�� �tԳ��A�S�;?�����b����	M�&U=��Z�J���L������98`L��ڟW�T 6>�Vͼ7%�<�]I"�:l�VO}Ŀ��(��|���0���Yg��mA}�2l�#nP݆<J��{i�/�!L߲���U%'*5(����ܢ���6}s�6'n杜!c��)��� �N��d�h��@�$�9��)��T4�=���;��Hc��~��.���va���I�=̔��jB�(���1���/�sz� ��_ɸ����]K� �.BF}��K���k��
�0x���r̈́���@.���J��	�?Ӕ�t�����uR�4c$T�P�?v`�^B����E� ��Z�/DJ�Ī��'��jC4Ƌ�K�ez2��ӝ����Ew��X(0݉�UA�,TTQ-=u�z�Cr�����i�!�|��=�\�b�!|u	��I��ۊ�N�2B�R�G�v�\���{�;v�^�ޗ3`��f�#�(�M1�f5��Mǭ�I�~Ar����PLS�.oʦ�$�HG�BQ|�\Mq���g|�GPي�����1��@o�w�6�ҫ�� ���}�(����-�Q�����G##�]͠Ş�_�P��e��8�,���h(
�&1�lf)��h~5i[iA��0I��`���X{~�>.#���͉���X_������B	(Ⱥ�캾��ܒ��ɴ~Z����hz���q�Ȝf�S�F��k�,<��#�]2&�W9pZ��ʡ�x�VwS d�G�5��I���{���1�2�+2^8J7�;���A�[v#қ{���wY4��p����g@�Xf���V�<r?�ҴЖ���B(B�֦X�-�h�o_5R;\�&���l6�	�Th�h�g�ko�.hsό�2(���sA
�̴m��=��7�qLD�!�f*%%�C�@ �,G�$4��6SI�ngޖ^1j�-������m�E�i��~�5g�v9�����2��8"�cE���A����Dck���6�#-~�.�����d*���Bߌ���w��y�C���;���V�&���ԛ���N�um�@��r�� ���fc�2�X����,fS|&�`%�L��(�װ(%�c_h��/�it�E�y0��7���g�L%��yr���=��Q7��=�
Y?��2:����_Z[�h�(Ş�.ip�	Of7�]���������������-�~�0W�a�� JQ�6��;Ի[x�u��ų�=
@�����n�݊J*������{gL�r*��xG�H#r�!dʎQ����d��9S
>Y$yxaJ~X�,��s����q߯��j���>9̇��C���5�\E�p6����~8��@= �.��AT�0e!ȫc�ԑ4� M�Π��&A�q�/wk(�5��ڿ0�]��6'��P���U��囿�(��f�>�A�W~�H���ar����ae�� ���`�EYAO��X���@j^�	�ϛ(ydwzҁ )$aɃ��|c�D搆��}���v-�tM���ʘ~�n��3�y����ߩ���������
���%�h��R�{_c;�q��ԭ��A�V��g)�	U��$*����"	�4Q�y�Z��V?��̟�� %��و�r�?t��w�h��k��[���{N�|��S?Y���8�QD�~gBT�6�@���	�����츟6���_��.)M
��y}�&��g/��G�^S�R���$�r�7�M�'xg����N9WofbX��/��?N+p�*gG���5_�7B�
�j����\�ޔ����\�]��������c-ެ�3KG����:D�Я���߯����}��F�4c醠�)s��?�ZVm��bR֊�uZ���ЅG��v]�������;��q�i8(��S�Z�%�לn^���*������(eu��.��ixJ����t�Bֽ�#5	+�%��#�%/�*1,�Rfݺ I$�҅����$��б�J�Lc�D�Gr��O\�/�I��y�L���8A���R5�"Q�)�$�鈜j�\p=���e���i9)RY��L*@s�(UX��&�;��h+��1Rt����O��|n����9��T�b���f��O��?�)��e>V|�(�fZ������ٌ�7X��NU�Œ�6��~�y��ַ�z��G����^F;Ntv��5��Q95��������hv��{A����e��w�f���k�v���`�]�A_�{Jf���	���]K�Qp�l6�8�V1�c����h\�V�VA�>�Q� �ْ��&{oN�s�T8�Ϫ���H�V�e<���+0ӏ6z�uh{5�����R%b����|J�P ��C����B�T��[��Y
ޙ������;Vv��sj��p]�b,P$V����q��s/V���G����?�3K�L��$.&�X���g���n(] E^[���,U�H����!2*lF�ɛ�g���x�$�\�D���`0#�`��F- ݑ4�����ܾ�K�G䳊��0����R�\��d�x�Cf�.IC]f4}��)ƌ�UK= �ΐ4��@Nh�)D[(�Tt�U���u���F�`Pf�]����D��A�.$�h$_F�������1h�仨��G=�Y2~6vSSJ?��}����S����uũD܁����v�*M��[B���'�Z�m���B�o?��A�u���uJ]� B�3�I=��3���ĳ��]�2W�./;0�d�-����h��n�G�8����vS���k��&"پ����M͉����t|u�3��y��HJ�zPØ�HЂ�iQ+�Q2��1�HK膉��~w��1�᩟|.�P�֧��'J9�߬�9�44�&g��Ы�W�H� ծ��4�a�(�MLa~���[$o
�5c3��w��RT!r5�p�3Y\ʂ� Gʺ>����<����+��@�@QN��@��3���9Bw���7��}�}/"C�YX�Yꛮb� �4v����3�����Jc�07	,@ �-�Ӄ:�/��9b ��U��
uL�%�v�k�q�5a��L�nV
L���K�k�K&*����h�l��i��K�UXM�0)�q7�`��0*�rU���-ޑ���xΜ_x2�f6��m�=��}��NB�+WX��87k��l���ѺF�T$]������ݗ���6EД�>����
�^y�	�#�{��U�ă���3\� ���r}�m�t,偧�����t3���(~%�-���/є* |Q�W
��R��7�F���jb�4���r�؎!�҈�� �@*��s��O�+&����7c�潸a�<F����F��<�]E�l}m�{H܂)3ܱ+��R\/F.	\����
b�.1}���5�P��ֺ����i�y��R��<�D��m��"�Z�R������v���"�[�1`@��o��P4����]R�����jQ)�2�|�0-cDiӿ��c��6	_��Kgn�Ua��4��2hJ�%�x�mw�}��r���U)���4���S5T������0��T��������A�v ���E6Џ1?7�lx�؊g'.��Ar���y��Γ��k܅R�>������]�,����TT1�9�"�e�SA?��ظ�#TyVߎ�����{y��u�$�n��%Y�im�4,_\��+�76\�o�� 	���	���]�-��x[�� p]��
c$�Ν1��C z
����mE�/0���5`�X/u�qr[����g	ײ wQ�0�OWO��.'X$�ɘz���{ �
tH�����$)�ٙn��Ӕj�Z�ΙZ��{P�?�eG�e��!�Ya&]LC믞Wf%��q����u<	�2�Me	�Q��pwU�kw@ =� ��ԛNN`�[bv�0>�8�b����l��(�,|r�oP\�r�����3+�Kz����Y�ǯ�?�w����U��X__91e����c�g��ɽ$�Y������;*{�S�J���t�� ������K���D/mMHBV%&y�Tj���4NvD�J^��է������_��=�7��5y���S˲b`Q��N�[�� ������� �i{>���q>�ڱ/y�H�[H�W<e����,l��p�a�� �1%� ܸ<I{�U� ,�����(g�}N=�;�8iM���&O�pPO,y�8������T3Kn�c۶�QL_
K�C۞�4�����P��D�H;N&��䱭�-�a�բx!#��/Fh���'|AZF�-2�*j1E6�I��qWS�Q_Bs7�.��	A��q��br��o�m�g�.�s�8���0��1�({��\=�+0cO�s�*�^�y|ջ�T��>�L:N�����(�(F�\���[��+��q4	�<x�~x��9>����N�q����$�����%HO$�>�z����uE��D����T�E�H4�ܹ��ޝ�n"J`*��rزʺ�Ded�&I<���|�GV�S�j�'���T���N�����0x��+��ި���-�p!� �2�r�>\�U���Y��e��;�/�O���HQU�uV�<����ƕHN��pͽ�UA��T�^�x�U�u�>��[��q�Ԫ���x�B��d�b��(8zH�XiY�8{�H�w��,�PM���e'�[`�Ƙ$�H[�\�Fn�K��b�<�W�� WU�>�V�Ͳu�2[����b;�Z5u�6	��X�����uhC���X��Z��Nv ���M�s�*��j+��ܒ*\���g�3[��6��A��]u�C�z�v����ϰ�&b�عV�M=x��20�*S��`��e�����b�@{��2��f2x�c��6x��?Y_d~̔����k�.��n����<�z�����=�U���c	ӟ��I���	jE��7Q�R{�%l�������HH�˚��D��]�6{B���v�����6�gc�Ӄ�
��n��s+yH"���C�m���]p�lgJQ޼2{��*^X�, �	��x�6��_��)��^ނ��$0,�/?U��j�_�G�'f�J"���Zͤ�$�H~˅b��E�b��_\��۱0>� R���9g�6����Yi��)���Q�Nu4[.8L���;�WT����}A���40��((�pŴ�B_!Q��/��T����jIq*�`��껫��K|��O��~�L���*i����^f�R��d���b��k�
V@>ߓkɣh��u	-5���j���sA��O��5��HY�U����;N���#�S�K҅ �W�����v�ܛ�F�/�G���a=��\vt��>�z$�7˔�x��d|�}�b9=K�z��Q�a�-�SM�P[<N]R\2:̋RW6�F2`MР?����/�A]��ߕ�S��e���I~V�,K���cȩ�_�I���J����j��Q�+:^��&m�����Ce�I�D[>���n�����sc�>Z1���z�Ƭ�d�Ɛk���7s�>��Jh�^���b:E?6�r���#p�k�+�Bc��м������D��\Cj�[�x-�����G�%:��Ʒ����@����/���?WsИ:�Q�e��Z,h�K2�v0'��?&��HڔSi�ż�u��[�r���}t�/��`a��:�R��^<Q��	�i��L|��+ �DS�����̶���� ��Ŗ�.�_�]���E@�!Ϻ�4W&�<�s#v�}�P��z�}�12�	�����¥={�g�x�*�J�j|/��	-��#�	!�}���"΂(m����yJ@WEE"�y�#�U�YaE�a�!'�������o�!�!��-��4Ge�ӣR �?Z+MK�h��� l�����W�JՌ��/�����Xb@r�d&�v�YDf���Ә�ؐq��`�j�Y�*�w\��4���G� vS��qr�}9���l"�6�)I8�Ӝ�:>��P��z�ö�j�G�@=�!��_b��㷻���m.%Dl#I�	|���pM+�d��@�2��_�g����S,{c�/������\�����4���Ɛ�UX�����`�lf��r���v�L�jCP�X� ��!������AM "E�G��S�ݎhn�@L!�KP���gͻ���"�e�ޢ2��ZD��F^U�r����g��F�8n 캕�) ����W5q�V�&Uꃢ��������k��Ě<O�~�6t��-�$����������)���_^��0��w�`�6����{��_�*�H3;��>�ެ=V�hVS5v�I�5\F�Չ��99/�&b��b&���`W;WpQK�^��ľ�n��ӽyp1��_	w�E�%ݞ����,j�Z�N8q�Ȫǀ+������E��Ĉf�J6">m߀�O��Χ�E��v�_�P��`�SJ�&�JGS}�<ZW��ΰ��UDuZ ��E�%�_��,��#�B�ݫ�;������T�U��DЬ����˶��;����d�1GB�o|]�ڈ����|�5Q�w����|"MKo>]�P�ɶW��J�c�Ya\�x�-��[.�I����m,s��r"�fѻze�\~=�!���hfX�#[,��sg�r��	�U\��R����އA��{
4v�{k�D�/g�ݙ$X�H~A�֧�%bP�Y�Չ��;�U��z|��q��^���v\�l@�Ix`��.L=��A�ֳu�=���L��:/q7���H*���q���֑�oXj��B�G��4#�����S�����j�,������p |��pu�XK���������]�	vg#J��&j_¼a6��R�}����}o�T>������~S�	���9�<c���5~m�}F�>���A��f[0��\���N�3%�����ªP3�~���Sl9�����5��C˝'Js(�&�I��P�����+�/�r�e��Լ<\�1 6�D�9ك�f�{%c�GY��T�z�c#��xp�}Ѡ\ � [Y�^������;E�M%�1��ă�z���$,�[I�Ǵ��5/M΅/�\� ���W��3���Wm.8��H�Z"/#�mZ�]h��3�g�Ba>�rD,��\�B��.vt�n�|��^��F�f��[
��i(���xu�����tTm�|#��F-uɛ��(�C3zK��o���kun!յv1��x��Oj4�0�١=>��<Ѕ�Mc_Ns�]��G� �=0���n�i��}���=6��z�Ȗ�*�1��3,�X�i�� �pj����nt��z�ZCW܏�Lbw�6l<6�Z� �r�� ����Y��z�X���7�	؀�υ?7kƂ)��l��޲�0Jx��i��H-�ȋ�|F�B�{��Lzt8����{�9 �#e�G7\������>�]�P�A+�-l��ƬX�>6���{�$�jP`JG��к5�:���b%�����ݬij"���p����T�������~��aHW�ʂ��Q;���/�M���h�m5<�:����=�Mgi�m�O�*U�_�XWQX"��.�|�~�]���Ў���&�4rY�y e���!֏h�ݿ�Ab;��RY����aAKx��S��֢#H'����K{;��yy�V"�)�`8���W@��Pm7�����=A�N�?1v��}+~�% ��������b���Ʒ�¥�i|ŭ"�k��M��ۋ��R�/����DxQ�+�}�����A�����44���{����A��8'�G��kU�&��)�{�7<�ػ�Y1*z%�dL����9;���&s�wz���z�����oc���f�1�~��lh X��q@`�ϵ���`��4�[
�/M9d��1jW���R�[R��'���y(��߆�����UǶ� �'�.�'UA/"��o�p���!?>��G*��	?�?��3�Ba3�)����󫴯�0}��v4���:V���}+�[�2���{��w�
2��enǺQ��E+�G(YU�0�>�@ml����@]��!��h�_+���AZ,2��N�_��2&�U�d��F�פ��b��f�}��|��9�2�b�?�\�w[�Ė��UM�h��jd^�=���ok�����t�����Y(�s�%��"lgv7�}Cפ#2v�_����	��n}Uh$I_t�M��=����[V.FX�	p��_��kp�W�pU�@r���N���҆��QK�~1(��O-������f[߂�gӖ��[�OO������+n��s~���
x�:|�Y���i�j�Ǆ:�2n��<HmP��G�s�O�u���{�Rv���E�~����S�p![Oş
~Sq��y̕��`�x>�d��V:Y��̠c�^��gG�, �HkK����� �������	{/"�{F���W��x�%G�v�S���S���5
5��W�ܻ@@���h���C��ܹ�h3��v����;u�n�
���n.�C��/HQ8A��(�:7�ګ�c ��M0;c�q��=�X�w�����r�DsTo��6���p*�0ULݴ����݇��qE#��L��"���f�Vx˿�����!����-"�Gb�7��"��Gx�
	��b(k�kRl�6Y�1Hd}�Ç�{uL��a�e���	��}� �&�~�m=�K��ޟ�a�}8�k���8����U%/�k%��Ք�~�_�W�]��&(�a��Kya��ކG<Wıf�wC
��M��kZi�#x�)�BƹJ^�<�$���|7�`�$��v[�^~v;m��f�S]�4�����xRL�J;�� _�A!�G�LC
�`�:�� ���8I���]"�v�/:t~�
�8l]����5G@>G�g��.0��2�ygD�8�qc_��8DI})�h.�֥1N����J�E�!
�]��T���U�O�j�*}D�*�6�-L��Ȃy�
I�o}����d�ϪD6�{!��̣X���R'�{)J��&�B�$� L�Qk�d0X�󊫰o�ל������Z!&/�����7014FN9��'7K'(VժM�����@q@�9��<t���~����j:�E�
np0���F�{F9i1������S�������/�dR��o�J��1W�ռ�¹h�9���;8�����Z,��(b�T�����5�)6CI�y�`Z�g�g��*	�s
=<��Ĝ�Uɣ�i�S`lB��IZ3-�∉�,q�$�>(�ģ����9|�榉�c�I~���Ha8�e��~����\a���]uX�D�l#��]w��ג���E�ۭ��7�3���ٍ�b_m�7qY�]���|�T	���za�9[��(��ٳ��f�:pfHtuP;�N���mZ!s�@Ǌl;AK>'U䒝����c΀���;�P�x�<r�~,����U�Q��T��H�y7�;�ۂ�ĝW��WU��	b��w=8*/�V.R�¬|��j����W	��t�b����\�_R��E���\4�3�ٮ�-�,j =j���Êl�	���8�Jc�q}Wx�����,R�@�%����O��A<�E$���j)�$��X�7
4C�!�~�5����q�f�ZNg#p��4�D%��V� 8-�@��8�i�g�2?%��4�Xy�\�$l�Q����a�/>�|ƭ�������uQA.�U\�� ��Pux=�����ɟW	>���#�������ƀe{�H���E�f�I��$m�y�$b�]��ע��Y@��d�t̞��R���[��V�ェ����*�p��Ho�"#C2!Z�%l����1@1�SQ�I����؊fP�����b>K�?�b�"�~@���#�H.������{w�����ְ@���	�5��^JÅU�὚��\Π#h}�5���<3�#���f��3iU#�M�'�@=������fL�$EFv��t���Z��x�w�aU�Ĕ���w�#*�.+=�y<p��t�5��9�E3}]X��a���T��D kq��{�]���<.��u
�HS6��T��v.�=;}��<���=P�i�� �Ƀ��xtj&��o�4}��h���G�Y&#�����d�����ƓUu$���6;kh����h�O����Kx/�D�'{'�WߧJ��&�V�	��$������@��.�:�[��`��	A��==��¿X�{�<�9���X�԰5g\��EqI��3�~64Rz+�:������<
T?T������ʾ�>	��VE):	��ގ�4sRs��X�m}�A:�����ہ��c���Yy�﹵�!
ʩ�|:	���Z �U�K/b���?��c��:-\�`B|^������M�H��v*��9�l7�������<WڞJ�+2�T+�Ղ� ���a�xx}N� ���`��g���9�钄v���2`]�I�h��Ϡ�����Q>�ߴ��v�*��_.K~�gS;�|�e�U�as(s׹�Tݵ�`.�[N�?s���-��x͜�<�T�����ߩ\�}T�w�d��EX՛&58y�r�e#��Pf쓑��&�k�	^S�	�:+ז�F?�Q��zYE����t�: w���O"�[����<�R�`&�܆�g�K\�蕣u3"�/.DA�����Lq�b;�i'�sN!�&Y�=�EY�`eO�-�#��*r���A�h^#�&�	ңXޛ�*�	�X��Ӎ��D�M?��|�n2P�ԍ��Px�\G2�BܴG��A��1����L� �(���Uk�<Qn�5���������Hy��n4��pg,���`���½��xB���Z��ΝC��=���b@��8��/\��"P���Jk����y�F~hY�=�2&�v+����d�����nM�Bm:\ �J����Z���P�|y���;qۯg$F��t>����̓3�Ԏ��9ī�-�����ـ��#����j#�EQ��,��V�:�-篐���ݣyEо�,+�/L����Y�e)�Ã����vae���2�n�.v���oX��~-\��8��OcS��ֳ��;��� M���/O�(9j.j���ن��s�����]q���r�?��2=�v`=�E[�N���N�02�X��>�� ����c���N�T��2H��RDəII���)y�+ z��^��JJ��]���Rsqi�v�i�(ݕ����ޒ4} �`IU�f2n��W��6�xA�~��w��7S��E���Q��f��A~k�ׇ�ON��� ���x\�����O'?C���P.ܦ�ڜ��1T<��"��Q;3#���8��U��̴n�@=�	���SN�2�dP�	��l%��,~Y.I0���zN:����+K�U�k&�?���̤�Ey>W%�H�z�F��&y!�0U�s:�Ѷ�2���������I���Uz�T'�%��>5�;3۬,�U�}wol��. b�p�¦GD9z%�ӶAuDK�����V�0��A��..�#���e�8+S��X����N�88��9Jyc�J<d�g���o�����G/I&�E/5���]���%!���zw���QT�AmG��J<{�����j�=��V>�R@F)G<��X��)�:)�����ڂ�z (L�1�����ryY��1 U�J���xpW ����+΂����k���<���Jv��c��p5C���NU���ԩʹI��+�lA���3x]��_�\�>7J�h|큿���Av�.�C�	%l����5���e��㉆�^�b�ش�d)F�ᙧc8����v���ü�س�h~���BK�������=�]�y�I��t��Y��^^�M�,w�6�m��ƮH>?�zL���y��>I�.[�?$�z?�#�Ȉq�6ؕ�-�ea�g��}K U̫�܇ �h/6%.,�Si���uZ�=?�)���XH����@���]�����S��6�[]q&i��QO��SJY͈��n��?)�|8k�U~��e�s��E}�4�����2.[C���}����zR�H1��r\?��j�����d�&�'
E����=�U����_�g�F!m�43Qx��x��Y�?$�3��T{
�{f{�A�Bm]��i�'�5#�y�EØҜ���Ԅ.t�*����,��xɛ�=���r���ؘ̢֝��6�������di� b!�d�\�jz 0����b0ǴS��Ns�Re��rOa��@���Ķ`d�Vna�:y%��s��5����Kv���dz1�Y�
b�-�D��(�vQ�:���h�V{�@J���3�@|�ld ���b���y[p�=@�Lƨ/h��q�$U�F��sV$z"���y�#fhكO�a�}ѣd��-�>�Ъq���[N�1}iY�]��X��3�J������O��n�IeQ���*�x�<?.uV�܌P�ƩeX��@�z��П��*�B'���[_I9���̢��t�0k�{5�����J69��;%�q�[�uyD��!����L�h,��j=�ew<4.����Y��y��+�}3������3�'xʻ�L���{M�����ޥ��m�ϑ�{vp�]e�ީ3�2�����˖�;�O�G��F�s7I�nnl���6
z�*{�%���Ea�+U���0;R�ż�-����2�+��x#�4�!�
���U��H�d�`��,��?���]sO���/�xGI����I�n$�Y�*�^p����t.ը51c�C�8��R^�G$� l��3*`�u�>C �L @t��걋h2�Q��R�d�/>'M`�	�q��x&I�)z��q�/�\�D��Y��c��sn����N�ss�nZXIM'?�JES$�޾�t{�h��9�+*��Psl۽E��<P��A����:���6�e�K����T|�o�������HP�:Б�"`Fֺ�8�v[�&74��ݓa��d� ���[�����S+����Nϸ�X R�|��� ��S�g=�3�wd(
��m ՗�p�%P"\9���&7rſ���Y�l�)�B�f>�����w�u�����+D4�<���o���6��N��������#��|+�nV
��Ҍ�ɬ|ut��#�80)�p��(�8t��!����t?���X�x�k��
��?#��*�HܸEtf����榟� ����}ϥ��`�gr�~�����(@�ל X��xo�҈/��[ƺ�a���P���hy7�e���֖b��%%��NX�ki�Y'���\�D�%�6�y=�n�g{�T|���ֳ����A(
�ô��vAd��?�o�4�&��H]����8���p�3Ξ�H[5c:���ֵt����s��k��� �����m�]=
�8�3�E�8?
*��a/��b����0��Qf1�.��	��[,'�x��1z�=�l5nh �U6e �_��(��nE|��P���/��X�C�mR:�
��􎲂]���/|[�Nw��[��Vv���F��5W': [/���᪵+>�[�%7.�O�=W�yAV����w���jn�ޭs;��}[W3�}?��hX1�Jy��a��3,���ť�6e�c����ђ*�ja�{��^�tؖ�L��U@�0�"��Oeie�����H�]I����l<w���UN ��C}!�J�ˏm����2���h\�L:V���ŲP�(M��Nß�c�~q6u�&��H㝺��1>�ϓB{Ӗ��Z�(���S�X�=KT Q�>��H#������ �C������s�<��ʧ�R�*8~.���&�\|E[�V�0�Z���`{ S��)l�G^�`�h�}1�̤�Kqm ��kyy�,!z����6 ��Yj��U�F�[����)�W7j6ݸ���_�\��2k�5��}2Q_�����~�I����@��ߎL��XkT��{�˲&%�8-�tw	GT}��j������%�Od���(���津�����[�=�����@,,3�=�]��<�Xf��(��g�p�ޫ��;�c!�i�w�qn�ֈs�����;����J�cI��o̝��_�y!�*T"q��E�6A���-y�ϋ+���92W�m$�� ve�!��A����+'{��Ч�#�^����b�+��B0u�w�[Ad<��~8�%vY_v6ծ���z����H(���7g�	�kb\u����L��  ƺ9���'�*�@G�|��H�HT�8HRE��˛�ʁ+@P&rȱ󟿐�a�8sͬ�	���T�<���+t/.���U�q��l��l҄�b�O�i��c[���,�d��m�6��U:!�Yi�W/��~b0c��ixW�6�6�$SEޥ?�1zA�s0N,&t�.��﹝,��y���'��RL��ǚ}�,%�	�&;�������O𡈉X���L��i)׼X���gU��t��1�Пa��q��1*C�u�~�l��CwǿqΎ���a��J댻&��B�O�$�]���0�R�"����:�H�\o%��WM}>3a���Q��'4�t(u�HB�C�ti˪��U��5�)0^$R�%X�He�R�2%��x��aH`c]R����S]9��
#)BvQ�O��K��,�9%���Y��a�����V#Z"��T����-��,l��k�w�h���Ѷ��d�)��z&��5���Ǒ�('h�x�Dȭ����d[��Ҝ�?M��l�]���h~��� �L47����J?bR���+�3-ŽMơ2@� {w�7%Z>C@��¥�����ʻ ��9U����/yPB�zĵ4��e a��X��w{�����ȒY�YK���z��s�޻c��5ݹ3*'����鍀���jju����=c}Q�*k�i]��K�̄S���"V�	��c�3�.Oc\V;�=B0�&�F�_����E�,(��?9Ι�T�c4b�`�(q�X�.H_�b��@!Pդ�[@�N|��w��l5x+�8+7�8����6��u���>c�&�4o��\N�:zn�J���W!�w�ltϨ���5V�1r,���+
�Sb�H�nC*���2n1������N�|8~�������^oK�c&��!,�����~]�Oo��vs��8fm� �/a&���3D��$D�����}�n>@hќ��<|����>���s,��q�UĶl/[d����Mink���� ���Z�����t�х{OE��f�$�W{���������:6�V����-
�[�|M�א,���hB��s��'܊���j��h�?�S5J&DF.�O�o	�J<4������]������d��Xa�Ϛ��H����~��\^��.G~ã��;abÌ��%��4q�5���M��E	 -x�Y'm��s{(�]9�C��N�<���;��]ϏY�c����fė����I=���n����7��3�.��A�sA�����9��nm�M?t�[�}�.p��S�9��ZՒ���~�V�w��8��H;n0*�^��,U�(:rg�������@a�=8|�}_����N|�4���2F��Ki7�2H���������^i�O^;rQȳG<v3�-��(ڛ_�hSZ��ۃ���w��Y��*x�J����G3B_1Fb a.3���h%RFGrNœ�^�S~��LX�Ň-}z��in�1gDZ��lRuv�Jm4�� ���E��x/�Px��R��0�{S�e�󜐂~I���	�jf�Q�,��5Չ�i��.ga)v2�zM�p�o�_���++P��2)��+�,3Rs��~� C��}>Q���x� #&w��1���4RE��!���ܦ�A_T��8n�SҁX�x��d5����1���D�V���Wv��"2�~�K������3�o/`��}�T~t�ͣ�$,b^w�JH�v6�[G�3LR�v�O<�E	�ǌ�O�O�W��EV{e�/MR�*�f�Ac�}���=2�n{�9(9z�(
����
�ZT{ʎO�ʾJ,>��
'�N0����9����a9B� 7"�5���Tk�������b���85�mkN}�YcY�E��❝�*�cd1�x��i�{�/v͛2�����R~Ð���/9�6�P���G�Y�\d|�N����K2��ʙ`Q����2�l�N�ȟ	MU����{� ��'��t��ԇ�Yt��G�I��Q �]]%�	5)Ϫ0,J��KQ�?U��_�Nwr����~�l��3r����y��(m��1�|~���粑sr�B���V�X-�:б���lU�nE<(��HIP�+P�H�^�y�t�gw| �W�n�y�f���ܽ\ٲ�!����k��Q�U���4�7��(� �J��,#�^H� �l�&��u���nD�Lŕ�n�՘2�o>%�C�~����ܝ�w����6E!s�7�v6�G굕��׬ҳ��a&Om<��$��m� l�;Bv�o̸-pp�O��� ����_8�B��W{&�u��k$�� �K`�N�0����m�!G`���G0�ᵌ��p��z �]ә^��K��*��X�b{�����kф�GVڒ��=���e*��%�Y���K�8F�W�&QMЦ%�b�o��Iـ��ބ}�ba�V��&P�g��>w�72UIzh�L|��RW�=�F�믱����i��v��B���yr��g��� Ϲ3w�x�����0B׳��,���ġ8�{��v�+)��c՜,<���R��%G�o��K�o���[���$��}�"\c�94հz�;�i��vk͡�|��Ζ?�5�&��Z�;�:	s$A��K+��n�#��
��B�a�h�$N(2>�;EO��T��hE@q�a�t}!��a��_T,�d+����o�}�Ԍ��w�mz�y��!7	� �F���Ƃ�b�v$�am�7�� ���ы����������B�F��._#��.8������1��k�ˤ�����<�t�t����4�X�,�~h�:�g�n�6��6�c���BV&���풖��k�kL�K8�x��M�����T��K�"�Y9�jS~3�����_t�P0r�T�qLS�ؤ �aT*G��9��-f%��h�Y�����ϵ\$.� Da�m�#�#{!l3D���� �\5�-iu��f%�PT�lڈ[��X!����R��k��bv���8$�d�m���7��{f����5l�b�B_����8��F�փB��],�� :�v���f�vL�c�M��ш��/��I��Ӛ�ֿp�J�;�P�i��پŲ5�"�>�����+�]�3#���!���1���'o�NU�/YqR��.��?����-����Y��L�N��9��zXe,wP�{�?u�j�l��\"���|"�7��"�S�F���	�G�۷J+i�9t�QAQxe6&bd	:v�3�a�������=��&0�}}��T
!����f��|�b����[�]B���6�)�y	[mV=Gai؃T��I���wM�[��6Ze��獠�(��#��1GT�i���5�*����kŁ��u�U�Dë�L2����6���[��p��L�R��s������X�T�3��!�.7xˋ�4�
���QI�?ϱ�p�8���f]F��t����.>��~O�&���e��ݰ�xm� i�3]�Oi8�L���*-���R��S'��sct��b?�AG�:@ڿVE�l���(D�������e�X�ƭ�?<��K{�X��7��u�{:a!_8qa��C*$� ���6R��ԢI�r_`?A�O�ц$ϥ:xS̬�Fs	�\���&��5��+;gF���b�ԩ�Z�8Nx�S�w2��7b�:K/1`��v�]���Ʃ��o�{_�c\ !k����ӣM�<H��Cĉ:O��K�3������}s:���M;����C�,bBM�դ���`7����j�*��p�h�κjRj"�K��U�x��T��]Ujm�[N�&�je��@�>�~���5*y��U�,#�c�9��ii:����vX��r��7r�M���x_��~�7�d�"��w��G1Q,�tgpєRs�H ���2/�8U�6d�N$ʂ��YN2D-PR8��f�	��_Jp��=JD��u)<BS��*S����ȼw�7�?�䊤��,S|�:kr�\��$�<���P73��AuO�V��M��ހ�&}��V�,��vBYR�|�M�j9�y��*c��7�.9�+HU����o���|h�_T,��Q�:#O�td ����D����Ɇ'Ȳ��l��J>��0�+��.�x9"C�[>��֪hr-x����߬���2��uo������}�%�O*�<|fVs�Lx��&�^���Z�:Y���Ò��7m�w)ia��V���I�̘x?qR�!
v� w��,��0��b[��b�I��ŧ5�U�1m8��v��Q,Qud��M��H 8o�� +��'� :ru|h�0zGy:9�8R��4,�'?}(�h���T����l���8Z����#-�j��*k�`W�+�^]�W��Ѐ΄PT�%����a�p����-��!�"�"(�Xv����^��G}�냆7�n���>*�q��;17],����f���L���OŋFf��t�j"���MܟX� }���~K�4p8<
����JW<,	��:QT	r}��Aݹ$��n!i����˂��wQ-Ԍ���/S	k�F�
v�WwR�E����'�K,:m���I���\�&�;
�>&��Rl�4�#�?�Y$�r�Xa�nݨ�tҡ���[�'&JSC�$S[W�oC-|�\��~�3��,��o'�8�B��}�א/�RN7��+�W4��=[`}�h�? �5h�3K���/u������P"�O�����������!�hΌ�K��9T�}B;<�/C�5����ɹ/���3���7�
��U�� Q�Zp[�m�7��-5i�K2�Z�l_iP����Ӈ=�Up>����BBMEٷ��z��Z�>/p�9��:<��6��SI�|P���B��Ln�	YnUD	��S�����b��i�^0��(��3i!�$��WLd�w�4�+��!����F�%���HPS��]���N���eYS��l�S^z<�T�Et�Zyp���?j�K �����A�P�l=�jE�O��$�Ĥ8+��2������S8?
�o�����ݑ��b�y��#jD�5���_�~��<��^�L�64�Q�.�r�����I>����G�x�UR���ko�pc��]����#����ש�vo�%��$�$I}o��x�丮<�����k�`ڹ��%GEv#)f��6\�(��6t��"�V���] O�#,��<�Fs-#U�'`��KX�)>Ņ�PR^-'��S���`�Fh��T>~��F��<ƿ�喝�nK,�=O�ly�B�2e�ņ8����l�(B��L{,o#����wV��֣Ss��C(m����o.:��� Y�e�����I�-�XCH�r�T{�}+T-�}5����C�R����c��B��,��l��X�V�D4!�����M3�w��3Nb(��VF9�EQB#�OZϷT�cq��@��|߶�I��T��� ����lֆM�(���/�N�	����}ev�S�=|�},���~<��h�y��K��S��t�e�22�K�y�U��~�����W���.�@���l%%�E�h��v�8������ž�-�������(�%�FhA�M�[4���pGc��QX�F?��uu=��%<�ڨ�����p|�����*q8��1R�lQLj��R p�b�;�iW�dԎq?!�(��q�q�_0A�+I��_���f^�e�s�0���m��;�N7�4Z�����o�O0a7�Ҩ¬`�����W��-���Y��o�13��p�Qʡ�_�8�i�����@fŎI�ZQV�4��u����#]1(��G��1�Z����,� #��ڥ`@Ĝ6�����tK�</k=~��wc�~�ת��ü,Ҿ�B�E�>��!6���@:Q���%�E�>& e�����7M��f�������Pҍ%�,*N������[ٌ7����/�{P��eQĥ�<����g`V��A�^i�rn�yo'�����v����.��΅��!i��S�	�Ra���
����}��9��p�1�u��� H�U�\��V�M�SFXw��蛡v)�u/p�]I��O��FY����i�r٪t���,teU�ѷ��8!TT���w�|����NIX;�T��E�\Ih�l}ǠOd�ˈ!�JՄ��a��AM�C��KZ�U�Z�	��ƫ�M� ��.���{�0���P�D_"y[C]�$\�6!�b�4�p�c���5w
􁔄l�����A� ��q��p<Q�Qꞕ;�`\j�9K����Z�&W{\����&�/X�-Eď�\�˙U!�EWwd����V��|�!�-�4�8���>��~�=�;��&i�zB~��;i���������4�!,i�i��t��E
�����]7��Y����4��^?q����gn1�(s�޲�("¬
6����4=��V�����ŇC y�¸��A�t/}@z�� \�у�ϼ"�A�q��/Z�}�����K�~2��e{`���Fڽgh�����Ug��Ɛ⽩a�,�.�:�%N>Ry}Tǐ
9��Kx&[��E�@mFp&��	���ǢB�����r��ٔ�/QO�>�gO�A�5�;L^�C�.�u��/׊�+��������ͤ4JZ�����'��e(
�1�Y�j����GǏj�N0���u��M�\��1�ϙ����"|����F�Ha�J�]?g�헦�
��C�����#(�Ʋ���^�ngG�)V��K1ُ�i��:&�q*�fj�,_�@��~��ꩤn v�1;�~B8!v��xe��pY�,��Ƞ�F-��u���w?��l��R}iUWK�0O��ɂ�	>��J9��\6�\���ރ�Roꆲt��.�4=���C|��"q˯��(���㮫Os�����~[���b��L	�$ml���\=�ha�eMX&�U��*�х�^"�Ƨ���D������;���Q���,�![�/�=le��{�_�D9�>aP���o���|.���u
xIQ�:�$͢4vo��c�2�u6���L&���0��z(��̾CdR*����@e��=���Y�1x?8t�c�S�
�X�����#�[���D�)�ʌ���)�%M0M����8�����q�����|�'�i �� ����GB��=�*A�$�Hq=����2�Ƭ�$x�)�4�~�|;�,ۄO�W�a��#�׬�����Fe}LZ�|��ً	�@UO�LCмA�N^}d�Y�{^GrC�!�l;a���H��N��T �}X�_Tv>t�����p)���I��k��{��lc��;O�w$"��=�ӄ��<���s+�s�����	��
����#%�ʃ� ��w�:�v����A�l��+o���+	�MQ�Q�T������O)��#.þ�Q�� �y��̈́۠�0�z�"rG��2[O�G�`�kH{�A�������2gl)�����e�`g�8�T�Mvщ�9'T��	�[�꜊���#1H�;��T�=&7���,(ı�Ə�;4W��:�P������K}jV�#����É��Ż}o�V��3դ����>�D�]0?�#L]u��X�ػ�=*{�)������=���͒�}��Q���f��R�>�{^�=��q<�\������H��jˮ������\O:JX�塚�!��R�p"s�P	}�1Q%,d�-h5�@ ��%4��ݦa�~��dI�[�m������2������}A�1�nET�"�M�l�&G��T^�#�輍J���nS ૾# �C�4����|y���j�︂�&��<ah�nq��J>��`p�\�ܻ�cR�dR�7�ȸ
9�	Nk�UIw`n*\����(�V��Op�Mpݼ8����*���A���{��N[�� \��E��	Z�yղ���O�ħ�.��MR�aޣ��kf��E�~�)�|��X�(U)���A?e�a��W�m_��YxE4�E��6s����'�:��*U�4L�\g}��ʖ�̪�+��\0�"���k���.?�e�A�g˕��-�o����&�áVY���No��׽��fʥ�q�xl�`y�=P�q��ϙl���zK8&e)�խL�Q�PFq �8���c�x�+ � e:\��6o�m|{�G�:b��aAdO �/�c�sUgVZ�������1�c�Ts�1�Gl.�
�����翛a_���z��ǲ��%�K�C����);�Y�x�JI?�'&S9��L!�Q׊�� �P�|�����ű���i��u�G��va���z����u `'7����m|�vZGLWq�ӆ$���m�QW�O�A<詽��bt@�wOL����7W�;O6���'�=[�p�D�ͬoe_�b����y&0n&�K`�io�e���-�1�낦�y����|,@�+�|.�j���7�d3�����;��4@��������C��_\�pp�m�Hl�g�K@Q�
��blI�)}��*�A I�.�qgY6΀.n�06r0�wġ&?Vq�͠7�cf�K�GMoZ��:2irr���g�K�t=��g��D�'e�;�|`U궿i�@,���sW��ꦞ�Y�P���x% d����j��.����,D��VFth��/	��evx����Ӫ�7���]O ��as~D��W���a�G��q���e�\��7:�㘚)�z�1=!p�-θ%_gY�4q����� b����:���o�-�!¶�<��������#�R��? dWݵ�DG����=�۲r2����M\U�-�
�����E.8.9,)$��`;Z�z�3�\Tn�G�Y,�'!��w�4^SQW�����@Rֶ3��@h8t�`�r����|˟�§e`[op\OH����,@����U��s��m�x߬�7��1�#�vRB��An;��`���-�7�J���z�8l�-�r�������]�:0����Q�tk��3_k�j�^gVV�%�L��f_T���#�����Q�f@��sܿ����J���G�4?$F�4E{�'=q�����y��F�b���q���~�`�Z�����f-q�q�*�E[��\n�@x����OV'��e*��z�_)?��w���E�w�EAZ��jb>����\� !Eờ���Hɰ9�����z6o�F	8=�{�T*/ͭ��2��I,���|���l��i�e��F��j2׊�栏��M��&��/��?�n�5N0�T<B^zȴ�++4'�p�����i9�1g��Iwg|�8a�{�I�,4ٕ�EE����O�F2^L{�R��eH:�Ɂ�;?3N����m�EN��Ԭ�����h����z�l��U!����eYF�%��t��❹I�4�w���#�Z$[��р9�2L���
���k���g����+`��m���%�R.*W����� �S=)�i�-�K=�}۲�}LM���s��U@�h��)�� u�"R��}�A1o>HW�ۈ��Zc��iZ�ꁆa
���'u6J�זjs�bD�rT�C�]�]�8ۘ�@���5���ـA��5�n�	�z�]5�Y�]�*b,�J��,ʿ�O���`��������DC>K�4b��+Gl�(P��ڕ8c�'󃵭`>��I(^���p�]C��[��PB�Dg�(A{����Z�)�#DѤ�7������H�X�� �|Gٜ2R��O��60۩QuwE���I(?ct�a�f	�L6�R�1z1*2Py��!Tǂ���#�w���͊��>SzNvT^�MB�4V��<Z�D5�"����ܧ�Ůܥ�����y�!��&�,���<����X�[����B��]�=n��P�c�z"&��
!9�b���wU�O����WJ�Y��Y����b�]l7b��=Dr�y,\x���R⤠q��'<�"΃�M�@�P�hؾ�2U8��faWXpP����-6�m�� K���B�eq�Ė�!�k���!��d�\�0���%��q'I�WC� T��_W2Y2>} ��b6�`�N��}6���&շ���뱩aa����l
��k�0��n�nTb~ҡ�c�]�;� vu)Ct5'"��U������53�zL�5�ok�G+���/k�v��|O�_ads��$��$ &�"V*��#C�}�k
����փ�Or�^�:�>��Q��uXW�'�E�:0SԪ�kp ��p=�;���lLc���%YM?��ez��K�_x�C���p��_��ÐӃo@ɦd���P�n�tws��gM?ơ�*>�_�>H�$�K�l�>�}���#��A�B�hP���'��7L��$��O�QSxb��� ����u�tRh-Bs�k��5�����e�� Y��1��׮���D���6���0����Q��]���;m�h�d,
�U6=S��(5��n�����=XV��HTٮ�.(R�g������y����L>$��k� ��0܁��VN_����'`7'	Yc_|��g�4�.=�X����<�������9fB	�̏���s��r��Rd�t��S�I�w���-�Ƨ����/�	#����-xM&��p��7��h{|�2���:YA3ҺD�_�8�
��J�In5���L�� =+�_px�ހ�4�_��Jfp*H(�g���wä�3\��Z��^ǜ�ۺ��[/��Qf$�}�!�����`�F 5�&���ZU^����{s� �_G�ĺ����fM���:g��OAd*#1��Q��!,��;��K"@
�+�N���弩w�[��:��^b����Wb!�ʊM���&�a��Q���� ��B����P:����E>�aB�`��i/�[~*zm:5p��{��aQ�+��3��1q�Z{
�$Ų�5RL�U�U$Ny���oέ�� �'��#�N�4E������+&B(ҋ��fð����X�<򖟶�p��]^��w�7F�11N�"��c�qJhf�I�r����@��a���n�۷{�� ��yMƭ1`����&y�za�P, 
��g=	��NS��.����p���5� -"���s���3�&���!���x��r}�,֢cj{zg-Pq���H��?l����p�7�A9��R~�ߗTO��9U��h,�k�m��Ħ^"Nw� �j�7D�n/.��'��o�C8t00��]#��W�Td��c���1#%���u�eې��vrܯ
��e����9�7s�i�R`f#���T��E�5�Þq��M�5M=��`���)�5%�y��ib�i��aڈ���T��E	;�J{�r��u�isk(�U��2<o�g�����e�D�w��i�V���3W'�;(e-+גOQ�j�25�AUN�O�����ѱ&�\RTs�]���rI�E��Q�/"�M����Ѐ�P���ļġ�֮���@,����s�
�p�n��.=(���T��>��	f�go�a�cq��FKzRG�Hf�/V�2�l@.�hJ@L������ǋ+�f���ȌϪ~�, ՗��L�S��}>��ڻ2�*�T
Q��V�J��%��h_�9��މ[���a�������"j�I�G�_<�7��@��4xސK�}����3�2��2+�v�HU�	9�e2nA�"��ߣ�LTT�-�kN�1�����X�!u-do&�����]�q�^W�ޅ�����v�Gco+�j��f��<�룜�?�E�8b�$�1���!�R/8���z��[�]�A�c��T��dV�����l0f�����&��fV�qn(�}̗'�ҞV�r+���\�Ǚ&U^��w�ϙq��;#e�Ii�����t�
�P�n�G�ŁP]>���� M�j�5d�I�Ve�T�Ě�D����`�jܙTl���I;|���Q[Q��_���X��r r�������|�Po��V��kzX����C����9kX�zt��1��$?�O]�ԁV�� �'��ze�e�g�����������Ɩ3�wY�����������.�i���K�s>�J{U�-��H4�v;�G
�F{Oeg&�jVes/[�@`����;�M�u�s�N9������Z;�,y:��LM�2�3��4�'	AwC�D�H�����G���<�P_�B탵.g�o�.��TK3���e�_�ou�JH���ݤ�c$��]ҩI�_�Ȩߚ8]�R^B��/�쥋���r��[�fψ����݌�,���nf���i=ռ��L���qcTD������oI�|}�S���OӬE�6�l�Mb�a�y��+'9&�rPU�'4����,���R���c�%��Lʵ9�1�"�nÍ!�mX(��#����;4_zv�+�|s:hz!d�vl�U*%�*J�3��L.MJ7�ӮǄ�=����[�!H<-��\������E�0�;���мs��Y��&�J8'�@�:pS>���ǰ��J�A�V`A�.�Z�Q*��u�0��&5�zc�@CPWu�v�V�DK�o�[^
x���6��py�����l��pHɅNtl( T�-���$�p�fB�����u���L��L׆�W= �Z�,�J���O��p�P#��	dopoPdt��Fʶ@Z�^xv�����ԐY�:�TM7gv��Bb��������/�w�����B~�i�i�8��h��N�k������<����!���3h�J���9�Q�>�!_�{ {�e��J���y�g�|K�͔���Q�-_K�� ^�d`����r �Bߋ�<A`�`SK�O��i�q�*Kp����=�m��-1��W����"�n@���J�Bpm��b��|_§��!Y�k�uwgiw���H
�*�nd	�q����H�A���L�k���D4p�sRW�hj�.�[5g��#-6X>��� �}��.}��%��)�mNBp�rI��h76Dl�S��_G��{�!�	웩4���@*���'���e̔����We8�V��Ȗ��l�XF=}LF�7�� 4�QGfV�@�8��˽]�KKy���<�Ő�/"�Ԍ��2���
�����H5�$P��qO���V���R1I�\%�3]���\���[s!�k>�Nh�����8���y�f�*�:�shwA;��
?��f��:�@Yga{,��tC�5���k��1{���W�{����"�a"�o�#�Y$Y�3pE3l��}*"< �.#*��C<����ڰ��S��X�l5�QLI�����9�Q�01� #�3I�5��b~X���[с��ׂ��X+4��Ғ����̃�dҊ�F��Dѻ����D�"!�yЪGy-���`|����� �ĢY�J<�q��k}� ە�˫���@�%����	f'J򔮮GqW�8�a3l�B��Jc��x6��^ƅAp2ߋl<X|!�\�72��,���@
�x�`�VV�)*S�<���6��zfu�_#��R�&������+��|b�t���-}�Xso�8=M�	�w�j�z��
>5�\P4zf����Y��G�8�KD9�.�|PBR>?�H Z	V��M�gq�Wf��v7���	�+���������W{��z%5Fg?��p�G�;�u�Mr{�4��П����Ԣ�J����(��oP�T���́�1�Rف��i_�)N.]ߑ�Y>U�Z��0�]� �DZ��ԣ��>nZ�Z�u��N"x>�&�Y�:�s�����%J�`.L^����57ɟV����-.�F��_y�(r\�9�*����6��z��Ν��G�/k*v���LM��2T���H0+{�K�����W���L$Ӯ�ӣ�鎩������؈S	�)=}7��<�R0����t���$T5N����J�
K_�l1*�r�2�l�%z��N��Ӑۣ��������p���Y��`)�M���2X\w`��;�F�^�k�z˛A��K�k:��R��+�^�#�3���D�P���y^�;kOgֽ�Ϗ1�}�~Yz3nm��馏��l"x��L��TE��2m؋��\'�T�>aԇ�,6�j)����Ӗ��������l��139�R���|�g1B$��9P��{K_�W�@��l�7kC4G�	�Sz�hbڷok�g���d�Rif�O�������[w�哳r�n�)�\����N^63~�-
c���]�BwNױ�^{$�-�dB�6���f|����� R�F:���yjd�W՝� *-��(��'/P>�Ct�[/O���&"��W�n�`F�O�b|+폃Gk��0�2f�^�0Vp﷩�!���i��"[ZZD���&��c+��7#xV�x6�\���H�J�aែ�g��:�9��~���?�=�T�2�W�l���C8�,�*�fy���\�|�����j���RI�OԮ:D��� [����s ��F�TfJ�T��X��<��M�>.�Q��F9}�e���J�Q~+f]���͊qA0���%z�r/��c�u�շ+����NI'�rH�I��\��?���^���f��W��E5��b�j��p �$S�j�<%#P�t���M�3 �$d�J������	�=�����K��������%��ؖ��seL���� uE��L�"V� �g�&4�0�6�?�3�gzoA����l�9������8p&!`�'���J��X����|�K�v���|X�5��kh*�<8^]�]sy��xC�	d��H���Ő>Q�ȃ%]��J��[ 7RO1f�m<��Fm�J:�%�����\M�j*�f�0]5�i����m��Ｌ!N��T�-).�S��˒���q:F.�&���ȋ�>)�|F�q�'x� -��t��HQ?9a`UGvt�4�IQ�E�C�{%�{��n��'�V�pc���(tZ������_:v0����(��>�?��cȬH}Y������� fx4*6�w���{�]�%��l�p;��`N��v�`A�wj�u�)fdZ��n0yҼ�����;J��L*	��br���1m|�keY-,s鎵P����0
��킅����n������6M��q�Dݮ{�}��&�e��9��l�z�Vϒ{��VP�@,�"�s�t1�H�eSq�nH�~���a|̾t0侀T=n�<d��98!��]"ԕ�dK�b��eO���P�YexL< ����+-C�bh�b�d����!;u�F�u�8��'�ig@��]�w�.[ ���%�+{}T?���Ō�R�f�GX�Pt9�H�!�)̊o oS���83h�L-��g�	P�/l9�bGP*��m[,�a�F�f��S`�΢M�j� ǜ��*����?�~��?��BXo��١N:�-)��o�����z= V:������7$���;��1�@�Vu.ų;.Bk՝q��\�v��
��!�Y)œ�Q�lA���q�~"3��ŧs.��$I�D%�]���5���-�XW�|���3��Ή������5��8�_X��/U���O8�n���#["�4RM��g�I���6��[�Y���А5q��N�V���2�Y�+��4y��d�����=+Y� [߰�Ǧ���"���_�?@����V��5� O��H�l�S��T������N��/-���o�`�iF���1Y�L~X�_ �N�T*��W�^	C����n됟��C�嫄���8�}M �$N��෷#A�@�pIm+��e|�����`"��(
���X/��νm������|+�Ү4����1�c#;�A�$�ϥ��� !��e_s�q�~0?�rH�<y�%�[�U������vL!t�n� ��6�B�۞��a�,�|�ן6U2�0h�=)�;���.��O��l��_�Q��,������|��vI��F�� ��F��/�4M��	{-`��ERo
����d%��.̭�:�g#�.�?F	�q���Y�6/��'6�`D���%�0���V'��b~8�r�gI]�zk7��o��9oe���/�"���L��\E��@��B��9j�� p�����=�y����PP�����/6�����*�.��0��|��ʰ��u��8��˝��pk��*�A%Zg�L�r�٪π��O9�C�V�ݔLB��%4v0��m�/m���KH�s��	�R�=CI;�E|ω�����UǊ��PM�yx�.> d��G���ͩP��L���?�e��s�k�s��Y��	�� ��\u�Z��i<�?�Ж(�q�8+/�Ts��]&��m��rNSz�J�B���:л����NJ�zZ"���.tM ����N�h�U�@"7�V�3�;z��}yf��6��v�����828�*%RX�φɄpkZ0�N��v5����'��xV�b�)ȓT͠d����ِN ��G1Ù�W��}�������ѽ�T�?U�?�|�[+ҁ�
�	���11T�-��+QE�~�>^@ߩaT(C���1�ćn� �T^��^��e���¥%w�y�����
���׍|^s�i���F��=M�]�oM�O���!W�����ͬqwA��1��y
�Fbx4�j����E>W<�&o/��\p���e�Es)g���>4���;_X�@�*�}�qST��Ǜ-`4�v#P���/���+Q�T)	�4G^���f�S	tNP�nml�T }�[��r�-��0���k�̖�Wg�}�Vф]z5d:��4M�wy�|5����c���hA�ϣ p�#�� ;%���������{L�@*y�	�K��D�JV������`EZ��������5,�����YȠ�<&�#�m�<�+b�
V�ݻ+��i�mzQ�J���@��wf�s���x\P��?�Y7�7��v*e�T`��Td��z��5=�v\�ه��dϣ�+,�}πI%� ��Q�&��3�c��j�ҁu
X�U���FA� i���I\��{�6���!����)�m;�2P�您3��ZS��H�31V�|o�PfoW�6��E�g�;X�p���RX)��U^�g:?`���J�Y�c(���Z�v�nW���Ӭ�ל����y�A�WD>���S��#:GR�"6E ~!��L����l�.�����w�6��=�&'Lw�g��m�c�G���h��~�[J����fG�n�,{rԳR�h;����Ŭ&1�T&PEP2UE9��Yy�Gz{��o"�(nq����?ɐ��ݤ;�h�������`	�}R�u�AK-���,/N5UvVPR�}%��g�_0rDU-c��@M}o��}j�>3{�M|\�J��zl��7�s�ax,�+�7N����/��<3&ؐ<G�}�H���p�e��ȿ�I��g[����(� �{FV�;٨5Ť���z3��W>�ū�kwC��t�ĩ��tӬ3k�R��nK���I%�r�����\c%M�å�yE��旕*cGӎ?������ζ��Y�s�:/#��y��|�)$%�%�l����������$���?���k$�7�_9S�-Z���Qy� o7Ylo���U��I�%������ ��w��
p�0<v|�|�M������9u+�;6X|ncpR,����(�$�1H��Ҧݬ����ΠnxØ����y�0*��N9�3�B��4�HH���g���P.���p;�	ۣ�=�7�y󚏳��\����(���3���z���&6$\�6���͒�\�������S ��|�'�uz4����]{��H�J�!�qX�j/�?�5&e�j?>J���7j1ID�,�#��wp�C�n!-c#�T�{��\�BN���	-���y�I�'�J��X�I2���^���/-�
��g��SEk+SŐ �>tD)I�E��Ek !�ĵ$�`��~�f�GxF��\@b�9g%ni�Q$�klB2�KO�'"`�5���Su/=w)�����-��dlSQ�C����֤m'�<���5�fا�k���Ƌ��	[4r���b�O��l�<�޾����R���/�Vx�Z�W�K����� ��!���/ G��>{M�S;�Z\J�v���2�i���:�쾈K�����k�.Z��rB)Kж��;��e<{X&�����O~MHc��Q]�r�l�px�3٧�U��F�l�!٨�&��%���/ K���̹���:�z��@l����sTVf�AF��TG��}�d��/�[6p:�ia���4"}y���H-��=��Y���>K@��1�Wn����9�"��� "͊/'����8I�;@���d��2�h�L瑏�q��^24���(^�P��ʴ��8S��3]z"��X����+g�A�ga����"��4��U�y�?�����,:�0F�+��`e[ĄJ;�$��S�M;��:2fH�DC��-�ߴ��À!�w��k�l�r����*!���K��0�X�b4P`�$$9a�«��\���J����.n�����5t���ޜ_i�H�l+۸�f�;yy����agyk��D%�#R��JU!��e|z9זX�j�cC~��eKT_�̗H��	���@�@%�7o�xKO�������Fl;�֑��a=3����5j{0X~*�f,�('0��;��f��g����O�p�{¸�'�ӳw�#���T�).����TJPO%�2
As�wǿzĕHc1'=���grs��0P�+=d��Q����j�w5eZ�n3����I��@���qŢ��x�'*$��m��4�V����=��!�E����B��6cr8�m��Q%1�v�����O�ј���"�'�:r�w�a��%T�S�#�}� bx����n�2��sO��6�D�������\x���1�ZKHm�rF)�9g	���ߐ��!��.�*�D1[�H����� &=���� �)�y`N&'�+����N�x���]��Ѵ�.c��wP�����s�f��)R\� #�D�ݴ������4�*b�Z	Ę�����K���H�z�+|�J��~�1��Z9���������g�9)⪡S��IU6
�SQov (x�Ƒ�6{JA�SE���>�g��c2�gL��sE��*���L�$�"+Ѿ,�����]�d�)��dG�
�ʣ`�X�1*��B��q]|�;���"!�9���`��G����gʻ�k̦Y1�~[O#g���.%�[&2O�A���j�Ѩ�!3�C�Ij����+~��P㣎�B�K�{��l���c��=�Q��	��/5Dƭ��)��R
5��Փ��o膈7��8ɇ��B�M�Et�����X^��U�~�����	�Z�o�@tc%�|�l�A�';s�Z��	�g�TԸZ�a$F�cR������u@��]�vy��B���M�~!�Pc�_�����.��������:��3P\��r����P=&��qO�H�dd�|��T�vƼ>-���3����A�M��A.*_�9�#_eRB\n�LK�x��C]T|�,���e��.4s��{�?Sl�ӊ �t�z�܍ϔ��!:82lF���=���1|x���B]�q�d���q�(�7C�b��� �)��ci�&U��fTRW�M'ŋ�ϭ�.\����t-���Z�0���T��m�ڊ�u����4[If�V6%�_��U4놉h�\�+����!�7��A�,��L8)�1�[qk���V;]���sA�����{����{�ʴ¦���]�[ȬA-B��w�D?CV�����uYu��~�	���k��m,�4@��#�Q�����]+�8���<�h�%�	1� Z^��(�Ǻ�􊻬��Ӳ���(�:��������D�%d�����~��� R/!N�IVf�1yT���gS�9��q'�Ⱥ�9�g'���oS�dd�}�Z�{$��xV8���)O�"�ۃ�|���랱觤 ��N���|y
�"w	A��uo���֤x8�ϡ�o_�P����� �X|�b�&B�Mh�����L�b9x�U��T;�,�_N�%�wx����{�A�����t7��`�W��I:	e0�:���� �2���H~��`��į1���jQq-����p����9�p�Τ�a��e\+�k������v7"4@DBv}}��bD
���e��������J���VV�%��ɵ�c4#�S��G�
%�;za�{Q+�^Z�2�&�7(b]�~��<ܲ�������������zo<1���#���Y|ְ������)�3�V���ZY��m_ׂi]���ь��;���i���hksF�I�c$��|������F��K�E�^!Fc�� ��-r���uj�j?̝��h�tU��)np|���gaG�cMm4�rX:X!)˚h�U���Zչ�/wY&,����wI-"BT�A�F͛=����r��ĦcYT��a�h}�։&��m�1t��e���ڽA�YE�qg��p�,���Q�'iZ��M����pZ�S�Sƾ��+l��]W��_vD����e��F@�IV`�󽤵]���7�oI��?���ԣ-��R�*��Y"�a�)�Ru�iB�C�(�����q�7%�e�W�.=��}{� �jv�ĉi�n��3b�����C��Dgrޅ=���E�1�����qa��c�;����,[X���� #�\�>�*��m�:����\�2���j]�[�5%�G���Z4�^��u]-E���(r���]}"�6���hG�����̒&�uvBy�2e�rU[���W -,��)Ƹ���n��f��k������ut�� ��v�l�R���>�Ѹ+�E��V}71�[F��T<h"�*7�Y��{$����EY��:g Yė��k�(�~�j� c�֥�5\��U��JJ����:r��s��2��=�)6R��0�0q��:|���|:���#�\�Y���S�CT�|�U*�� ŕ)^����zTq���V�2G2T�=��~EC@��rm�/��M�����ǧ�A���Б�ȯ�4B���*�P˻V�J�g�<��`���K��ė7��χG�<���1aMf�XN���p�^4�ŧ%�Bt��ࢩ̂��a��ݮ��(��F$jW�;�� ��	�^�#<���gT���w\�9���Q�eᓫ���k��u�bw��ܯ�=\�6���eD:�K��g�l��1TvE%fZ�,u-��ӈ����R#XP�g3��@l21>�K��l��+�j�7�b����a���x����+�u�C���DݐM�C$҈ؿ+�a�a楶Avơ�jl���Hu��OAj)1˖� ����X�0Ȧ���2������K�!y�:�% �mR�}u�xI�Q3'$�c�i/^·ÃJ�Y0A�P������Ua��,{E�*��X�Z�! q��>3�E��Ф~�i-=��
*>�R�1w��0�Z�����#Bks~�� �]wv�_�?�H�� 
��|Q�!�F|CV������Vpc���(��+�|0T��D�*g�Nn��@S�����L�U
�{nNh������NP��B)\4xщ�vsi
¨��% ��<P�T���V9�N�c!P�{�#��6�]-����L�Sf��S�m�ϒ��f��k�-gK���^e�6�s���":���匨��JIe�η��\����0L��J1��(�O#������m�O¢{@F㬦�;��<�Ș�E6�M�����c�g��jh�Y�S�'V}l������th_)��/���Zz���03�ݫg�y�u��@��%Ff#���.����5�jFƲ1満�ifAX/�-�ϗ��<����xUïx�}�(��"�k�O������ng�=��#�]d�%$���͕P�H\��X�-;s���X�b�uC�j��&_XdB�|bu��A�Y��64�`	�cr\�<n3�|�ϡ�|���"h�[�R]e�t肠����S�pz�����P�Q�[�Uc˪8�e��1th
�%=�вq� ���:o��74suX���Ⱦ����|�uˁ��p�:�G�y�����5��a�:�3��(J`�kRd�۞�%�ju�&
��!�@�P�}&G�W ��W���ṅ�[�P��oU�I�������F�b�~�U�}��<��n��_W�$��:]�m�Ӣ��#NB��6�o>"[ס$yr�?�m�6�?E`t���pkP���'����g�R�n(̬B�g\DA�%������)�ռH���t�tDt�L��x2R��Q����3(*��ݧ����2�������Bk���,D��*���@`�mo�������W�r��~s�za����������$A���~w�҅��Bݙ��<;eCi��h�2"&�>�+��/Mo��F�J��sRWstiv SiPn�tMJb��"��h��m顋�RuL��N:0�qn&��t���DcS/�e�x�m���l�T����{(�
�xYD�ϛ�@��'����3F�p�O]߇���D��bS��"����
L�0��"�d��;;9���o9/:�p��(2�/��J��L�C�#���#0�qC���f���G�>;���a��Ty��X��'F��
�11�,�L�J��}�8��*��3�eҘ����\���U��s�g����B/v�n����*6��F��Z�Y�b{TD1r�/���׳�g�t�k�����4gR�G��4@�q��USqC
5ۭ�Q�,��Y��iV��CS;���L0�?F �!P^[X�u*��s0`���N@��`Ʒ����������a��%��[I)��$x�Ed�[a����p8L-��ѢQ"�#��C$��xAH�f��=mT-�j��/�L����3p3r����u2��6��'yM�,)-����&h��_r�&HJ�o��(ܿ��E#lѹ�y�Y���Q;��x-1<�%荍�g���V����2�h��U*$�ۛ0I6�]p�@��Yj��|S>�P�~�Gsf�@j�]b$���"���,x������%��vi����'r]UW9�.� %AKa�s�ZA>h��}q�s�5�s�~l`,_�,����)�׫U��EcN9��qI{��W���w?��jr�����˿Y�$���Z�b�y��Ӥc�S�aN��q�_��# VC�)Hz���8�����ͬK���BSJ�k�K5~.'_@³�`(�چ�Ӱ%R�Z�,:*�u�%��;8������]��|-�R�?wJ�A�#����
��N�*B}b��s4�;�s����?�1���!{��r�1Lг��5�F-���T*�Z�,=zw��ё(�~ل�ki��^5��JIP��_E9�������-(�mg2������M��ߖ���g�N�d�hms�6^ĺ�ŉ�WE��?� �Z�6��h�5[��X�Di�V�f.�/G�#�2x Nz��h���GH�w�u�����4��|$(I��oF~�\�oD�Yk�_�i�sz>ڃ.�c���!���M�� 4���1Uc숤cxC<@�����W2dw�{�'֞"�p�H���\p�R��X�g\ܲ��3}�e��|�?U���FR�~ 	��(>����}��]OF�-phT�43�f7�\C�xZˋ~��;w�k�����k)}[���ux`JV	Aj|�%�������Q@,/�Ge�i=�b+q25B�h��%��&�#o!ڙ�����C�W��])<��7�w�f���Z���ㄧ���@Ԝnq6��bu=�Fw��g�P���ʙ\!? �;�<1���@�?��-tGw�4�w�*bY����vj��n�%���ǓO���'F�%��t}��w?g	)pe�ئV��O���>��Õ��c��Ck��S�%��ʓ1���6i�F�B%=O�3�2�lLe�H����Qb=�țU%c��j�p��L:c�M�FN��R��k��a�j�c�P��1�#e@��l �Z��Iz�TyjeF��bkҼ�������$�#��;s.1Rxn	��e�%����j����̓�@tv꟮�]�<�%�i�=��u+�ab��!e|<O0����V"Xah�2}��!bL��I�O��Y>_sQ^�!АrMW�EQj�����(�u7���a.�����z�f���/�(�N�[cG�q2,QA�$��T$-7d����d�Y�j$%0�\�!�?Nﮊ+��l�PX&�]�
:����ї�.�2k�L�qh�2"���w�afXv7T���H��)��%�๘��wQZ���U��y�~��2� ?�m��v~)��BP���~���'��H�ͦ�8��Ur�l�ԗr-�����wYu0`H���m��gk}fW���L��4���'��d��l��8y�O\. ���j��O^�Y١�A{X�|E�@dy_�FD�r6A\�l���W�� ��WXZ�����0p��J�&�d��}Z֗�P�����:��gc��m�_ ���N�_��ʉ��LS��Մ-��+\5HwdTf�,�3��@'W��������Z��,N\��+3��IĿ�]��O��1V����%����S����ǃvD�U�$ܱ����6s��W�x��s���ΰ�|�]Q�.���W�U5��z{K��kp��Ѫ,~ H�U�~�^[�d@F��<^n��!�Ym�]�q:~��=��}���U��[��)l�8K���uSxW�.�8<�h����D:�?�&��Į�V��w���7�������JtOb��w�pL{����B�#��;��gv:�.}
 ��q�6{��r\/�-K���vt���9.�7��]���]u�v�mj�z�|���%@�@q�������Y���o�鲴g]�1�-��W���� %
 _&e�z�B0&�+��c~�TRQK�{r�/�L��淪J���V����I��a-4Pһ�<�KF�R#�OGݐ�^�_?��{��2�\�QmV��)����ғl�K����4�Q��V�q���?5%�"�`��d9��+��gB�*�&{��2��U`�K:�.DZ"��9e(	��Ҷ`.�T��+̥�d��vm^)��6a���ڂ��_�M�<��)8�����/��>M��H�P�آ �T`��݃$t�t$�**]�m��
;l��\�aj���6˾w��	%�pD[�n������=Л�do��-�.-K��.�e����F�:���ղLz߉B!�h*�lW�U����j�,�A�������-�tg� �!�Hb��Uz�z�nC��@���9ƴ�gS>Iрޞ�e<���XE�3�~ �|��C�НyoS�M���FɍўO��n(�ᛏj��ܦ9����n�v�ݞ��*�^�i���\�_�q�)��$qfi���
)�N�4n�P���������+�g=�a�A��Ը���ie��_�}8Z2�6�*!�AF{�
^h=p�̪�ĵ�c0o/u�L%O�FR�0`Y8!��sWjՁ���3��c��'�:Z�aZre�0=������K�F���-�~_�����0�.�%+�h=I�Q�,�%V=��A�kc��Y_���h��Ұ")�Qw8�{u���fmۋ����(5mS�[X҈L��5-q)yy��*��w-�5g��T-�{�P�,�m"5�|r�M���܍�p�l�PޗgA@�W�/5ʏS�[�%V�&�F�ᗒ�9l���UIV�6X���W��i�H����8:
TUq��fK΅Wݒt15@�aJ�W[�2����;3@@���+U�η��x�b�XP��Q�bC�t�R.>1=�&�\����'X1��o6��T@�3�	�;U����UH͒��+G����UK�p�|��ٽ~����*3\6}���#�y>��3G�f�����U�w�H�.6l�h\�J4Ոsg=ۙ�X����NBIb�� ���}L�eY��l_�%���a[�k���x�;L�F��Z�i�L�_��q��N���'�)�(��^���ܛ�ۣ�+R�W/�&��棲��Iq�������a%;�T/b�>�<W���AFx^#�֪�'��f#�H��Gm	�p��P�A�AV��	\��.���[ג�y�/2	T�1�;s�����~_��c&�b�\�&��3_x���l��bʣN��sx�l�<��b'��^��$sSEs��Z��´����d>��~@������E��eH>�Qk����ɸI9��(6_���,?���Q5t��v�=�	v��bl���"oʔPx�K��lQ]%��6��,:8xT��|!m�C�k���p�MV+���+�W~5��l��r�����C��P1vE,,��^��I�F�_#.*-��n���;J m��U[c%�r0K��m��Ro��P���wr4���eRm�@��-�؄��L��pn�2=f��ޕF��Q�."2>�Xa��Ud��#�p���{��]�QR�We�p�����g	��s'���>ސ��j�o�Y:�(3餩tX5ȾX'οz��v�S�Q#Zm*���chk.���(��:l��|E&o��XJ���9Y���_�2����w�>��Ohc���ȩR��"'ܒf�/)�l!@��9��pu�\箛�O������ƈW��X6�`�w����Pȵ�J�
Ɔ[8>����IE��Lh���Rkw��bHN�L0
31{d���l�8H�/�+�&����h�Ĭ�x�?��+�ũ4BE�ک����PR�6
oГc���qUz79Y�OnM �����G,�҇�O�X�@7�I^4��Gn]"��.r� ��i�n;���^c�=�nɀ�#L��<
�7W��B�I��,/�̿�+�x�>�R��%oJ(
[h�U��2~y����	7���ֳ	G��&���-���|%[?�m�(n����59:P�f�	co�-�䒴}Q�y��fM`:��-��/��#����F��]#�ɴ@�,G��b�m�iQۮ��� �8U�e8�I3pS�l�qJb���V��"�8�4�q`���%1�l�1X��c����7)�!����:2#��L��S�)q��X�kϹg��2f3^��{�'}��f��P�׏q�7��%T��_��i��}�1�����~*i�w�](Ҿ 4��r�]@�O��Im�L��?���.C,��:p�[����HV�je���=��/�fm`K�W�z&��7l������Yf�M��*5C<f� 0\���ִ|Vٮ�N(��"�>����c��\$2u"L���x)]O�h�7xL�"zB�řr�E[�%\���dA���׫&J��9�L�P�i����z>a[:�6b�cy�h��f$ �+z��7%oЦcw�u�Z��+%�ړ��s�+�u�n���Jz�|�9L���c_x#�ݳOkZ�0�|"8jq�,�gm�ޙ3b䎜vO:7�\�$��b:�i ̑����k���!�8Bm:��2��x���C�,b�u��Yr�fe�����>J�o5`���47L����ϓ�^S�Y�O�iI ����̯+���u������r�6N�|��ZQu�O�q���?��M�q<�)$`ӽy�We�ąt�V��[���#���^K/*m�:>�v�=�ZZEH)����.֯Ԁ7��oX�`m.�Bu���2G���.Kw���~�kH����	�G�4��'���D���v�Uó
o2|wW/yˊt@�����?�%����8{^W����@���!قf���CV���K�L�p
S�oB�̗��²nv�^��>�m�8��;���o��fR��hK+��ғm���U����	�O4�{�'��.�=��s.��Meo���o۷Ew�fw\;�*�˷ �=��V�q;�
=�C��1���[�a����=�93B���RS���M@��C1F����1�/́ɅIDx�
�LNI�.�%��,��>J��
c �z����< ����m1(�Ce)a�"����^�2 	"����nu�:�Ǒ��S^P���
�3oKHP4q��Wo����ʤk�*���0 2y3?���g���҉����tòxw��ʦd>�X���TQ4�2u@��3 ���m�C����nY�1�0�F/М�	��.n����aΧ�J�83k�8=�z�,����>��s�I��p/�^�O�a�E��Z�s��L$#��3�x�C�~Z����u��D�7 `��I���դ%���ITY��,����U��d�ځn �6hU��o��L9E���*V�h�"�n����4x�0C{�u�{��Ϣ���Jֲ�A�6o��a4ar{���%څi^�Ѩ%/�y�Y �l�M��p���qh��'{� ؀��)����C*C0�Y]Y�C�=&��W���x��B��R��U�{K�O;���"I�i�~��6���pE�(�F�\S_,��~�d�&iv�?�Y����	���0`C�z.WM"B��j�ߠ���-)�x�P8��hz�^���Êpg��%f;��o�v��;�3(~h�����EqDvt���l�(�/��O
7���s]�B��P�}�V���n�Ċ�κ���K�T�x���)��M���)��jx�ڀ�ǥ�]�_\���DY�&6^@(�����=�>��c�N�]�~��ӝ!]��O)晱�3����	A]~�4��j
�8r����Y��<{�	x7��_NnϑTXuՐD��p�F�+�+��p奓`����o���Ag��S��`�sL�~�j�q��e{Fj����2QE�;���>�4L��"I����-�6cmV��P��&�u���ձ�@Z<ٟ��n�����;�08�����8��r����$�o�M�N	�A�1j�.�we!�z&U*.��葋~�佲;-�C�ٳo�cd7)=h�9��<T�E�Gc�y��(�t���'n:�!�{sG�&�X+�XL)2Y�T���0_��"Rװ=e�^Y�?hޣ��W�!�c�.`��XD���
}=�/gh�Ob�B�g����Xgy	�cӘk�~k�Σ��Q��?M̂��u�%�8�R.s�>��� ���}�r��>Z��F�JE�H��٣��/Y�����ѧ������O�&$���ृlP���b����M�P�D�L��0��@��IL%Kl�����["�Q�q����z^�vuT*Ȃ"�;\5.�X=�k�I��y&�7�x*lV�l3#�j�6���,�*k��:���#eǴ|M�R�"	�I�`9�ꡜFİp'�b|K�'PUט��kVJ�FXe�-��0�����	��5a�M��_4K��xYF|�����c�N���_/t��+��~b[��l��%y���S�8syAC�"9����Xn�����lօ�ʿ���"zAT�d��p:Րq�U��=�.w�f�&�����#7k@����4�¸����CK�k��i:���$��l&��Gt�������k�8����s��-��/M��LD�C�R��h�ڊ
n�/T�̿�F��b����������&c@�c��r���i�z���_02<��� �~+9�r�P���LSw�
G��M�Q��	����"�@-4:q�w6;�B��o�[Ww���-����E�H#�q�i��BU��g}�_�ƻ!w���P,ذ[�e�o�")�l|��̷}����4A8z@/H�92
�7�>E�a�Ύ��m���%�LoW�q�=�������-K�	f��*D��_�1��P�W ��S����l�v�' qe��jdiFw�R����;n�nC�h�ro�o1 ]M4�?�#�%K���_�J�q7wf���0�$/���5�11g�����.S�2��*�}a����p~�;(5�4.�Y�C���f@kv􃆎���Ŧ!�c�?��*����nVg�ķg�Е�� ��5g���:�/;%D�Rѿ#m�%�e�c�0��"\��8}��6��iX�vS�����2<j������ʝhh � n�[@�`*�S"k��ޕ����#]��4�W�r��J�5�����b&bS\6ii%�lft�0��'�.������I&�X,�S�ǧ�'�'1WXM^.X_5��jp �f�0\#{l��Tר�f2�����̯*�-0v?{2u,��S�
ES#)@֩���EUf�_���{ǫH+^�gz���D�O붸�P���A��Oݺ��<���E��jL��`���la�3\�5>��j����U�����njȼ����]�qC(Yqf�8����Rcqz�K6cl�e>.D�l��{�iЁ�v�@I�ws�>�1ǉ��CU�H�W`S������s���#�O-I	��,��f7h�ǘZ�Ʉ{�j�1�(��uaa��ٝ(�K4=�:�\}�X��(�����+�э�𕕯� �e���?��Ra>�Ht/ۯ��Z�Q��$��S�Q[`J�zR��qB��8g�ߵ�Zh�@���4;�J���:����w!���s6'>C��d��\e�w�-���Wnr>l;$Dy�!VS1�@/a5͓�T�
����gy;��=�f���}��I yVke!��^^�-P9�^n�oA�WV.�~UE�n̤s{ܷ��
�c�J����@�ªv���u�t<��g�n���hG("'꺂K	t� m��hܦ��G[�~�T�K�u2�|�|VI�Vf�;;x 	~�݌�=�F�a�0X���伫t� 2\��M&�w�s%���q�P��$���S�j�����'U��ڕJ��Jc:�u�޳�¨8w�~�N�f��"�(� ���+�{�S�-!,� ��l��y ' (���96.��u�\29�
:9�͕�CT
��RD�h8��h� �ꉸ��#�Ø��8+}*q���JK��;�_s��j	�pm��FM�9|���o��X�w����?��]��o���Ԯ���끢�)�6r}Oog�Bi�ͳ����{c�Χm�趌>ߠa���iXXͲ� /a,��-�!���"Ȣ#>$���g��I/����@r��0Vd˜�E�	#���������<z�[��/�7M,���6_�5r��r-cpʃ5/�x���@�Q��{�W<��Y�F8�SH
��90ɀyȨi|(74o���G5�?�����%٭�L)0�2^�x�y�Vi���y<�"�Y�[����w̍�8�)�<�Pۆ���a7���D���b��b,�2d���X�#1;���~?&��$���g^��o�]�ۥ�`P��ƅ]�rlKU����G��n�CI�m��t|>Q�,9#��k��I��k��z�v�k�]�^�7�4�ՐTU4B��;:D�u���Γ�!*w���e߀^����蓭��
U^:�൴Z-�/#�1��uұTn�ް�B9�UR�l	�2aXD�PNqF�Q�bSmP,}*kdͶd�eH�`�2	f��0ڍ� �T�~�i�yT�ق�Q��!0U����Oc�f�n�m��X��H�{=��ΰQ��l����]aa��J�BD�I(]s���+�yR��w"v��[�B]�� ���s�{>t���]�����|8FK�����q���٠������Z&��o��1�C��z�s�pƩ,�Jq��� ��������(�µ����zP$�8=y�=&�z�����_�?a>����.����4�*�\p��m1*`�}�o�sk(�VN��lwIPd��8U�����llA�O�F��X¼6��h�DStw�«w�	1�V5�C<�)�1�/�ӿ��v�{��Y�����ysb�n	35�Ǔ�9�X�hVO�m�Ri.�Zq���`�2�U��������K�1��	lԋ�%J�9z��]z3��;6����Y#�a#.���9��SV�/ja.�'N���K��M�h�,X��_FF6�Y���H�V/=���2���
�\���q�k�P:8 7�L���~ټ�3k$�y�n�j	�:S�%q��\���'G�c��ߎ9�cr�X��R8�5@�u%�UjL/��4��_�kvI���S+��D��TF_��6�Q��W�\��Ti��o��x羡lm�l�֜Sh���#�(=�m.���WP/����]w 46&���e=�tզ��t`/B��H�������������f�R�z���x.�A�Ņ"��E��^���G)U�IWD�2VK>�:��<�r#;@��;kt\�,x�F������zj�Y��F��r3.)��a!mꐎ��O�K�-�G��H.�p̽����.4}ʃ$�������v���������.��<�~Zy�4S2��a���:P��U��^M3>��������]�C"	_�*��ڶ �՚1J�!-4�B�S��4�I(f}Y��MN�R�~��K�"�R�l���nR'�y��v/ĖgLM�HlĥCƥi��uע�q������n���fzL7Y�P@�E۲���[f�z =)%_83���e�����%­K�-��A�4d�*�E/CtSE�YtV���`v��[��DUy�|���)����=|�����mޞԶ��>��������!�4���S��H�`�[�{�	>J�]��A�8E��M���/�
�_��-'b �U���������,�K�՟Sh�E�@8�n>�j������E����\z?�'���6K�:sKe�����h�r�]����"�UQ|[�f�<uc�Ԛm�C{>���n��&�K��$� C����5N�W���qTW)�.����EI��B=j>lq(�O�|f~�|J9���*�)7h�x*� @��}'��c���_�fg6	h��L�K*r��z-��W/"tN���Huڇ�Zk�.��ʏ��)��� 嵴�F˺�L�0�15y廟�7���5�U��7�-L��j^ϙ'Z�<����w�A���{���(�ZA �lE^/�X\�#&����.�E�.ӆ���o>��pJ�N@E٣۪(�Z�|xK�i�k����A��g��+����uL�	�j�n�`W�	T���Y�!p����BL[��Y��
�3B�s]��O!�d��t-�F
B	��x*�<�hW�^�xp�뮫�=ء���=�	��l�i�U�;�B�ݟ�c{��/���}�`�����Klr�TT�2U2����ry�Q~8%4��tt�rH�o���w�(6�5E@�i)�Kg7�Ĳ��ߊI�\ⅲ��Ԓv�7��vb�={�z��{�d~8*����rp�0S��;�N�3Ѷe	 .b�q�X2�+��Џ�:�u:	�B��O�����v�):q�HxG�=�ERL�b�&·J=�bs;:[^g"�r�\�R�A�PgT�y��3i��7�������^�G�&���/�VG����'�`k���*���׀���fe�.�G��?�9F��g������rΪ�����hޢ;$Og�D~���f��%I��M�]�$xX���<oZz<`@lE�N��$����2	�oqƉ9�_Oe� ��u���~��Q��� ���~��Y\^D�*�U�3�0K��y�C4�:����e×��<ֽ�N]<�z�J��s�fO�܂F�o���+j��c�8D�;��þ�5�]?[��<;F`O��������sPv�'��q��G�h�H���\�,FW�v@���r���b���.��M�Ǎ�����v��#��#�!5�;���$�Y��95"�޾a��w�'sg��>k'=lq��*
�
�����&z}C�H��r�� �!��\}���p������v�o���� [X��,�r��'�%EJ��,7x"	�]*9r��F���MbS� f�������]��_� iPc&��'���`���S!Ħ?�8�,J�a�[W���@�(,�d�0�Ã�Wt�SI�!�1J�z�e��C4R:'9KM��Tu��p�-/,�Ju���S��,��e�B@G8\�M��C�B���n���O�%�Jyd���Z%FO�ٙ��3�k��S7}³$ԣ���`� ��'�1��gL�t�GKzW4�&���H�$�m�ۊ�ޟ,=�F�(���43\���b��۴��?�T潛�`M�H`�8ބ�X}������6W�kG9m�2 �hLO�k��yp)1d�u1��h	����Ow�X@��fn��R�`���M��QЄ%\1�e��W_t)N��t�X%��ݼ�r�����J���t,Sq� M��HK�P[Epjy�ut���(��	��ڋ�N�@{�R _Ŗ�mIB����j��۝�]#Íz���}Jca�{���@��9Y��*V������7ת���f�	����H4��a���K7��%S?�&t�,����H����g�t"��L������8���qc�TSH�aV��(���2��?�,pŇ�@��@Ժ�wC���S�$K�����q'��F�.Q
w�����jV ��n^����P�{�vA>!$mҌ[.G|e�*s�Fl�1:�؊M�K�y��z�m�-�k�L��=��F�Rkp��U���E���}���Bw1+3�Wj9*!8�;�ڈ鏽��d;'�a5��e�],�ڜmxP>�Ʋ�>@5&�w�:m(�\@��FG6�X��'�܊wma�kD1��FB����(�\/#�M��1�â��֓8$�/5���p�?>���6�{WH�A��#��U�@�`�:��]��y���>��XѺ'����).��*�3U�������&4M�}O�X�`�E�/Vy��_�p	#:�$�����x��[�FO�9˛��0�5U���?(� �kB�<�Y��)�n��p�M��UPf԰��I3��;GJ�c9v����V���g����:X����A��t�7��S�=3{p�o���I�����k\D]O�2%<��g��j��z���K$H�j�S+t���X�?��j�҃�~��}�Nf\�y/\Q+ <nYL.�Eu���ٵ�xyy<~�|T_q�C
h�U�<]�����\?w��ٺ��3�����l�S�u=\?
�eίtj�w��߁/%��6�ǍE�+��� hm d1�L�m52�o�\���,GU�t��u!1�b]l���GҗEvִ'�]��)o1�3-�DC�ḽ&���=�"�[#��I�3�_���fg�@Bc{y��a%��;/"�Y[�k9ǧ�=�]fͥ:��!¹W3$�-V�rIi@9B�҅3a���rŧ#��hg�$�G`��(c��՞�������D��`/��4�h^<|u�����{�jOF�`i�ɝ��BcՖ�t�~>$UKEB�C��m%�g���L�%}>
�1?Z1��}��*+?��f��&�RT}��"T���&�8�8;��f���ϭa����RRW*��������xe}��uEp(�r�㹙[�c�U�g6y����?Z�.6���o������yɣg��?�M6�3	��_�q���������'�p"%?�f�|s�W������?�t��?0����/���?-����g�b,�I����:�~�d֣^{�C7DE��^�n�ry�C*V��:��ǲz;\��;���k�/q��t��1`v�ˣ[)[�|݀V���5o�P[���|w ���8^����M�U��]������/K�a~j�i޵bG���j���0�řw��(��d�v�����f��(�ZE��:SR�\3ꃎ��^Fb��Mr�ܼ�F���!���%��ps�y�����c̠-%C��rjO�sq�0�^K�!1��H�����c�b�)/�	�#+Cj��F�S���5nm��0�3�,~��o��Դ	�2��m���=,�L	��I�i�M^|�!�
l@�n2|%���x/�3�x<~�"+=s7`��/�Y�0>��3h*���'ʇ�!l'�s)R��s�� a2�	q�K�&L%�!�
*(���\�q���9+Rk��7����%��6KSEd ����KTo�������Y�oB�m��<����A��h��K�~%��N:�l�|����Q#�1Sr5hV��	��P��rob�d&�ӟ0H5,��ul�}�0rhՁ&Y�Z�|ى3vhɬg���#j'�<T���q�R��J�s��<����$^jHR$�����r�jɪ�PH�	�4�e�;�p��N,���'��*6�.hyyd���i�=������Ij��K��,K�s����W^�X��^M��C�Xܗ�֞�a�_�H�����,|������f����\:~Ela��L�h�f쐎g��m�������!>3��k��i�qy�*7�e
յ���ɤZW��ݍ����_o�ѣ��a��Ak��d��/zf(T$�*~��7���l�Yj<��Ԏ>�$y	��U�e�H�̬�&��Q3Q�Kf�������!>tͽm���3!�/S��Sy���J��V�@;>B�r��%`d`�k�ɞ55��:�&.�::��t�ā���$m����x�̜�wT!����+6ݕ��#)ANwW�~������M�?��Z��=����ٻK�O�z?�tI�ԧw��vn����7�[Hu iŤX���$���
�h\��E �Z����r�]�$^�N h�` R��%P=��x�� ���j�^7��Pc�s��3�'�����H�U̒��/緒���H��?Ԛ���#�.��A63�"���G'�ǵ���8O�u�~ݰ�6N珋��������[I�;�W�i��{�w�rH�~p4>�kt�7m��[j�n*�Z���zK� B�-t<U�G�g��%9E�?)f�s�^��تzH�����Z�fBnZQ��8#M���?"����H$���\Hv���^�Y�"
�0Oն�]�S�kvw���IJ��+d-�(&H'=͍|J5��W2�!\s��/�8���rGJ�W����]�\U�@�'e�8J0)s8c%�9�T��w�&�=��Gm�{C��q3�ީIE("�ٖ�;%Y@�&SOi��E�\������G1��"\t�d�}�Ek��xfps�#�yD��o�"�2���`�p���o��-�֮N�*jeq�
~�VhC<U.W��G�P,�����ĸ{i!���4�k�Xq��uEq9.<w���/�p��q���)N=���,K7+?D��Y�v�}��$|9'��$���T "���JG��h���8�!�Ӓ�[���.�L���e��Q�qޢ@/��k's4�q�;YУ�U�	 ���8��EF���)#��	%����l�1>k����m���Z��^=�*;�:X��D����ݹ��9�T(&��C�����s>Et��{= )u6���r���B�9���g�rS���֐<x�O���S���'��C7�9������[|��H���P�{�U�q��)M�}�攥)Kw3g�r@>�����Z��X
@��d��}2�偘3G:����E50�*�������[�D]��Ar��#$�BR,��GR�2p�Ed����v�/�-����j��Ղ��yrݶ�,�
~��������+��A�a�N�8�<	�iݐ������u@'�#�u��`.�����]�VB@���ᶺ��'�/���X��4l��S+���6�n�����5?�F����w�}���8ȳ�@��mN~V��.[H���{�e����]��������o��6ev����D�Y-`�u�Svl�Љ��4�y�	�C'�wn��D�i��b�\�Kt�������#nYH�Q�Tz���S�"�yu��@H.l��_���PTk�	���e�g��8�Y �G��*=D�b҈��[%�.��|�\�a,��Ƅya>�b�S:��-�z���hX�I���;L){�tBo��8ش��n�D�Y6��eL}?C�`�+��ieV�����6t-:Y�m~T�� ��&w�A4� 7����x�8}�!�/X����͋��_(D�3�+9�_K[�Qt�U��!x4�tf�Vx).�����jl�,X��mp�iU����֗�]�	o��E�!ȕ�.�������B\�`E��)����70��F}O_F�swv�(�[�	GG�f5Λy����E��²V� �yJL;l���'k{L�J�\����`�6�nV�Kn��@�:���W�8A����	�/1����Y>�+� �4cY�f5�?k+Oi]��S0����ìq}�#�Y0�WA��1���sM	L���� �?O��&k�����r���y ��г����LM�wV��C�6�u^H����L�/᱇$Fm����ᗖ��7�sj��f-�}�̟~��[g'��k$}�3�D�)�^����W�7����mPc�w���I��2\�2$�|�2Z�qKr	�#L��o�i�2"І
7vT&V>�_0R ��3۽�Xi�ʨ�?��9v�ݻR�Azonb�/�M睁�t��:l��?h*]U��J���<M���XG�([4�`XҼ.�4�ZO%��Fڽ����\��T�z���:�eo����fmho�:������� BP�yr�4{��5�����U��[���YOpr�34b�3$�����PW�'������@��=r��5�R��xLP}B��j��h�ĂB3�1P�Fk�c���@($��
��������Q %!E?z8|o<B*�o����$�<T�E��ݻ�gA�L��8��->�kB�"o��!�}��aQn�z������W&X��x�?�y�
<I&P�������vU_����bP�kѯ�i����I]t�R: �]V�\c��p�!�,7����e�ae|�t^�?�a�� �2X�k`n��[|M�dA%/��-k�:�~�����Ê�Y\�,�S����/)k^q��6h�bi�b�P����o�^��s��=~�J�0>wݞ6�o���c<�֟�l�;F"J�`s��O��DX�Q�zڹx�?;��tV�H�s,��X�~&^c��k����.�Cu�s�G �]n/U��:>�ʜ�A#������)ll�،S�@Y��T�:�ZJF֥�޳�ɞ���Ըn�<{��K�ҷ�9QǮ��(ӀJ�3�+)�
A:����ڀqR�gu����e�O�*-;�P��é�@��(�".�"��e�V̥J���ϗo6���rO�L�U�)ٗ}� G�*?�]�D�M���E�!��]?Y��D��T����{���P1 ����p�'^�V Ot�_�)�(z��J�OyU꼽4��U���J"2գh"��]vG7\K��-l*�8�$�%=T?Z�Ԓn�=U�ӈ<��9���z�C�����������a}g����5��/?������q�|U~У���[ǘ9s��⼹.3- �|��E������Pr�`l]Ӗ3#��O���I�Y�j?��'ܭ��8�Q���� �O���B,��Q�Z��m���!V��޲�q��&�ݿ
l�$[8�"�s��{�����T�ҡ(��V1��&c�ӆ�Ǳ���I��4c���ɢ�G�1r)�YT�;�^�*�.�\���a�<���y��J���:�Ck��p-�}�+b���L�y~���}�ã��.J���-���O"s�0i�u�s0�g�����nmr?j����;Ń�|�f�c=A��U��Lu���aO�(�T�՗1�KQj3�<� �urGK^x�l���ʝ�b -de������)ٴ��+OQ��./بᖄ�f��u�W��I�kܠ*�P��w���mjt�h	hw��
���X�o)������R����!�x#e��]��f�0�'^��ǚD�;\O��v��"��7ůG���Cz�Sl����tZ��Èk@=X*SL��I+���!���U|Գs�)�$Q��;��s�&yj),� {�+���FQ7��8�rb�8�I'���r�t��t
�_�ܚ���a�ϳ|��C�8.!�������G\pd�<]�S���Dk� ƛ�xdz��@M�hs8q8[�κ4���l�O�P��ep�k���p	��S�\�q�.�i��O��fv��WY��|p/���]���Ys.V��W�>m�}���D��k��N��y��%�]�`z��iBFq��8���;M[}�8{ �R��F�1�M��.��a��(2��q�'�X�v��V��U�%��H(�ض���6
�[2�UBvb�J��]��A�=BHE0]�\��aO�>ߞ+-0����Z���&��i�����X��ǟnp�]q�]���[].!�V,qG�����1�Z��N2:7����ۣ�gBZ�WV-i�:���`��aT�?�p��A�ۈA��8�l�.�~Ya�.M�+�F-X�ky'���)�m46B_���w�)�J��j�N|�+������D�	R�;�tj�e�m/���P�~=�>���1r��X]4�c��K�8A`�����f-���-�.i~.^�|�[� �
k�k�h�%�Lr
5�}Nٰ
�����&�(�#&���Z�\P'B�[V��B�-����n����]��O�P1=�������u1>`;��ά'�K�-�o\.n�Kw��U*���������V��I>�;�COH+�y�o����}�h���k�Adx��dz�-�z�,X1K�.0�d�w#1�`�k�Q���ĳ�lN�%���=<�V���$V�����ɋ��8(	@��h �S��Sv� `8ba~9�i���)�:Ш�P�Nf�?��S �'~��&�?����3�=t�_'�
8��k*�L�F�ѱ �錍��m�sV���~�Iij]i
�VC���5U%5��k��O{�UX�
�6���w��;�����ׁ�2��l�'���H���0��X�!���x2����ޱ#���ks� �1e���������u i�	Է���1���#'��F�`��Yz8���Jd� ���ȑ�r�X�6�̟�ۂڭwZ��o�l���?C�x}q���6�\%�~�H������D����K��:���xL1R.�x}=���3<����\��Nr��'}��=OT�Wb�U���wov#�d�3�X0G��,yN�a��z*�vn�	*&�
}���WH�B�0ؿ�tIͦ��0��N?!f�?�Q��R�ڦ�Ȋ�S���{)E	3nc���BA$��Lq~ ��@b�0i�*8�(	���;@HD�S��qq8rVl�ʯ�y:W�b%���x�������w�xըV�S�o3pO�9Tk���!�r���%�j��hD,�� <�`0����b3ؗ�'1ϣ`Ļ�B�H��Τ�yY�Ů����vE��Q�v�j-�2��J�bѽ����n���GX_28��{)���<0��+iy�A��j0Nk�v�_D�OM��le�W��6q��2��&����*7-_�T�\f���8.����7uaZo� 8ډ[{o��Oނ!O�U9W$�\M��� �B��� ��=M�eb��^����9����(F�gև��a��w;�b�"��災�����e�j�0o@`݊F�����}J��\w��,��n�v3�l0�(�`rC�
eaUF��!h��7s���: %��ad��yr��aC���O1�&�~�ŏ�\ty܍�i0�m$���yU�Y�u�l�߰;����͆^�x��_��d4������^0(�(�x<�,=>=�t掳�t�ب��W�{���]�Q�LiX� TbI�mMQ�e�5�=��b���� c	���3�?7��(��	ъ�eP8e~����(<���XO��|�0�,i�7"��m����v�j�2h�x�"��ò��#�B�N���kY e����M@	�8��A0���k����wWa�Ck
��\��)�F����m��9����O����-�PY2'�d8����������?cC+4{L�O~bk�)�0e�2{��q*�<#���a`��_��I���ƫQ�k*��������>� �ڒr�MJ[Df0��������O����?��ߥ�Л��s��9j�\�t���n�ژU_pvKB��:Yʌ��s���9ˈU}�7��&�]���MZ�='~e^Y#8x`?6e�^y_̨P�߱��[k�E�Z��-B�,n�T���?�v����}�O6�e�Y����j�1b��#xD��2zl7j
���ڻ�k�t�ݢ��hL�/�L*���a�mj�����*�m��-��:7�R��sb^���y����ԋ�������wb�}������i�ry!�����Y�6%����^oN�o�C�V������a:�� \al�M��ԉC�-�َ��SW�q��/'����=��p�2p�UX�C=xB��+P5�R�_��eY�����bvJK������2(;�ۼ�Y��k�S�UH�ZTR�6ϫ�Z��9	]�V�ÿ5�p��U������+�����X»�&�!�
T~��b�W3˫���4c��3t��Bq�0 ��AS k�	�g.�c���s������BC[��w����l
?�Gp}$��(~o�R��0��tuF#��b���y4��,*��lM��Gv�+H���e݉�$�q ����t��]�N�υ����spw`<Yw\�ۄ"9t�2�᫲T�w=P���χV;����6�Nl���70��=�},� ���Ǟ?#tt������#./�ۙq3�a�)�L:Q�䖂���7@a�/�hIT �j%N#�)�	հjl�"��D�S�V#�A%X�rR����{�R��a�7�j
.��u{���C~�Q��H$�dI�[I�s�U��#v֛��r/�
�OBL]biUM��=��}7�����:���n)���AXhT��<����.z��kk�R�̯�/��q��6E�
j�"�MV�᳘\�����WGH�W��@s��ܿ�]��7�;	e����;�g>�"��!w<j��4�Ț�_�^l�w��wx'D��0�8�mS��]����Go
mLF_%��Y_�\�������C�\��"%- s��*�c�4�~,��:Bl����%�'�@�rb�w~��)<���ƶ�T�?.������^�m�85:Ff_t!R���V6�L̪Hs��.3,vC����t�0��6k4H\y�iB y�
ӽ(���kj?���EWHU%e�⬰�!�E_32��h�(�7���85�H�T�h����'.[�N�G�	���aO�]&�-		f���~:���;�����F��e�6;�]��9��Lp�e<v��d���Q��7�R�V84Ldh3��2�Ww�^Ȳ�Ee��9d;�(���}����3��>ާ[�?�Ɵ����Kz��|�o�^��\���E:ZLE�����	�#�a�<�X��}�����]�\T�òe��9rڻj���54��WA��v*���^0l2K�)�����S��Ԭ�CDMd0��^ ��r8T/X|h�<���yG�GӜX+on�}G�o�(�Ǳ$��ƽ87V��ͨz�s�i(/h�q��m����7��Vv�����CK��s���Ԟ��E�n�7_JOQa���G�ӡne���m����
 ��G5 �h�j�����h�[������NRJ�\w���z�[�
&�@��
���OQGi���n~�I�Q�1�����A	%�_�\v��a��8�t�oz�Czq	H}0����U��.l�������@:������96F��k3p�0o���o"bEH"�9��5��!���g��w�u� ��D�ht�]󐻲-Ch�{������R��:ǎd�V�fR����PF�9�f�./�Ҙ������|���p>+W϶KU���3��Ls��D��:cz.A3K?D���W.�l)	i��' �hFq]��?5�c������^g���$��2�����szn�BPH/P8c�8�V~���DQIgx�J�J������y������4a{=���MK=B��P��65u�1���P�`i�\N������ �*��(��*Nq����t5�.��UO�v���W�S���\�5�&P�=�y�l
�5�ו��h�Y�V)�k���#���ޡ<C{��o@^��
-h���Z3�]��{��!��Y@���M�krQ� ������ī?h��:[�`ޑ��~�=J�rs%�z%;M��ؕy�����k�P�6��yU�v�c;s�~���-�ɐ�ɂ�g-aE<{J&b�23����J�C����.�}l}�`W'��E�~�ظ/	�ɘ�*��\��͔��Z~�#����j�)XW��H3�N�z�3�ՍtJ'𙃦��r�3�sJ0��J1+�%�x6���^�^/_�n����.�:?e�Y�O�]��:6�pȓ[$�^�N���0�ׅ��{�Il�MD�[1�;��A!r�����(��8t�f�U���h�������=�.�F.Q$�y�*� �0jg���!����zY�lL[I)�v}>�iL2R�b����y�ۈ������U�o!y����zXmc����\N�m�*Y��"���ơ[;�'E�g5�`;J�__wД��@�r��v������+a	FS_m���1�!f)C�*��x��c��Jl����/��!&���+�~�N�4ֈ	�`�� �Xw�>|L�:=PV��S����k�v���4�܉_a����Ì�o����W�!N��N��e��n�B��@������P}Ԅ��j݉�̮y?8����0+b�hb�h����^�-��{�0iZ�,��F��S4�����'mD���9��\iz�ʠ���(1�?+&L��EXr���f{�]�N�39v`�k+6^ndj��c��^粴z1j{��Y
���҄mi�%�h���}[*&��֜��VW��e�Wi]7���%�v�DO���(Tm��TS���Ҝ����I�+]
<�:�_�nF��������p��k�y݌�����`��&X����(f|B���ד5:�KP�$���_�#*R� 	.��	�bn������ws�٩�ĦLZ5����`(zK��D�!�|�(#Hi�V��~FfJ1�R�ߢ���hqN�v,Wӯ��Nd٨��b����L����:ڙ����R��9�c�[�hp��i�ESA�d@j��`P�O��ww{b��|�?6���x�a�К1�9&�Z��ǈGJ�|N�|�i(}��q(h����LnJ�(J��i�@��{^,JJl���N��J5[�\������q��Wu���82����pZ�A����
 0$��pt�K�	�VV�'��Nq�n��r�@Sa�Y�A
D:R�"�N�y���gy~e����ӓ�g�5:7DgbĀ�љ��!�
Vf�z�d�XY����M�Q'l����n�(���Q��/&�>��W�����R����=m0�)�Χ�߻2H@ZK?�%����д�9���ѳ�m���j����<tC��"��^�7Faյ��K�0�L��4Pf�Q��Z'�E�r���8�[\,丈�6g�	\�K�؅��!e�33s�z�:�*����{ҧ�[�>Fr�Ȑ��Iu�t�:����JQ"n���a�G��6G��x�f�iL�I�v�@D����<Ы�{�IW�}�"p���+-D��3����%��k;w��gsP�z�tH�����u�c�A��[fI匥L��(�	�6�E�p�@�*�N�������fe�����7�_�JK��d���h�sP��o�;��N����*��1�('������+FX,P�j���zR����tH�w��i� 4F���7N�p!��@4sk�|:Vʙ��[Z���n� �W�Q�e�e��5�5R�Vx���ӛ�Y�-Ï�+@�k]�JXS[2GX��<�1���3ژo�^��)J��n2�}_�wr�j������ܝSpI�'�q[�&��z��GI��1�H��"�돻�prɝ�G���SBE�%�#��y��t�����Cn���72�h^����5���L}s�N���'���/�C�ٕ�4���&'�����8ux�'��8�[�AT�/��*�P����?��o�hc'��������b�L���0{������7ˡ�]<��r�����k�����g 4^ I/��B��c6+�rܘ��~�s�~8>�f�EL��
�Py��!Є΁��jd�	,�������c������ÞO�ص#�7I��e�Cۙ�'�o�Q���¡�%��h�뮚s[-͟O4ky�o���b�7wLa/u��WB�a)w	^X�b�����1�8���E3ێ��;�������Y��j��c�x)�;l�����h��o�?�h�~�]�x!r��68��"kW�u�j��mu�v�0B�`�;�a�hN�"d��晴;�8 �@2��;i�����ɲY�]�R}��D"������Y��䂧��)B8p�Y=�芥M���\�b���G����;b�Ǉû��d�D)r�Rߩ�ގ�]AtK�G���~,�aOߙ?IVW�Ɯ���I�.�b��\擜�;`0�	��`5n|X��L0�����+��I��*S n�F^�w:�e�'Ӎ;&O��TZ�\���(Cp�B1P����^�n��x���"�W{~{jM־��'6pQ���Mrm��M��Bd��uA6�Ii��)"�?d���[��AE�v{P��п�)����RW���8K�Y�	���Kϸ��o����#� ��i�4�1+9��_]��ns���.�#%�n�r8��6�a�)``+(�Hbb�Y4~G�뒅�2*�A����p���N��iĭ�"��]/6Aa!Y]�Yj�iI�;z�҃Y"u���!���0UWu*�y�g^�|KGd�n�*�0yOY��{1̤��|Rxw��d�c̤�~�+͑��h�� ��˺�ǹ����^���0oAޡq�n�HlHw,Nʡ	~���rV� �l7=�vGP=���G8 �;5�j<�_���L22iR��8��:�+/�.�����X �Ѷ��p�oc��4��H�u��o|%)]uk�׎}��OHiȃ�Ť�c��nb���p�#�K�bi���� �q�qc��$����N3��h|�	�������P�0L�Ņ�r"�����n�y�LE�am�H"1��8�
6�Z��_�'^���S�2���{��Fݪ��`����>�7��Nج�2�=��ۿ6��K� v~aroQ� H���4-�Q4Dʁ���&f�.�+0*����s5��S��r3��m�20�U��g����RD�&;)�K�0�`+}SJ	�4�ؿ~�����<b��3q8�-Π��!jj��ݔ��$}�s:����4 }P�J�u�/uФ?�U��O�a<���ZfP�p+Ɵ0Fi��1�u��a��RX�I��)7��mᰶ�@�G�&d�>>)���X2�ؔMI�����tj���~fF8(��먊�V1��h����Qx��ˎ�I�0O��?����T-��ya��/��o,�J�6���
$��<2�@�A��䣌CK���0��Z�����E���Ԡm잙�/]/����*>]5�f��Pg����5�� �k��<�G����m�ɡ��� ���4���wiԤ��(9.S֫��j��M������`n��>���Qq:��e���A<�ٯG��1������Ű���f��Uvr{���L��,3�5��?�x2���H��W�L�Z��a��^�|�!n'���������Iv?�vB�U�&��I�G_V1'<^[�� ��+��n#�c������)��Q�h�H���%�/i�78h��cV�����2��}{&��jo���4��0�v�K6K�P^�jK=)�JR�3�b��C�H�"��N]�$Q'cx�~�*LE�mr�نO2<RX�� k>
I,5����>fӴ̾��U|f�K�ߋ���$<�J%�6������R�;�bg�"�ʕ�1q#�CO�Ę�C��u'O��o U27S��u2�����.����x���5ѽ)2�)Ժ4~z�{�����p	q_�u,�c٧^�7Y�	���[���A`|P���5FL��exfi
�S͊��g?&�ӗ'�v��DF�eI���*�'P%ٙ="SJ�tD�-��O�"Q"m���I�	�׃`��S�x���7��U��V
��lҸ;�\ώ�{�0�m��nP�W�ۊ�_�Ap4L^5n�j-��d�Pg��s����
D�}�ʓt狐}�T��b`9��z/��&�n7�#$�ï��/���;��"Ea���zK�dZt� ��6�}�]�&<�_J7��{T�:9в�@~���Y% j���
�!�E!���U��+t�F�3�ër�i~Un-�b.`��U���ja짓�$�_�h�Ŵ��E�] �
�΀QDx&���e Ww��tbx&�1�dbe|:�v�d�@x�M��.pOȭ�Z'�#������h��g*�h�˰ww՟+��Ә��}��l)HF��e%��_��{���I��OG��uj;�C��V���窇3��~rK�+^��Rc<(��Ǚ�h������G�
k���V�X���L��MG�=���oN7�MoN��tVv �
���7���@&�Sh	ӕꯜ���9�S5Z�U�Q�6�P��}��bç܄=*%�fA-��J ���n�(
%%�>�bUf��ߩ�hH*�rS%�5��� ����^r��<�!���/�s�0%��&�OI��x��2ø	Tݗ�,�	sZ��ո-	�R^��^�N)��5�ma�m-dݴ7nBuc�
�!N�x��%�S�/���a��n���2�_�c�W,���{��$���T�,�"�1�3C0-l� f0�}U���ȉ�ٛ/�'̅�Z	�f/�z��Q��3dT��y*)�Q}a��/[b��sʠ2�S����t�;�2b����ۓ��oo����Q��}�Z�7�Ar�[����P<���� �E#��Tj���8�!4�^�����>���F'�_`o)[�݅�p��*��)�d��^+C��W�KwG2���j��7�Kl� �M
�V^�JM���Pa�AF� �_���~F��@Q2�iʄ���s�O��������Rp���s�?۟�I=�f+������j�K��=����x�DX�޲�3�{�����`ZD�xJ�`�?��&_+P�%��=���H�a��?IyH�-����>y��r�P��̸���%Vx����k�Z� /'=p)��Y_sS~���͈W��U�9�1-!-]{��h�� D���Ix,a*���5�7et��F,q�Bs��(�t�^��Gӌ�2_�e�Z�T�����&W�F7�5��U�RʅUus/SZ�A�nA��"1�D9�_k>aI�z��tDC�	А�sy-�;doҦ!1헐���r��K��ǻ��w��6+&ҕ{�7��o�T�]$���}Ar�Aci@��g�ǄK�Ar��wd��,�+X�����'��V��.J�XW:j4�Z1�S�8&|�]p[1`�&�.{�
����9� �@��5��@ᅲg�cg_�P�&Z?<�#��Tى���(S��Ê�L,k�6�U<t����y�ڨQ}��'$J ^p>a�d�=�)�/Aor�j�@�,X�.�mxp�Ć����b"��+��z�Ō��Ƿ�@�WE�8���}Bs��'5�޷l*I�d��F8*������ZJX����������}��,��\�L=T9�`� ����L��7�,d�3��p���a�H��eYtu̒ �s�?��������N+<�r4ۡ�/Iw�Wb��+T���O�6@����+G<O5��"�{.D
~��7�m34�-=r��q�/�Q;�W�0��a��\n����-'C�ܷ�n�r�+�gj�"���1���]���'K�B81=k�8!�>du���h�6j<M.��A����7�]�v�T���&ij�T�{�)u�����`�/{I�FPx�$&��s(� .2�n7A��AQ��p���- uM����8�,�ʘ����3��2�_��g�F�)H���"�\���@�tU����I0���\)�((XV�Ü��!G����'O>[u�F\l���/z.t�M�u��Um��n���!/A��ɝ�<[&���[&/ �����S��p��F�Jn?`��u<��6N�1s�̽RM%��)��c��\�����*�d� GbM��f��$�'���0ʚ���Fg$�f����N5��6v�íz� �Q��-<�[��9"l-dm.�_�&%m8�5j�����`P�-��xSS��Ҝj�w���F5�gz�4���w�RXۅ�� ^��C:�06�j�]�+}}�i����N]��0��GT^�f���<���X	�YI�LJ� �c��E">e�3^��%�\�ғB�W�E���&%r/����{`�;�W��Jኣ�}��-�g�i�C�}���z�Y�&��jc��2Q�Ɂ�X� j,6T.EX�����YJ�%��R�[� ْFz@CM���]�$P:�[ʝb����jr�@�Y��
�����-��� wt@;v`1������Ӑ����O�so^s�"�O�ĸ83�� ���l�7:%H��k�qP�eR[ٮ�G���3��,�|����VC���P�`�J�G��jz��w�����מ�t�?~�o"F�-8��Vv>ݢ~gi�#ћh�����a�1,`]
c��s0~x a\yP���J1A
�Y9'h�tت"6�Eg��i�� S2/fi@�/t�[^����AJ$a*�JXD��w���sy�\����fGvp�cR{�+(��A����q�A�-�G8�v�x��XHmș��*3�u�+�HF�.��mQ]���&w���@ƙ^֚؋��PϮ!B-@�;�٠�bpH���ǘ��8L\�V�N�:E/��Ɇ _O>@훝¥Z�D�玠
�m��R�Am �Sf_ I�+y�����58��Xr�	�aR�_a�}tj^7��M�Ɣ9��TvQZQ�'t�N��z�c)|4��Յ�-���~K�D�RK�`8��lEf�N�4����_�X�%|�?5'���Hha?l�ۜl��ˇ�E�	����8M���|G�φ��I��Qcw�K�z�yWbLϗp���#6�����ZD�1 ��a�Jpo�h��n���KDB�#�P��A��L�:BYU�XT�K�@���x���8�Ã������K.�8��q�M)2�j!��Y��]���-?��`隼#�\sV�wB����;�<5��������d��x���Fo�J�����"�Ʒ�˲����Sa(+P������<� ��DQ*6�4�m{;� ������C���n�z�j�
/�y�/�b8>U�K@�LT�StI������'ցrO�ԙ�-*�c_��������&���yL��B��� �^W�h��!�H��J�p͂
�^��Z\���`/�����,��b5��6�#!�	�Q��)-��T{���9������2�E�*y�p�~"���8:����,�gg�
m�	�;�/p�Cs`lu��hC���2bk��5����2[t��ޔ���4����\�7Gq̧5r�E잣�+{- ��g�ﷆ�����-b�{:�as�`$�u5����3&�z��[���4p,4� 	�y���w���r�g�{/�/��z�'Sc=�Q>��L��Yӑ��vǖ�;x�/�������?;���-�-\��]m�gy�IJ�ʆdDV�hF�#���A��]_"w�0�$���C]ӹ:�����F�#��cX�������_=�K��
�4���������O� (n4���I��ʧrs���gc�U��.hӗ�.�o��c��N�N�7�S����=��9[�X% [4`�0jh�����m�7J�����ꑚ�_���A�{���6��yDx��߷ �\(���Gd@w i> ��q ��%�N=�x�@-/�$�KMτ�F���'����52n�tǳ!�2\֗��vÍ��j�M���B�WWۀ��^I'��A�|d2gr~������f�;ۆW;ȿ;�"���LB��1Ӛ�\���6{�3BR�mF!J#��2q9��s\s?��csMRt��	�R5	w�G�HhfX/°@���Y���L⿜yY�E��_��maɉ��J��I�pL�̃�!�8��uOc����Q���H;�PY�Tsڞhv�,k���g�s{�7Zр���P���!M#nGZf��7A$aw���6#|��iݼ0gc�P;]nE�X�֡��J�u��!��b��d��iKk=#��trb*`tV�N����]m��f��/�����0�&^[m���� ���QʼGC����)�*%��)�����L&#Y'��j�nM��ܣT�g��7�O�<�"	���j��z�9���&a�$��	/��o�j�=�o�0}qk�*���fv���?��� ��

��_C�Ni��Bj��X �O�:�Ik���Ů�g��I��J��o�kn#w['D��6T��TI���� o�%'VN��
b��k�#�e������G��ڹ�N;^���l{�ȍ�r���qUgݨ�f�R���	.&6��)|X�ژ�p�jT��t��`�4�h{��t��`��.0���|[�]L3���:�v�P�@��t�ͻ=fC�
�5�s#]�$�"�u~^�Ԅ�S�t���=�𤅈�aM��}��5�����Ӌ��ʶ,��dK4g�k�C7��������p�SKf"��Lò�d;�Pgۼ�X*X���m1] �Y�y}J*�-���@�:��)if���H��3��x���}�ߪg��K��5Σ���,�1m���QȄo��0��k6*��L�3�����݁��!K�Y	!��feE#��0z���F��!Ep]ƈ�r�0���B�� Na�� ��i�|O��F���k�mF��Fp�S�lU�\���g�Db+s1h��U�U}z��z��$cJ�?6DV�O惬�F���\�&���=��V�,Ǹԫ�Ԩ�~��x���0vB(w�A�D����t�%�bOmy�Ւ��w�h����y^���"���f������-��i��t��~�c�0ɫ�  ��q�����8I��픏�<�4��ط�� ��O���;+�?F���Qľn$k&����0��-�:�E%y���������-�P�6ax{��:���Zr��[��k3�d�@�'���{8�I� @q��u��)�SJ���.�Y�|Z7"�L�;�4�5;w�5ݍU)�ʏ�bc,�{'�1�&�5�P��ه#��m��|�8�33o� �y'�2�0�+d�<Sq��D��ȂF5�y�ObD�dű ��]�FRY{\�º�w"+ 5n�'��&� ˎ�сWj9��� �w�#v%�ۼ3l��
��m}�_�r��lά�⯦�`[;�����ː�eKj�LvY���&7����<KňOo(�SS]I����+��#���s;r�^��B?�H���0���{�HG$�0����tho��&s���l$SEV�+�ks��[����p1��M�:��Typ��$�zJ��.�LB��a۶��'�i��$�n FaQ���~2J�Ncg��+�}S����,������ڱ��
t+K��*��Q2�)�^���!�p�}��e[���UM�?-�`���P=#�1^��#*Aˡ�g�D�'�2�:g�`buS���O�X�#EX��6�;���m�����]���!�|Y6qUc�V�P���g�#֙,Ĉ�������JFlJ4���q��-�d�f�C+�9�Rp���S,z	��g$nZ$ .r�0_��a.��bS�M�������nc�}v�;��Ƭ��ߴ��Pois_f��Q ���_��3Ў�*9G����%:C� B�L��Re��L�&��T1�8YDy�����
UÞ�_�������d��V���L~�T�O0� A��=�o�BoZl�¶�"�	_��(U.I��T�9�i����쒁�afQ��<"i�pW�X��F�?w�O�~�=o��u���B�����%?IF����VH�pJO�-�o΃��cQ[(���'�	����9=Z��HԶ��|�����:�nF��^�ۛ�r��:PmS�e����!�׌�L�k�ͳP3Ž�;A�`D%S)[X��|�7�,�W�qn�B+�T3JVR�,���%ZQ4�x�s�H���� ,��=s�y�\�:�YP���`l9��˜�&�/h�l�n�l� ����n����~^���N��?d�1|0� �
9۟�k%չ�z�)�
��Wtq7��ş��ަv�c�*`��U��LY�=����9S�ʞ��Xs��M&䳉���E�Ӂ0�::^4�!5h�Qw��W��i�1��SJ�%�1������݀�{.m !륌�b	��ƴ�4��h�|h_���\R:U0�ˇ����{ޙw�`��*�~u̙=bC�[����e�^Ǧ�Q8�iT�bA[��ϭ���:S�fU���L�K�0Pb�`v��a�1[<w�������k����.��)�d���}T[5����j�u���mP�n�a��.��FS��ۜ
 ;p���!�0�FO�� R��G9�7���Wu~�P��>s
9�UQ'-�b�&��#ΪfE^.�� V~�Y�{��8Eaׁ!3a`�O�8�F),������E�0	���</\��l�i���g� ��N��d�ڙ�4��&;W��^6�d �p�m�<�_���2��	L��̫LرNi���?4Sp١��u����\��@�R�fa�ݬx�ڨL���#7���3������
��8@S�* �D�d<BJ7!�D��m����1d��C���aj(ge}�	c*`K�"P$��D��.�^������?Y_���mm�OJ��"p��Ze���7io� $f�)�
�j�ʉh��Q��vq�����ޠ� �޴�%���������;��t�k���#�l)��	|�sj��c���Ya�8By�������%�z�!HH��Σ��$l�٤,iZ��Xi�V�W����@h���<j�ܗ�e|3��-�Wdk�2��V@E���
�F(P���H_���ƫ�(c���{��a)"���+��
g��_5騴�)T����&!��|�F<�p�����V�yrZ�tqx��'F[jB��i<ڃbj�I��GWq�E��c�����:�,c�!bAM&GE|E�(@~==P�F]>n�^�z{=Ζ܍��M��X`s�&��iX���Ռѡv�*�6|��; ���ϙ�U8�pn�G���
HL[�⍌o�-�|�g�K0�k#Ew d5�G���� ������yRL����ϗf-�x�Ol��x�	��}�6����qsU.�˘��� �^�b�M�_������O��z�$\�+�(wF�u#�V"������;�Ƌ/�&':�2�͓)6�V�+e5)���3�H���<7t�^m_�c( � 1�ǻ�s�@OƘ�~~�d�a�ωTQ� ����i<��%��>��~�#�U�I��w�zl�kv�O��p\��Q��qY�m�"�}4���~�@c�=�S"4xD��6���_!p�	�z�����<����]�8׾�6��XWa�A�~���~��8��MҨ���G<3>!�� �����h�Ã�[�C�����YT�rQ띉����f�_Y�%g.R'C?r�
+X�T%a��n��e���r��{/�L�4ހ�<�%��O@K���>)�#�1�7�9>E�%X�7�bVB,�"3�2EmP��n�;�~\����l��!sׂ������,�.��mM�,>�yP��v����պ�GNÌEc%�ಽo�I��^�;���t8w.Q2�Y;)�X#_t6sE���>J����@R��'`H�QBq��<{�U�1�|���A��-3�i�n��_l�9˻�64 �=�С���[��H�fW$<��l[I��
� c���8Ҕ�&6�Q��!��;r�Bb�q�=�+�9�+\$9!���x��p���n���c������@m�l7��C&�,�͈��B.V�}�B��q�22P���6MEHD�ɑ�3��"�	��+�BN$���ʾ��o8��f/ʯ�
�\zj?Ғ���2�i9㖖��M�I1T�v�w�HY�?냯�����{͂�i��]?qI��p���V�?F����7�K��h�Ʃ�avPc�p8m.^��u
�a�����?�H��;�%�����}�PZx�)�\��G@����$�c!������.��s���c��{��m\�W���!A�O_��=u�wF2@́�O�PW�<�˟�e�O.�g���Րv�&N�P�ul���dݕ(1qo������x��2�sZ�b�5rra���az�c��^���"�y�����Nm��TĒ��ͮ����k%��H�L3O	�`���zU�5j���&�\�Rg�>����2x��o�M�(;�#(����YE�_��O�<�s~D&�:*q��f	�3��-h�l����p0�,|��Y��}�����!8E���h�ћk���
XR��E<|��jR}uv�	9@CL��?y���Z/�j��yǷe1=��(s��Ү��<l��!�P�"���b�u�J�r��x�~sߵ>E%����}��-����Ī l�]FO�no9v�K�S�h��&�#5��=�X�p�-������K14՛�= W �菟�Vҧ�,�� �Z�A���o�H��k08rk��Z���F���*�hd��ll�]I�����ب���DAw������U����2�hK�������'Y�)�L=>.۳�8�X���r��r���pZ���C��z�A��dG���C��ip����&Tze	�ɖc���:�@���'�A8,����sm68;9i���1�Agj@�g{u:X�7��k�:@Lj�4m���x>'Y��TL�8��� a�鮥DI��p��'`96Ƞ��K�s˦/!�����+�]���Eg�S�k���4�z���~59sR	���!H#�,����xع�_NF�5y�	Þ�ߡع��{��%N�Q�\����N#ҷԉ}�yh���R6���KE��^D�Af<g��ߑ��-�R�da"}��hzۅ⎍I��[WO�A���Aj�[��c�DgӉI�e���$+��u��کd%�vҚյ]V���Jq�����cɡ�C6^o`���>?%_H�sm$3�!�j����Ao�du�}�d�
T��+UH>���{7�$ �KV�W�J"m�}��M���~7J�"5��&M�����w�OiETG���8s��R7�G ���,}�5��>��!}��f1��f&��ȹ�h��o9�Tl����y'H��$З��	6:{7�������wYc������~�8���ǻT5,S?�w��z�Ӏ�a�ߏt!��ٽ�{�������)�Pٴ��U���[H�(��`r��֯��5����y�k|��q!�=�URY˕�v\���􏚬B1��N��!.���	�̀�8s��C������jfV���=��p]lVl�Xַʎ(DƗ,J|���m\�3Ii��[8��I��-/�n������ob���^�#�>�GBJ#r�:J�;��0���;B�B�^/�ȱW����U�v����rU�Ѫ5�k�!1Q����tmBsԯ�U���=�S��H���Q)�ܞ���3!xl�N�d����&���ڎ�W���U�ˬx)`������{H^z�Xbӯ�QX@���Uk3
���Ӏ�C�yg��W2���d^?<_�� ���ZX�Q��Z�(�~�Ʊ[�0����ϑ���>�BrC�Ff����`�z�����	�{�����[���\��O���ݯo�v�D(-M�]�x�Aᘻ	+h���wy�2V�z��XI�� ���	��+�"����U�x	s<���=�d@�X�[��?l(�5�Op�o(8���B�oU����{�~,T���a"���g�����ї�#�|(��������ƶn���p l8B�\2��*�̡t[��gnpmQ��c���8Sc��țU�lorf�Y�6��A:����,���/��ޏ��pD�Q�����xA�U��3�����=��lX��r����"Y�.>�4e�S��{k�������^����"����\�����UBj��h�������)�~�t���q%��3	���+Kk��>�ņ[�2�����ܓZt���M*9�W�;Q��k'��<�l�9&i7�kY����ĤTt�-�}����V9D���#���4(��c>����L���C��1f���cUf=S�Dpu�3�⁚��Y�dW���<��jU$�����>�������luε(ǚ�uÓ�e����r��FLlt�����7E�iY��7ܾE�G�VI�Y�CM֋���!�Q��a96Z-��c�8�:�9�,r!��*N�m{ �&�`̀�ex�ǘ%�N70+%��/��e|[�j+�'@��#����5_�;���m;��Ҕ��.��������3�bڑ��B����_r�0�����noO��?��"��	R�(D��)*��� �@|���_j�2~�o7t} U�nf�O����K�P:��@Q�Э�B�~Q6�,���W:΃Ǟ�o�|�٧��6��%�c1k���7�zΣ�\N
=�v�ˋh�]��8��_`߯8�l�����v�V�"�^�M�@0���G�1^<�<��gw�������*E[�K��^#/|��5}�W��uq'~�C�ߘF�3��E�.g����(���UFq���ט��tTC������$���<|0&^�}��Ng��C]�2̤�������?-����	��X�~�o����^ݕ�7������	2�&޾2K>s�'n��.Q#0�$�$��n^���©�ɀ�r�S���PƓ�qtո[qX���-E�~L�71�>�{;_�_`4'�z�-�������3اfk�޲���w"6���[ ���I؉��� �~�����6�9m���m���	���c	s16<�L��g��g�߷�u��O�y�4��}r\7!>kOa���<g[�����ORQ�	��u�����ݚ8�V�eSKl=Hf�T�`j�LDi��~�����hawE�S`^#��̟�
�S&w5�&Sc��`0�����$*Ѵ˕��l̠�ݘ^��DI������Jh�a�m���,D�W޷��]P��.��q���^��O�jz&�	:R��W�V}��g� �ؘ�*�s��$��K��rпuL�W7&A9̯4�G�uN�0/�XUm\���!��U�Sk�N�> �*�����䚂n���r�c,&�"��
�L���={y&�J"/���Ƒ;�&$���+/z��M�A��+�M�ٿ��X�ze���*�l=t��~���1���"�e#u�"Ӯ+/�0Oa;
 ��ܴ��H,60�T�h�`!���$^0�&��Nc_���o�ٱ
P��6W�(��?)�[�!̎"^�T{����GR��>���I<�#ʁ��9G�o�Ɨ�b�TJ�[i�2�8�O	�%�几5p��0-'�E��ze���z@p�_��nX��8O�X�*Lu��T}_�{�aQ�V���6��P���MToށ��a���j_ao�����1{�v�b݃�4�{��V$��v޽o��l|�=�����	=�8L�%�ze��ҡ#�K&�w���2�
y��w�t�?#04Y	9]�w�ؓ�>���|�.�����:1�)9ܺ~������O��[�R�ߑh�N�Rs%��)"+��̗y&7����:�UA���R8b��5Z�Z2�x��h���ၒȘ���P�G��Հ+r�C�4:L�T����L@~���Ǔl뾯������gûm����C^Y δ9���:��e������+�;Aa�\py�7V�yJV#Fc�����{,s��1�z�F�Ws����X���GBXg��7�:�_���ݾwU���b����"s}����zd����3�����v��8s�h����|��"	�$��z�fAa��n�m�4�j�m�H�^�jΦL�Pa(�ޚ9��n�Uw=��Zǽ/�[1[Jmj�CUI��Z���QIZ�,��a\�?u����������}߃�5H8�@�{�:�X�"w3p`�[�#%�v�����`�aֿ8��#jz�g˫ъoJX��P�9}�|abyw�qe@�dH}=�E~��g�t��?�~�M#Ҍ0������ ?�������	ɚ���j�Ka�M�Z����J�M�Y��.~�燯Y��6�n�Dz_�a���$}�(W	 �1S��͇�,.ӻ�1��BU���ɗ|�P��x���6d��,bb��A6�K+�,x��p�Jv/[�sݦ�0�|�ױ�_��e��(��et�p�
�J,�B����̒'&ƌ�ثo���=�e�w����H���U	���"�pi�Q �I�W7��
��Ǒmtp�+�Èz2�6թ0 0z��GP�S��\F�3�3-.�z�x���(<��+l�˧9���F��Un��R����:��
O�/t��Yg��,�. ]�!w��sT�h#�����(��A�f�urd����􄻧iј
��0H�*
����w��}��C����j=�3���?��@I{KX��v\���,���h|�9������K�9�\Ց\=�<2�{+��&cN�,,uL;q���� �U[���t4 cp"�[�~"S0␬ސ�㐬�h��8o�ꨦ��R-{h�9����x���N����������F*�2��H�����.�*�z�ی�`�
���%!b���Wh;<t����!�f�SA�Ƴ0�r@O؅���K 7�(���>�X��K��rm*p�̱�_��	��dWC��������"��K<m�yU���j�� K���G��/�?��&�PO$��}0�v
�~�ă���?�tpM=n�;߆�O�%��]"��$T���o� =�|��q��i���G��0Z�h�v��Ӭ���Sa<���8�Z<|��8�;a�#<&0jZ���&�]�t'�p��*)��������͈a`�C�_���XU��Y�S��o��?�nc�V^n���!��j��HQ��,!��E�ɹm��M'n{��<�E�\�mb��:*���D�=��b�U��Dm�Ŗ���a�����C�F���B9�.���r>ՠ)�+1#�<���e$��Z�+ɞ�5IkW쎁�d�C�j�z�{@ Q�\�ʇ�	`����(�+֔�[-�q����7���MoЀ@k�x��a�瓤Z�ܵÏ�<<?N
o_�=mh�:�Xo��:+����=p�����Қ�H����ms>� '���5c(�7�߽QY�xQS`6����l��8����t˗?+�j�6ĥ��p�b��D�����21�G?�mч����fUȲ.�<��<�:��ټ��N\�' -��wt�Ԋ#ٛj��Q���Vᶰ\;��� 8�/Ba-�>ָ�H���A��?`[ |�P̃�S/gp �%?�V�����KN':�ˬ�㑥'����'�<cf��2�^y��.\��Yr7��Se��TAUKn@�-Zvzi�V��S�Lv��-���/|���HNz����0��v�|Y��-�t��k��˙���l�����Z�>���~��t��H��TH� KIӇ(��|� |e�`yJ߷Y��� ���iɶ�����8J琷���$�]8�/	s�?�E]��VY��Gt��T�敯�a�X��%j�C�ߓפ�K�\�G�#b�ڒn�q|X�B:�9Ei��9��wng/8fd��w5�����x�5r2٩7�xѽȏ��ob3I/���V��J�u0ҋ7��|�F�����:��[V�;�����S6�C�c�čd��$���l�v-(2��1�����CᰐC����+�Ņp,X��e��)y)������$�V'e��Wn0HV���]�Y�j,!�'y8ȩ��-����}ٟ>�����-�wX��5G�觐`�65�|v�!I��tIΥm@r���ۺ���Ѕն��{�:�6<��hB?H�K9��gy@��Z��-DB�V�e��4�~�У��5���M�Ot�K��u���OD��E4���Ā�n?������h��b�K�Hno��P������u�3i(^�H{�R�cU�V(qۭ��r�$���<�̍�3 X#��A�rAq#�Q���w��џ�q$E�)4V�j���Yf|q9�Gv5�N5����:�Cm+�rd�uQM�9����Q��4U�Ԗ?���h�m�˞q���٦}+�i#�,KhY�������KL5ēB���d��*ݪy�@$k�Ggc���a�>�6;��:.w7�Ob���l9�_���X�D#Ș0��ẊB��#v����z��J������t��P�=����̂<y|)�4�f���}�!&Q�F�ܤ�a��'��" �͟�f��V��;�ɜjLU(϶\=�&8���q��GE�K!�9"?���zV+G�n�dXv5����t�}�f>Mr�T��5
�@��Hr�T��=C�<	��v*َى�&���^�C��
�����Ɋ���v��o�w(:�����B9W��l�%A��d�(�m�� �Y9����'����~:��1���Ո�� NђH|�%±�������>ϥ�wҿ5�a����] gnHB�>>Y헋� ^q�o��5���Ɗڒv��������v�d�h]ؼ��߉���
�,�_��?rV�$�gy�����
>�fDn�K�tc+{���Y��L*o�q&����6����pD�������/)ܿ-����#����'>��F���B�����p��?a�������q{�?�5�u��*ܷ�r�S��yT@`�M���g��䜱��[ęBI�ʛ_�E��rүDl �?{�w-�����u��`��O�,�x�T;��9��1ly��;���YJFƊQ������(�o�M>�4�J"@2h�Jo��:���j���EgNFX��s��kZ?��x�Kv��'���h"9�g��k�_*��2�Z̃ 0vBdW	9��Ϛv��fM��u%zR��bg��u9.$TӞ�/����j*Ƃ�[^TX�t"o;��[TS$�t�p�1�Ӌ����FR�4y�g�q�B��d(׌L�f� ��Vs��j��	[��C�+U�y��hp������
��⾙�v���d?�-K��A_���^�����/Yɬ�]F�f� ]���=�F�˽
cZ����0��
�vז�{��a��`�������ۀ�<a�Am� x�lx*JDr�0�r��B'��-��{�9ٛ6�S�~K8�ā|�O,�L{z�� (���x�92�j�|L����'��dy���5u7����L��i�]Z�ʖ�4�����R�ѱ �M���͆�8�����ptZq\�8�ӈ���ݨ���)^��kڳ6���y�g0�T��KGg��ć񃍲C�i���������s�Z*���?�t���tۢ��aѤ�k�I�ݻlEf����]CƾF�1}2}��A����2xPv�NtU��N�9*��f��hIqۇ[5���]h�By z�X��M�٧=W���'��v�t�I��`�[ �V�5:�ח��+u�Zͅlh�I����~����,ypcfi������(#Hu�[{�>^������\*�eA�l�]�d=��o�j�e����ؓ���8�g+`@6U��V�oPK_bƩ�ze�<�L/�;K�%��8jw��0�w�xN�������y6�nH4jb�N�Xy+��yO5�Xn��2|Z_����EѴ����f�3��
�c%�:�Z@�mKǶ�xdZ� E˵]�Nj����N���U&)�P\�R���Dk�}a��e�cD��Zl-v�Z�����z��c��t&t��,�]�!"�Qq�h�$Z��.�p�^ٻ��<č���:fQ���,й�VQ�R������߄R�J�����K�k����<�У@�3���Q,�Q��Qj�v��P{��Tr��Pѭ"�핲TB[Y���'���>�(�iX�����g�	D�j��\7[y�Gg�ف9��4�/����j)�jc���̨5XC� �� ?)��:�b�٭ ����;��Nd�ѦT�9̔�z��dO~iҥ���=�Cx�2E���G���`d�SA� �Ѷ>bHߚ˟q�m�c���ܕ�C��O�h��𧃆�C�3�K-��ކ�:�ȯ7 �<�B���0�7��V� ���e���u�������m��gȭ�$,p�0�/�C	L��&���31fǣ�^���{�UcYO`�^�k�q��
�B� 1֬:�M��7���T͛�	rp�.�h� ��w�|�s^]�C�#[b,J?��S	#��8�
����!��d+=�I�[bU>ᓖX�
ڞ�>Uq��PŶ��-�ב��ɻ�e�	�	q�u��)Y&�g���B��F�}ևN\g)빦a"��$<�/i!����q����ҿ��Z�+�9L�E�� ���e|���zq��ګ�䕁G�NL�W�RE�����/�'8�V��Ǚ�
�F)0�eI@F����h��[�:CCwŚ?skA\%A����5�m����ڶ{M%=Af�c�'�X�IF;`���5��tiS'��^%:6�W���yH�3�U䞿_؆G�����7lz�qX��% �R��)HCUQ-��g��Ǉ+ 7���C�6B~",d��XH���T�w|^�(��>8�J���į��j��X*U�<#/m�-=���S�W���n�w������h&���E`�P����3Hn�vA�p����p��<�ӁۅD�%R��~u$�{�FtG��g.���>���"�����z�W}y<xѴ�me�*��0ޡ���S,	:��F0T�H��-���V*x�[Ac*�*>Dc��˛�TC�~�����-�k�s!���w�ۓ/R�,�l���T�8�^l��}�C[��-P`Rc�]i������K��szߨw"hZ�z�є�c��|��)/�L��)������ʛ,cձ�:v��)0�#
 �fO=���.Y��|X&�7���6�$J���9H��m��2���"苌�R�Ck���|�'���]R#	��@�/���>T�?��*��o|j�JR�/�4��H4�,����\J�Xj�/�C�&\1��>R�Y��،%���9�^0R;	�3��(WW�6�;uP��[i)�HƊ�Q��IT�v���g���W��g�K��<8��	�8���Jz���Ea�@�]��	�tށ�ĕI���QZ#Ɨ�%~�i�(�:���i�I�����B�L�Xk�\I{�t{����M8r��zo�ow�xi�`H:�D��y����P9xUO��P	��&�8�0�u��8'�\�b��c|�`U�iK��;�c�6��e�	�lF;�4i���s�����<-Y���3�=r�#��4���m`T�������qw�N�v�����g#����+)�],G����2}uӠ�
�g�.4��G��EFI;���V~���������!fW�|��v�j����Y����;�%�e%7n5���]����/�H�*+E�����%E�l�.��m����ѭa|���{�DV��w�Z���t���|2P��=Z�0�
�q���?�^�n<t�FG�]��ܰ��,��W��� �l�e�k��a�;2K���./��&^Z��gN�YB�I �h�GCf�5{bE���(U��M�o]�Y�(p�{��:C�O����>dF�����%��7���G��t�Z�����J��c����9�JoΦ��3}l4ǱR������ů�z�p�f�
S�mD:�y'���W�~ר����ݘ,R�Q9nf,��αZ���PS�c L�x68��v��&/j$��T�Jk-�����^TG?��Mw�rHN��U�-��)� �����%�K�CD�"��MR��3*b��Ƥ��f@�qo��-������_�����oJ��"ƗNHٮ�K]y���'$΋�gh/q!�fvl����,-��{��f�����w�,5S.��f0�l�Gx���*��*�@]`X4�Np��%�7q\�D+��v�V4y��+�.Z�܃���<�	��Ux n�G�j��� x���P���V=4�~/�@J�k�X���BF��/J/x���z�>���K��E�Ї�C)h[2��[�#,�)�G��/W�3���+c8SL٤7d`���C��V���J�l�]�+��~p��X�k�F|��S|��ΐM��w�d�KϮw���?����+�/x�i�D�����s�6&�p[��!�}8u��B�,`H`Z���R�H���&�v�j3w�� ��[ZNTL|�S�C�T��#"��%�Ǽ%'���A��I������i�=�8nw��%eZ�)�sG5l$js�E��V������[�%}�Ѵ8�XQ��W�K���a3Z�S��j n�r�Z
@��@)��!�8hŌ#��g��bFy��:�@���noX̘�#�����D�9���Q�k�H��
�'Z��Qp3� �~��0��V�����z6i�a�~��b�w~T�Q�Z�T���&�֜H��.I�R�7��TC@���R�goc��-s%�7a$�ʥ��
X�[/�������*�%Y�5��u:H�j�&I�l��Y�@�a
���H�w�׮v�w�2��d_F�xA�ŵ`"�562�W���o�5�Ls�>Ih~5���ޛ��h����'L�Q�r��,'8>���&�3�X�ci+,A�{��e��t?���#+[b^n'עAd��,��i�&n�{Vw�.D����EiL�:��92R�5rgC��N?%4e�'�Hs���~59�K��8���`e�Aѝ�̛/O{��Ő��E�y�[ۆ�v0�֭�wsq4gS�W�"�����`M.j|��넱+�Ia��A􉷥0�q�C�>Bu<���9uir��c̯��������v�]¤z�#�G�
+-i2P#FJ��?�&t�6O�+�Je��R�%YF�_����Smcβ�ZO�� �$&ċ/!�L�˕�A�5�:�[�/�IK+"(t��]6�+X7Ƿ�[8�J.6@�5�鐿�,tV]����<D[]�_/��­'������;'�{�C-'BUw-��3v�W�ڑ�zyz�x�� @�,����RO��L�y�TLXg�����I{,�q �C?$: c�J��fE��ƓQ��f����UX�&_4�=��@d�fJ�w��Ö���s'Uz��Dg��Ѱ��M��]����X�St�$����Gq��g�6��s�y2Գ[�~a�={mKvp	a�\*�Zz	%�����=LԹkP�_-�5�>9a�*T�\����!�֭�n�F�Ԗ<5�~�Efsv�^>����f��ԇ�����@m�.V��P���QX @Y�-1xի��~?�q��I��Pp��ߓ�pN���N��� ��q7\��v���8L^xWE�R7�I�  o3j���\)�m�\	$��Z���0{K��}��S%�Kx�2�����ʐ�y�u��-:Y�l�J�k�."�Gt��c�i��K��4�%q���VEk����i-����)*)�k~�{77c{�VRӿ�j�v��F�u�����gԬ�Ǔ�@�+�RE����/���^�jz ;��U�����}G�?˂D�3�u��SJ�~��o��1�6���a��S索۹r�LpMP�+�Y�?�[���LQr����0?�,>L��9Rh�u�uuX�9�L��~V(���@E�I�9Nt�܃�y]��P����B=,��f��k\��6�f�3���z`u����j�X#���׶6�r�c^��`�P_>0� ���l�;����?*�7�ؼ�4v�+�ucgp�Dn�~5����%MzZ����k:5,�{��I�Cj�%6%mj���J���v��6H�s��,��{E��Qo��Ã���������VDU�q��+��d�g7j�6�/�3��fE0.�O���1EQ�)��P�|��EZOi�y%|ck�ʻO��}�Ss, W�*��<�'�܉D�����#������q��%9����pBw��Z�h�� 9�X���-ơ�f��A�o�b2)��Y��mS��7��:��4�dQ�h�~���5ͮ�����-���س`�dl����,��&Y��<�[���J_��ۣf��Ԅ8�o�@Ί)N4�hmn+'�0���[��#�!�EF��ESa+����Q
"�3�ĺ�	��OP����t=�|2�h�j��a�MⲎ�"���o/�"�H��WH!��龉#+Ȋ�O��D�v굥�Z{=�&4�[Oo[����"�Wr�eΈ���=&8F��5�'�ؐ]d'�e���.���GL�v�Q��8z��	��׸�gbzy��c"S��s�����7���V�:���	�+�"�Ӧi��Z���C��9�jw��"˼�d�΀4�ݐe@��e�R3r�N_�}���)��n�Av��{_
ܓ��~��b�X�u!%^"�'k��	�����>V�c�Bۨ��h����ں�C;��׷�w�������"����r�'���"wR�e[����]C� J�������z5=Q�s[%Q��`��϶i�h�B5�ktd�a�AK�-�S��Jg�y�L�\g����6��t��r�'VG*$J��� :��V�J;��<���A��	���T��G�,4�|��9�0�?�l���Q}uBI�.Ut%qJ�n���{�d���mG)�����R7�22Ե߈> b-�Ӝx�mKā�����w,��{��v����S$H�l~7T_�C�
Տ��Y'�<&�- �Xcu��0lσ`n��{��O�Ӥ�V��AC�xrFm_�rH��������WE�n���dy}��My��|
;��f��'Ve��;8���.T 	�b�~����89��Hsb�u~��\�r��T(��i}C^=~\h��<���u���)�K�]�Ed��տ�L*Q�VO�o�rU��;�9���uWA%�1�����d�xE�4x����B��I��[��d·�Љ��|-��m�d=&H�A4����K�&RY�G�Yu)Ve��:�B�!����-cy%r*D��\-,؝�icL�)�<d�9��J��� �͖�°ֶ��BO���D��йHkN���oL���"�K,����V�M�����I	�J�>ϒ8�;��WW|���Duj������tZ�5߸�6zZ &y�{�Ԇ�@t�",���C�5���ƴT�')�
0K�2fY��G� �����꿫�^�]K����['��J�%C~���m�}6/N�����R��a�n��x�qǦ|f��X4V�)�-��Q�6t�Yq�{
�b�Ax; %>x~�lc�z�j�5�ڑ�[�D�	�������{��_u��%�!`�A3�H�k���ߊ�G�����Oe֍@�6	������f�����k����=��R]�D���UB�f#ŕ�l���ƠPD-o�f5c�m���0�a,2 �\�[��C�π�C��.��n$�_HL'��2����9�n&t4�_�k��Fy�tYP��{1��k:I����������ɯ�i�i�F'< ������aq�,$~��ϟ�[��Y2�A�lx��r�S��iq���ս�C]w�6@�5﬽�N����D\�K��+~�58J�� \-�����fb@�U�[uū��{�PRI�M6��lpKc�6P��"$DCV;�9�H`�jӼ����������X�^Kn����p�G�(W�f�h�[م��� �v���=ǥc��9Deg���Ο	ZZ����@|�#�;���l�����z�ݪE�o���&����w!�|�ư�#ؓ�S��K��1OO��RG�L�Z���Ƀlzbk�$�F6�6>�+Ь+���hYI\|t*�%�S��α�(�-<����v�D�]��R���RF�%�I����r�?G[�m	��Y4��U
9G��F`N"T	��� �;�k�TW��G��t|����_���_EJ逛'͂�e@�ҭ|�V-+�҂;�@�1 p.:�$J���B/����y�z|^��D����Q����!�^�PU��HQD�?O�v)Ɖ�W��C�)|1��[-����wY�1�6^���CߘR���w����	i�����M9z"�L� �~������qzu�sƄ��a��q�Y���e��g� �ߘ"���-������mU�#qqE(�uko���ϩ\�)����ó����z�0��}��W�F|cLt����2�<��"��]�-q�,@�{h�Tϙ(���A��u�� 
z׷�^�2���<*Q���/�S?�a�E��"�~xF�	�ݪys��H����eDu���#���R�@�NÛE��e�;RG���F�M���Q���Q;C������=Q4���k�5K�?�c��AJ��P�~W�z�S�Y�ݼBswfM�&K���=)яX�.7��H�WxsWz�{���� 0M���Q����VX/�!7��՘Ѯ��k*���}s��kw���aF[�	�ɚR0�C�h�w(>@?�#U<�[\�U����(4�f��>/jpU�����4i��p��;a�J[�.���[�)�z-QTΥ�J2J�G�%��1��R�~�.����V����R��۪3	�f�zM��5v*g�����736W)��F6��S��C-O;V���}��
[���������&d�UU/�[������ӌҍI}p������Y"�t�������. �`J���H`������u���^>{n�GbH�	��H;�˸��
}]Z�1��.pk�S��9��k������E�螾��k���G "�[^Ŕ��ыܯݲ�-O����S�l�2r��rL�nZ$�7�3��Ȏ��3�Baf�<w��3aXk�?o�tz�x�����6�Jz��.��Ү�l�.���b� :(Ck�j�9���.���,�=�7��m�+�  �7*�<'^�����W�jB���ﮊ�7�n�G`��]��Ԑv��HG�{K-YS���F^�*�5�()�B
�Ҡ��
�1C��������`�5�3���"����W��E'�4���W��h��,�D:����Y���~�c��ܽ�L"��5�[&�E���Hr�/�Yt�Z���B�����Ł�p�5�2�̔h��@V��A�a$�+D�m4v��Q�k�CTp(��]pvY=����Lo��/O{��d-���vV'W>~5��'����-�}�ąp1���;2m�V_g�;�ޕH�y�˘.,ů���e9t��8Fz�~��&���W�Z
�A��0{~ǡ�� V�=�'�7��B�i�_&H��X�3,���ZEvb�
3I'�Lr8R�0Jj��h��kA�d�8K<΋���}	;Yu}ُ�+�候��!�r|�6������փ+��^��/�d�Hk�� ���IJ�m��+H���2���U���|�1���[Y��&� ���(�v�=&7i��ٙ�>h}�������0���p�JH}��<��p��������u��"���K���,�t�*X�1���-8־�үw�qY����� *|� �����19^�$�Ru��<,2��1��)�mK�
�ܱO�;z��~�'�����6i�`����C1L]S)$�ѳ�Y-`i��\f��
"Ȼ=�d��63�kxT��i��]�wb�׏�Ӻ������]T��)�	��p���o�Bގ%� q�^p�	�X���(��[�HI!��xC�˗䖮A�M�oO�?� ��dd\����e/5]B�?U`+7Pѡ!����/���A]����u��z��
c!Ii7��/PNk�=��M�ɔ��t�/�3�7�2�j���Y�p?*�#,XR�2�$#am|mNJA�v���e���U:T���Ib��R	�T���?Q������r9�aT��T��i�A}�	f#�S�G_}PQ��0[�%��[%w��&0�z���2�M�{�K��0�Rd�#��Z�v~�̠g0c��m�38+�_R`�ь����ӑ�/<�'K!zƮԬ�� 8ۂ�60_��8J��FI�3�2�ח�~��.��Xal�$�F�P�i��g3�c�	��ȷ8��݃�Z'J���T��\����K甫���'֫=��#���k��auհgH���5�ٺ��$2e��<�C����.+���Kmr�ߎ�I(�As��(�(�'N4M�󝺰��Wa��_�r0�{_n��A�^�y��%��P7֩$a^�&�ݣڤ'
0үc<�z�ڢ������3�>�V���a�.B?����܊��й¯�?�Ų�+1�{��F����f��
��o��2fD�tĀ�����t'N6$.��J�4an�c/�⨟ʎ�S+���-�QT�H��F�;���}�EJ,�
���e)t�)�
0����]1�hx~wڮca{�L۪!m\�N]b���}s�4;G�w+ Mc�Ge좕��5`I�����!,��h�3&"z�(�#��S��ӰgR��|6��8'��M�˚����`z�ʦ!� P��J�/����
�]+�{%d��GL��'Oc��g8�b��'�ťXլ���s��0��P 﫧�ܰ �3�OKf�}�5�7z���mpOy�Vk�L��e����t �f���Uoh$ƈ��I���;їA$�xt��$݁��KQ�I���o!�������u82{�8f%*����>�U�3L�y�k�zm(S"� i%��V�]�x�����l�_b����^�wuo���˼!��:�	�7�q뎈]�L��}N� �M�N5��� �t���C�5Cm�(�9k"IZqj^�U�[�L9jɀ�m@Tf>؝_�s=B�o�Wt��^+ �{P]0�R���(�gӗ�G�}���#��V�w��,zm��	D�k��u�]��ܸW��E
L�n�	n�>� 3,a����0?�;��G|�_?�uc�<�)Z,��~�F��4� �'K��mR��v�!O���C�d��p�&�;�єܕq��o�z��f؛��30P�n��rx6�p��\Xc�?j���X�S�܊�j�$L�{hj�V-Ѝ9����0��sw�A���1X1�m=�y�G�#o- �.��]*h��9\d�����
�;M	P�&@�������T�~@ɰ^8Og��ڔfh�lk$����_R%���T�z�hC�R}x��6�"�Dqa[�-���e(��o:\:�+����%���f�+7�ttS*Z�����h�ǠX�>`(P����ÑH@C���R^98a�=�|`��̴���1�#ڗ#`f��}���A���h�dLR�����_J��i*�,��b���g@6Y��G ґ��Z���!vf~��҇�Ӯ��#߲.K��D{\��n+�ul�7xڣ�x�AS~R�a�F!e�+�jK��Ubk�Ζ���ss��t~��8��t�%��[�����x�zv�>"g�OӜ�u����j� ͨ\��$7����uTW=+���B�a����k�R��:�xm����9|po�:jS�R92�P67����BM/�x=�$Qv��6�pO�r}�	yE���P+�g:Wl�z�w\��L�`&ˉ�-�q5?����uεf����je��h.OցKZ�Du���G����^4�ܓ 4���N]�