��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW������r�c�v�e�������Q�6�E��>��P�&�?6(���I�٠b�A���V��0f���;���i�c��\� ޣY>H�E��3Բ�W�S��Ÿb	 ���5��G��r>��T�CF*�{D�̟�[�$xi��:Ԗ u׳����.x�7���*"�k��c���a�-%}�y(>�hž���4���^�X#�f*g"�g�Uu��7Sh�	� �ƌ��!����盛"��q�#R�eTX����'
�,�
�?H��_���տç=y� ������Qt��x��.o>��K���=�&�H9"}�`�ouR����������DK%���I�.b4��e#�0krՑ�����Pi.�n*���-���^�q��A��x��V��u���_��0�߀��W�e�<o��;��罇m"�9�2ē�����/�gl��"��y�^��f�2gI�6�ﶀ|�u�isWnK,����^�
>�ν��&/˥q��S�p�_X;tD��+��ӹ�Э�rd�l[�7)a��T<�S2��R���/p�	�s��[���n��F;^�S�[�%x�_��rPTj�xJ��6�d�*@�`�eq����,_8FDuDjj�#4�'�,8�y��f����<�0�W�,�;��$R8+l_�$ �L�)Bb��*�H�{g/�	��}����Kq?�1�;�@#x�����p��u��"�4�o�+
� ����c��}������h��HDć
��k$�iJP�g�k�.& {Fi�֜�p����W�h;�"9���&�7��y
΁�xx&g?�Z7����A��P�h�vq$,e���,`�f	1���etf�����H�� &'*[�0���f�d�H�O�"�OS4�,�~Ig�-�J@;0���i�k*e{7�>����2��:T�3׏�d�lV�C��1���f�B䀎�%���<(�]û_J:E�#�� ���`.��bʘ��ι=�d>oJ<������Ԫ�h���!�X��Hei�Ez� Q���R�S��2R���m;Z9���������?%�>&�N.ET�'F$.cv�6��'��>gn��]Vr9h�1�rv:�?xM���'z��.K��ć�×��M�I|�v���)N,��hL��a�m���<6��\�~z��֑ h�2k��u�H��3Dӳ�E�r~q��V��W�CY[;פ?cr!���"	GҞ^A'��,ɖ3_��7�$����\>�D�s��AW�ɏcz�F=��e.��P���`�Ll�`��ٱ_Tg�׭`�k�l���է4��-H���Gɏ|}�O����>�����g�_�Uڝ)��h�{|��/��:D��/B���?y'6�wu�H!om�[rռ��_p��q�g�;�2�(̅���l�0�$�����ɳ���|���
��z_C�LȌ�N��増�J��#8���]v_�Jdz8s�����g*�Q������J2k�84��T��~Y'T''�M���z0��+�o����1��*�W�=��oXD/���;A�����0zup�?�n�=*�$����eSb�Ta����{�/|�e[ɞ�S��Ӡ�y���uA�LsݟUF�V�z��rٖ4��I���E\U�>�O^`�"s���zjpwk٦��O�g��AA�U��j��K$-	6fh���9��iO'�� G����A���W8�"R��t5q�3}|�E�ׅ�g�D���]��֭�#��$p�}�'�pqJ���c�]�5�wI-x�vIi�̏���u�6�w��OӰ��P6[^?��]N�\�p�
̃{����HÄO_��\i��f�w_��g2(#�a�l�!��a`�U2z��Y��ߢȵ�;�������d��$`2S-��������U�n(p��N��=��5W���3�:2f�A|R.:sN)26^iXv�]ܣ����c��b�eն�U�*ywy�����P9M�7E"�'�S����%l�~b;ݴ���o��Q��{��#&�<�r�W�h��XZ�Fs�r����Ƅ��ȹ���~"ݯ%;�I�j��ؾ�� �}�wN6�$������OB4Z�S��gQ�@ 
�<�u��O�q$��&���ϔ�f�7���̓��0šW)��R�7�����oH$G���V̰-S��n�=f8��;>eY+�.oZ�&��c����Vc*��c{y�8A'�L)�j̈��ǏZ�U颁��&4?f�V��Y����ZH���!R�>�3`�W!w,�U/�~����C�z��)���Ƨ��[g��e/Kv���2s���h@�΃���[k*����{�c�5[�K��3w�?�+��&T��멎s����D�Ca�����+���XjU�!�yP����Ua��?��O�U.�꿥H�Ǒ3X�_1v�`(c^�+9�V�\D��V~ם.���L���Z �Q_?�.,Q!!�3�t�H��Cm5�k)�3�ԃ�ѾE�ִ[��/`��5F����P:$�L��p��&���ڈ�c�(���r�)���G}gc9MY�0�R�um>��u�js��O�C,!�5�Jr��(���mi^-GO'.�S|�.уB��i��,��<������iU��f�7�,tC�1&ܙH5���BI���T�|p��%}ұ/~w��#�	b��1��`^ڂ����6�5*�-�-,OS��@y4�E ���zb��#�JC�����J��H��˫m"'���o#������Þ�^ۚ���s�J���':�P7� �>g��-�/��T;��>�I���*�s�p��Y[*�;��5�X���ϝKk��o�.ڏe.CH²��׮.Z8����CBٜA�k5=T��8�"�S����߭��n�ڛ��k�q�c�tbف���߈��<����M7^�P(�V�n��;�2�@��rS��8#Dip�b�Q�ל$���(�4>��)Qr"Of��].� nT;�����3}����4��HŸ׶Vr<evb�Lh�8H2�}�%�O(�F����-��0�5��r��=(�p�I��b�,������6��P�{���F�ȏPq�U�h�_�*v.��9�	��.竊;t����Fs�6[��k����z(�=w%)���F�:���%G���x��0�۶=?�xk�D��>13���C���.��"���Zn�
s���*�*<xy�ۇ|��No1���!��J%1Hy��8/��˽-s/7�s�y��c�ۉ;�($��E*q� v�U��&��
���>X�^�0Y��]�͘��xFPg�0 ���\:VY d-=�r�8�O�b7l3�꺽��DO^�O��۹�5m���5�"�<<����8��7�#�!�+�F��랐��u{H��&�RN{�{���@# ���ΐ|i�Ҹ�,a�
�F|o�B�R�'����,|Y��2 ���q���v:��v�`�.Rzۡ�;a���W?G��L���R]����BE$t��*3�6�3�c
GU����%E;��Ě��XJ�1u0�|>)��q��%���|
�^��c�a:�����q���V���C(J2�ǂ�����{%�ڢ(����~%�g��g����l�>8QT���P���z��l���������Y��K�d�uC�UɉF4(/,�*Q��9 ��~�0Zƚ? Ur辊g����|[[N��h���\�5D�� 9�T��S��mF���9�W���&���{��)���\E�wҕ+K�GT��`[/5�c�\2j|�_q���:Mz�l9��~��`^��]m����.<��H1;���C�-e�S�19��){���X��k���^#�힕�<�&��=L5j:�5��,'_�R�Z3�潸��Hr��
���WO�)1���f�%A� cD�}ȿ��/�ӫ����*ƭh1���`���x��Z#F�|y���Jb&ф���ݞ��Rmw~���@�>U�c�^�&ytF�꽣��c�]ӷ}7=�6����O�q<)sVU/�,uS
	k��罔l
 ʐ�����0T�.�n!�Y��_�ɦ��;$�-��y�EG�uOLФƻ�+׊�w��X��S��@"{hOy�cf��y��f��vD�e������kOJ�D��Ǌ
쩠�'rV��(�J�#�ֳ���-��w�Vd>��:J�Ө� �:I��PS=�]��\*�;���
[��}ݍٓ��q���y��j/&{}w� �G��$Cz���d�~��>�M:~�2z��4���|�HsU�@>��o�^��\�ҬTQEC�d�� �~)r��M�G4I��˷�~;Ȕ!S
���L��@�@*�a�mԳ�A���A�N�p0�ͼ�7{����N�	��z��K��bZv]��y�b�8y���~��q��Zʠ�>��K��vE���>C}�ZL�Ge^����X�oI�W~����Xw���3u���}Ν�z+&'
�?\^\+�ɓ���r� �aǙ�kM.s=��CGB�7�����i��-��>�T�_Cm����0z��\Ns��p�5��a��?Ȳ]D����Q�"z���䦔�)�rsuDH�By����K� ���\�2��7�Ѯ�J6��zJ��?��@D�t�g(Ϋa�z��%z�`���["��_�ʇ��Ǘ/7���[�6���R�;����౒QK���r �B�� ����-�I�Ea{#
�M�t�&7�Nr3�����l�N .��6����3�n��gn�_
�4�����`,��b�@woʏ�.�Ǡ��r?���*e�2��j4���+���1_j�=p����I([]�e}�z�U�i��Wձ2VEtL����~���wTdez��=&�n��/M��'�zr��C��^K7<��8E<�\s��[|�3(>rU�I0�����}�!U$ߪy�	voF��G쐢�ǔD`�a��v�0!�.J��¤{�'_\�����3����^2�ӹ�fHi�w�&�Ћm8�M�e�.�㗮�
'��;曣E�b d�0�Rk�>��kM���B+�Mx��6��P6����\<�������h����4�z���o��q9��#,��e"��v|�d.����d��KF&�Q1�N�u����K�@��I869�hx�hu[/Ov�a�TAB��t�O.b�R1(7�A`	�$�fJ�.���mȠj��!1۸+b�ǁ��/KG��VY�=go���Νߒ�"l~�X$���V�XTd,��I0�x�t/���J�%�j�`$U�*�F�o6?���L���~����l���$�3�6 �Q����r��~|:�ۃ�*�p`�L�zU�^'{* ���!�n]����66?����+Y�7��P�s�cWf����Ya(���Ç�>��A/�Ԣh����+N�/�O���|+�w��pQ���и���J���?�<���9��p"w�H�hM���-x;����(%��9L�t���C*�*IݑKt���S4jz	���NKj�����U+-��n2�	i��.ye�H���D�sJ��+Z�yQ�S����ep�'��m�7�a���0�s�e�|�*��}�O�a��/��!�m���[�m��ה������N,5JO0�azAt�%�k�1;)�v��ٳl��>!aܫ6sM�J$ߥ��n�J�פQ�b�jl�_��3�Ojۼ$��J���<� X�.�O���,��}{h�y,sC/Ubp�;G3���ܽ���joP�V�)d�F��K�ڕp�i#G����t ��d���aޗ�Y8}㫯����|ugYym���<L�����_��)�/�t��G޹$���X��j�y[�CMK�f�	�6�rg��_��̙�>���1<#���q=+�s�hM���^�s�����q�IXcO�C�{g�rv�)�h�fc�x�����<h�"��܏4Nn��"aL;�>�)�;dqp�`�O%�g�n��:n1E�V�L�5W�%��ю"� ��S��H�j��x'[��N鯋��;{�~b0	��4��4*��u����!�}(��X��
���{×��xp��y7�_��ԅF1@�P�r���j�>/��z� �K2!*�<$Z]f�HT���<��HF�ou�x���sߩ��@���K��X� H��.�y��*|���������ӝ<�����i����#�C��z*���P�=�_�od{ѵ�J�1��4�-�%QCX�e�Ӻ�����NH
�~dk�kb��KV:Eɿg<��ҁ,iY��Rؚ���^���藊i����ތ��Nc3/~��`<b�Pv�;B��Ʌ��2�5{K��߬�޸��W��R��9[������ۖa�����:=�c�_�E��ط�N�k��q��%~�s��l)�����;S$pQ!��:6,/�6V�	UФn�o��h~�ͣ+�A��Q��0Kx��s���s)�s�$J�5���q&"��|q?	)
���m��-�H��;�����:��t�z�E�R�Y�w�׬�<�v��<�~5rS�mg�U��f�v5j{B��%@���X����)�T�l��ΰ��&�"	�h��<®^pP!���?u��\����
� 3�����R3��4�3��&s�ڧ
~h$�Vz�)G 6��-� o͇���L���KDA�l���"��0&"���8�*Fکd�U]m��*�� ��E�&FȒ�v@A
�Ϣ*�]����2����$�3���JB�r�������Q�.'�Xd��4�+�Ϣ@��hg<��\��Nv����K����d�RyR��.��*V�Oh0�J��ے��&)I��r�����f[X#-�� �.�i7���R� ����c���H�!��=�`s�����]4�q�J'?N����"�_�T`�UEH��n,6܉�A�]_�u���p�OͰ�|J֠�,T�9�b[��bM;W���^0$��^xL��p���WH*�D=�>�ڥB�:���\�h��
M*���K�����%��{Q��Մ6-��o�L���L����:DQ���⼆��ޯ��ʶ23>�}c�~�L�g�N"��("Z$UAɹ�NN�5���E�S�)ӣL������p/=v�u�b���A���_����bcx��;�aߝd%�3�m8�>�2z������6�cg�-xr�������.� ��D�S&�~�q�[�}�`�ڔ�	�Y��1/c�T��O2U��%���.!(�4�
i���!��)��Ni,ޜ��y�fn^- Aנ� �������K�^�O/ڷ*�r݂�<�!��hzdoti8*����
G���Wq�iO���N@�`OP�`wӱ��"Rn�B�N��(�?uqer�u.�������ȫ�]�񽖦o�-2L�� /�m�͑r.ű�D]���
�Wr����2~#�n�="�0\�:+)���Γ�_7Ý�tst��NyiqA�&Z��]y���>\����;~���"F7j1U�,������Ea=��1��|���o�;H/�T��ОF6f2��m��ݽ?��!�	�a�T�X�k\�V��b����\��1z7y�7�������v��d@ԙ	��
j/!��sF�Mn6��h����ŰB�D�|�D�{���ee ��Z�.�/0.w�Ti<�+膱>?��t�o��#Q~MI-Ha3�(^�;-gQv��U�U�MSL|)ϭ%|�k�麮Sf��X=�5\����5�nU�������\܋A�yR������U�h���x<-�N�F�݇���̬Z;�6w����bv�J��Ϋ�֜!BXH��lÉ���o������|Uޅ�;��p�LdP1�>�
��?=4��k�ۀD�P��f~��9L<Hm�PK�"�����R�w佰:�f܍O��&�W����I����c):or�ܢ��F,���t)�aػ��Z>��i�L��d��-ښ��s�'��MX�8�8&���7���P�4�H찪��W��Y��:��/W�*�&����߱�jߣ�..�	՝b61���z��jع5:�	��+7.�|��veV�x��Q�7����,�=���ǝ~����WN��M���fy ̄�2�"a�,!�fPr��]^������j��O�/֋�!N�?�~�����܀�;�]K���e��E}8Km���9��|ķR���ˡ]X�Fa�{C���4�ѭ�ǰgL����rTb������6�?F7<���:����cx%�3�A�&����i��)�5^�u���Tq�W"osH�������Fҷ�	yx���~qM��r�Z"ʐ�;���.5f�F@Gnx�C���q��Ζ;�	�e���Gr�a��i�^ˆ$ڿ����t��ɱ��WN%}>�Ɗ*���w9X���iN�4Z/�5�II�:�.�Y\r�� ���}^/�D��5�55)lv����w�F��
�@Z�C��򌆴Į�
�����KQ��������To�i�d_��}ݴc���Mh3}�XvWAK�i�8a�D��S��u�P���D>0p	͘�h��� �'�d���|4��$�g= �!(��kkZC�}�z��������];�Pz-���~$����[B���Ic/+VD����,�^K#4`�j]%5U�'��G�Г>U�n%���Oj��� �����,�nK�������z����O"K�hN#C.0�����R�ϛ*.w��ۍ�-�����l��d	A����]��	�U]��(�W�еV��!��K�
N���H��)k8�*]�Ƹ8�ڪb-�O�,dU��9w%���c�ѸߜH��W�\7�RlH�l����-Imsc���Jq#v�\���p��R��	2��y������b���������F�gǯ�>�\��A�KJ~	��4��(,Vo�\����J�����bG߮��5&鋌������=��Yv�gd�1�QՎۖ���5F�ly�6��U�?A�,<�.?y�uE�3�����k��ק��~��皤h�7S���Ta +�ހ]��tH���~x�M�����,��\�n\OY64ބNpj�K ��!1f��+_��3���4Qdk�K���y��LZ{�0���(gePT�!���<-M;�ԁ��|� �ҳ&Tc�ꥠ�����ڎ|��b�'-�	ęZZ��-��L�I6H�/�������[����RK����߄��{\�
+M�8Ɓ&C�˫/���3r�%7	�)�e�X�:�����\\�����}b��8����	5[�,o�5G3�i����{8S(-E�����~����-�K��w��ܠ;�y�M��.�b�$�m8��Y�S��`�#���+Q���3ՙ�,�a���0|���&��p�U�h�;�����J���3<^�ӟ�iN��ob��DCU ǜ~J�9;�BB�Q��S��/8���W�;��1	o'�z+�{D�H���k������[��3)*l��=kCU=.]7�c��x�ƚ^���>�@L9��CPsF)��'q�^��v�ԗ^�}0�Cp}�z�E�Qx4c�<�ٵ$�x�]i�FG�rK��δ�D�e:~A�q~J��1@eyiف,~W���y�]~eQn�������R��cŉn�1�A4�s-��v�C�=b���ET��ztYi~ئ�|���D�^�򳭓���a`� M�T�Ƚ�W2D��
*̓�֒v#D�7�#L�}^|��t�|s��s����H3�8�U�n�� �r�Ǡ��/��BG?��Q&�DM&A�Xb=] �\���Lk����:%�1⑗�
�[X��k|� �Y�����$sP�����z�Hw��#��gE��9�#!{�ٝ�O�5}*$�0.��G�O�b�`�]�*��*�l���/����p%�ܔ�;+j~�In�)p7������|BBv�������e4���X��������1k�3KmI;�'���ye��y���&���X&x^��`�r���u���deE��58�
nTɕ�{� .�o�tò�ױ0�x���c�>W�Cf꾣��h�d�E�?�*E.tL���¼m>�Vb��ͅj�FV+��ab�0��jd=��T�K�F�li�;?ߜ���5"�;=e`����_9}��:�`�/`!�$P�oX�p�$�"���8�, }4���[LBS���Cu`�bq�Nwۉ�x� ���l�b�� �9m�iG`��E�(�9�P���ů�1�M�L_�֭������W)��3��;f�k��ɟ��;��6�
3��t���U��e
��~���l�&~#��OčZ[L6g�,�"�t�~l�"=W�@Gޝ�黁^}�M��M\�7�m�<��/Rя+�c����Mlu�hwL���O�Dq��V�W�H �-�+��?�@����Ydh�X��̙�@|G�-�x�x��h��i�E���= <��^�̽<���C���7�Y6Z�Q�N����*aD��L8��&�� � �tsպeCt���}&ٗ���_�K#\�a߱�w\I�M�N�t݈w�m�?�����/T��Y8�T�$Z^�	ڜ���8��-�hPbpm~���/z�QO�5��YfK1�|ub�bE�.s4�3氁E`/���y�����dexR6̅]:��	e"W��#)��9�j�?�/xɟ��oP�`��7]��p��`T2(�L��2֮�~TMx_��!Hӯ'����� ?�
J�\���)[`���TD�S��ȭ��`	pKr8y^\�"őp�o���lf^�=�\���y�����f�qP�BA�4�M�ql#9��9��.�[J�?Ε<����q-��$�CBJ��-�������E�6��^�����k�/C6�G��d���M5z�C�ũ��z��̱� _���p9;���38�P"��������T����J�����a�)�ݑ�קr����ё�TNmҪq�����~b�rb�
��V�)�',��}� �U�_��$<��@?ya���������q�h��6�\�	���ic���$dq�����=�2tN�=��atb���o�Sb^�Ka�݋��� �M��%�eёu�����W'�����"�z>�C*��>���*�ֵ�"�CBc�YdKKD@H�y2謰d���m�M�D��x�۟>Ӂ�x�5��R�B�D�ֲ�����Z��G����0�z-��%$-Y{�<::
���� ���t�C|O�\) lk�k�>o��n�{d����g�:�0RN�Y֟�ZPIZ�����ׯ����B2'�����7��b�0�4�x���Ka�s
�f���R���|H�����7�cD�g�~ߋJLƈ��%��%6���.���o��xhZ+�*�ȗݫ�RVָ�&�-�EQmu����a��������a������CJ5*�Nl��z�[��e��i�V��}��"�**�	�����&t�e˞'� �����,��� ��C9����-�Ү��4e*�UT��z��ʂ(�M[�����3�����Ԣ��4�����K���Zm�75�2JoX'p�a	��n�?Dɉ�#Z���Te��8���C��<�)5�p)��^8�ո�?���^d@���xi �8ΚPm�T4� ��
�r��2�eh/��0�)}��_�/��?�>�e�L�l�����"�P����N��IBY+9��f������J�:,�\�xYi��n��!��=5�lq ��9�3�ގA��F:PןQ��|]4����
>eDҝ�l���h���:'Y����K���Q��nO2[P$Ʉ��k�e[�sH\�<B���/]��v�y"�`�I����p9,����.ğB�~(������Ӥ�oR�ӌ�=�����g�0��nK,��y��$�y!]�G1K%�6�"erh��k`�m�(���<��V��"	��:�X�]�� �b�����&iZ���K�Z+���j+����8�B�ި(�% F98|��S����=*pD�xu4Z��o�%��`gY�j�T"��hm�O�1�,�$u$��j7qn"�������z����ퟶ,nxr7߂��HR4�@(��ia�,T��z�(L|SR�FC�����Bwo+��5G��B)��a�/,yE����F5�9q�������P���/�IY�X$�v�z�-h	�gf�y�{R�\��tj^�v�Ơ��\�l��b]��sU2�)X�6?ug��Y��~�!ӯמ���V�j����}��ϫ-�ۆ�x��1�����9�oE�+���A�~A�3@-|OcW�k!x�.���,R��.�,�G�0�X��ޖ��gx���lB	[B�~׎�ԏj ���m>�k͔B�d9��;�	�S���x�n���l�[��V��V�������Go�Ћ��I��F���)+B�ꤝy���)��P���j�)ӏLPD�W�q�=��ۂ������o���*��1�Y�pb��Ť�}V�I=�������U�x4��j&��I�<̫~�J��p��Y���?m�O;n�	��@<�x'�fs����.b�.��$a��`�Z����"�.Z�βZn��u> 0Wl	D�����4I���q�Q��Ю$�F�e���)�����f����xe^C۸r]�<��qE�%�����P����V�� �]���M0�c���N�B�鲦���x��lD�&4��ط쳼�ӭ����DP{���tK�@��CLjz��v���e��t���iU5�]#A+2
Ue&��x�����5����)���C�q��ʛz&�[{6�)0�z�P�����7ߚVUB��B���ϋ�>[M�o#
F���������q�";ϧ����o�^5uV}�Ȕ'E�
�=z��FdZfhGL��4�T���;j^d�ou��oG�����K�DL!��2���� M��l�۹|ȳT@�_���>��o�e�B,�~�)��
y � �~�D��6�l��*'�R��l9}��MK�v�@Պ�������I��:�r��k��`�l��WI$���
���%�a`ZR׮�g�w�����(�E��t��`���d�9I�^M�Ĵ��+%�\��-�߃Ư���~9J^=Y���"LT��!���TR�Ϧ�"���i)�@<�-�-&�c7LC�Mo՚�{�89��늦��uV2F�=9��F�^�����z�)����������Kθ}��OG�=SG�z	MY�[���Ʒ:���ʘ����T�33����+q`����I����2��`�hѬf���0-"z����
}��>���"��܊��ʚ ނ��\}���F[L5p�M�˷���Z�~0Ã��i�����ŵ�!��|�m9'/2�N��e\b.6KΒWr#=
��'�bO޵@C��|5�kC�yr����j��WkI��1��� ���^ҢIɻ��~>�/H��.ȅ�L�ԫ��J�O�,^�g�R{����*S�>@��hy�<�U���lL)��mm�����g���:[����ܭ��z��ǅ�B�4X�;]�U1�'(��+	���̟�'ղ�#;L B�no5�e�!�!J�giJjO�&��U��_�`�ɽy>If�N��Zk������~~���3�{z�z?�f
.��>�-�9C����c2	q�ܔq_V�:��mj���c�|�j����'F�l�<<T��z�`-�p���ABHq�8n=�NҳԦ�������L��bAj�w�|���X��n��f���b�@k���m���'P� ��Ć��������������陗9>�gM}��u.�^��ey���h%z4ƀ���}���y�AH�$�9g}$:{�����Zg�P����FjK���l�*A;Q�����~D��M�I�� �?	��g&b���k��B��7G�^>wd��3��_�."�vI�������!Q0�F� _m�P��Yi��%��R#YL
!�$�Vt�r�p-0�d��v�5,,ey�;������3Z <���L= \ ���:��i��d�2-���,�H���N	vm��@�ps��F���H`W�o�l�MR::9C<���nL�9��)~\��L� 3�����,��-��Ck��[�$y� ����9�2�3SS�U֍y	�'�D������w��}�O����������r�s����~�C���"鮥e�Oȍ	������R�K�uÄ@�F��Q�Cj���N�Cr�=cƄ"x������?o�++�]�J>,� �߲>#;�@s�;�cs�6q5Lo��| }�1$%EO���h�"ܪ<�*4_�RB�~'D1��m�<�ڈ�%��T��ͣeaR�!�8;�+�e��m�{�ݕn�V�uU�J�[�G%Nm�f~� �=��C�D1a�\��\�0`�D���"t��ر�1�n��RR^Uu��:}�+��z�'đ��� O��?�u>N!cvj��Ԗ��Lq<����GH��f���k"��K�Ys]b�r6�4���-���
��y}��@��Q�ᧈGt��<���Q]�.1=�|�r
�,i�W+>��؉�O�W���c�}x�5^�����a=@�ʑ{,%��e�6h�����F��C] ���m)"����&��/��qz��@Sz3?v�n�RX�]�ى+��gט3aPJe�ƞ;U��E�l�y�������Ц�	n�|'h��{j��[^�YWMW�D��ؽ?�`�e?5�/vj�_~m���^�
mG����c��EW���j���ez��ޏI�����ty#�G'V��߿��`LL�*!Ѱ��t��Յ�^Y##����,����"�	c�9�*�^�N�yq���G?�����ӯK�Kks�TA��]Gˉ���r�:���8uD�v��4Z0��c.��8D�`��;ת�W�#��[�'<pw��,�A�&��f�����nP~�jjZ6��n�sT`�G���Ii�C�y!GgX�)
��G���|���,��>nO�q��|
��f���=yR�y�5�?E�YG�+�آ�
Ԉ��5�Y�檨/~�KA*���^��-�ɶ��M���m�P��^��7��s�C�o�ݱ_I�GHx%�4)�l��j�R��4��Z�(�J�ۥ*��_p��ս �����IX�I!H�8X�#R��;�_�Y�
�����F�~�5*�9�O������S$���S�� b�?��P�e����Lm��>۽�G�^�|�tˊ$W�
��!65�:� ����S�K��F&�C�a��3�	�G��%�.y�f����� ��+Nd\��!�*����⯬����9An}�1��L)�"��ӵ�&	��$m��7&���w�A�"C�|�m5�B'��7��f�q�X�
#f,E܁<;4QZ�8:1&s
ᯤ����c�A��ak�&����/�}U$���uP��P�� �"^y��	S��I<rS(R�w� �)5?��;��TgIo�_���G(�;2��|W2ғsE��f	x`��R�E�w�א���R��3XA<�k �H���DƤ���Cw��� 4�0K:	Zϯ*�]n�W	m]��yD��q�����?��mi�|�㙠��i!t���6�M�&і� ϴr�}b3�_�8im(׍T �D�h���
�B�*&�T|O�9&A_�F#��ٗb���c=�E��8���e��\��wԛK����b�n��)�hV��a����韘��?�d�P]@�#A�;�7�ň�ؼ���߯%�����Ӷ���t6\=:��S����O�[�6_z��q�Cܿ�p!ၤ�9@��¼�)B>+��F�׃�OC��A��g�2�]J��� �p��3s2R;�ـY��z�f&vIۧ���X~�#�7�O��O�o	�����?4�8��s�'�B�(�֨lMr���Y�x9w�j#���h���ը:�K�l��p^q�޷`�����EtT��"'ǥC��j�j��Ҭ^���,���ﯶ�.�*��>�H��a0�,df�CD<�v	�v��>(h�TD��6Ȥg�n1i����Q��ĉ;��a��IRx���,/��^^�˥�����w�!�C?NN����K1��\��$7�"Rf��y���H*Pd2N�n����[�L��K$��$&�P��7�^�>�p)o�h>����r_�����C���a�è����0C��������q��?�&����\&����f�)�[�F}JA�(����b������y���=�y�`*-���ՄȘ���PH[3�_l���� C}����[��� ���4�]�͡��XQ~҅�`��]�x"4��w�$N�X%nc%?�I��b}{���7䚇]yi�.�5x$:C5����ǜ�w���p֎�.�o�(=Yn
��za�Dg�L��`� ,�:��7�BVG��9&�+�i��EP�?���G�4��hXp��/㟺;��CQL}8�R�����#������HÈ�		ɱȮTi�i�^3[\�C� ,I�M�Szy4�.R�-�+n� ��LJ��������2�ܽ��N!;��X�ԩ��6�p��ٹ��I�f1AEHy�L�� �k�����}=D���1�@7�.s����g�d�����U�1E��l���-S��F���h{t�:'
�qo�7S�x�3?�'`�C�	��꜑�|��`�ӤI�[B�ʩX4��6�Y�O ��`�X�*��Wr�:����q�!|�*��S��<���7[�` u��͙��hW$*ڴ��B�8�EH~��+"l�}鑠K>
e$�P�4B ��h�`v�,�U����>AB�(_v�xJ�T����)i�{"�i01s��u�BӦ]O�X���
��D���i3�"dM�w��Ŕ�C�AñFj�F	��HA m@A�!�y�ϗ�r��l@Q�/1w$ =:�����MN����p�N��t�'�6�.�����]�ԃ����w��F_L���u���0������9�9@��7��G���NĎЄ���w�Eqۄp� ��yK�BSm��#[1s���S�W�aP\R��ۋ����A2�����ϯb�/��5`�ױ:Vg!+ZU�(��`I��Б5b\�%�;�Q"���$8Р|>`���h=�����-��L�C��#U�',�=��?�$�N!׋.h��rT!��,�q\�yJ��ԜP�w���xL3-�,��#�b��m~�տ�۷=B���юy��& :�;�/���Y��$0)9�����<�c���SY�2W�ml��Q;������GN����i���?�h{@��+�nO1=Y�aaȅ�'�����҄oD��4��������"�,�ў�?)� ���i��~�[���%���59Ө0aP$ڝ8}�~���
�"���X0����j�"�C�=-�E�J��5c��yr�'?�{:VnA*/��Aў�^�(7��U�'�z�H_[�3�܆���:�L�SG��N,Ki� �>�>	�{}��� I�:�c��V�y�Fs��ҵ<F�m��Q�<F�L�?XUa����2� �R���ng��:T��N��x�~v#iN7�(��c&7z��M�	�>�l�M��t�/�R&���t��T����x��)��FƵ(�����0C�1B�1H�=��w�c,!�Np_�۫Su)�$�j��(�K�'��¼Nܺ��­)�1��3�1��h|4<�3�%�B�D ��^�O�Pcl��X�xTi����s��Z��#_�.2N>2�d����yh��<��g��_��B<��@�F�����D'{ݱ*˲���Fq��ꈭ���h�+�qR<U�J�Mo&��+)s��[δ2�GU���#�.:j~ێ�*qYԐ��24X�n����Et��������n:>p�[���!m���)潳Z�ȀՏ���ī.����sԁ�5�����s;ҘfG�N�Ͽ�92��ɓ��o{�aK<Y���P\�?,h������M	�3���x��*?��A�b]j'���\�놁(l��dR�EQ##�&11?lnA�iD����x��C�c���	���ϟ�5Be"/'i�>�Vi�����'u WI�jm��}�9��S�J����B���Fb�Gg�ٟ4iƸ��A��Rn��k���,l�l��X�a�}�����FI9�F�Z �䪐Ӊ�ot�kii1͂0�JL���O!"I�t4�;N�;�#ӆ��4��O����kp��!��.�h�}9o���ᑻ>�]��ftK͸��a٘��r��xֆ�h���Ef��R�����������$(KZ�8�c�\�R�E��NXqBGV��j��KMC��	�z��gB��S��8�Tϝ�T.��ղ'&�#�����#o�}�ʛbDj��s-�$,�+9�7&Qc�U$�"���6�}��}���Pp�!ހ�ǵM�XY�)��<���JjF�A}^��`��S1�����{&f�Ҕ����0�s������*4HQ]�𠒬�k��G�n1Y��=O=��|
!�u��b�3����U�Y*Vj��h�p�*�G��`�IZ��=�z�o�䑨J�����a�\����n�F�j�55o�z�t�EM���e������@bO�p�%�ILг˕����iU��a� �����LZ���I&�S�!��ft5���ծ�3u�Q�=���q�Z_t�U.����Cs�׋	F0��-r8�`�%���1~pSC5<Y���U�A�͜�ِL.����Hf�a��C�]E0zi]3Z9T�Ƭ� �C��=�'�訤�(�a V�8
򴨍`�
��$X��J|_FOZ,���"��{ŪP�AT�8��ag:�[xc�¡v�gI5M<-�Zӛ%�t���\��ڭ��)2?/t�?H�/��J/���3nu�
#haB�QN�;�w'U~|xІA�YܵݳM��1�6T����.���-~��rS�[���-5�3x�t`A"3��˔��4NN��,f��J{e���;1�}��������G�����	�EV�'5#[��p ���19E*�K�i�A3���}�.w"��!��v$�	�@�'~#ߢ���\L������SY|�s�q(Tҝ~w/'��M�d�l�n�m�&*�&5�v=s2�W�����G�8&@���N:&��=�0�X���v��\ zU��E��.�//O��ѻ�d\VU�c�>�!FMQ�}vI��
ؠ �?�[Q�S	6ԗ-��P�#��7�,��[��I��+�����;��qΟ���+&[����|d��*�Cӹ�?�Ҡ7��	�E�$��������fȞ����;�MM/��@��6����)"��8	��H��$x:���ի��9�҈�5�#M��*+I�� ��F�)�&���"��QB�oyK^n{5;�D�fR�J;�s=����*xA�qb�r>̈́d��	l�0�i��EɊ	ʿ���0p_���@��(!M���磣���\	H����reb�94�����%���uZQ���e�~�:�
e�v�]P�G��gYt}�M~4�����}��=l-1�	�mL�y���$��� �m�u��<����]��U��kљ���&OO��.>(~�H�����*��Y���8Q�Y���Zג�S�y��Bi�BƉ�
��(>�n9�Vw�^��4�����>s~��
��H���t�[�JQڽ8J�'C�-����| �N��t�?�N7	+�R\�sD��4*����<���K���h?+��pI�����hş&�l��������B��.�3�Y­��9�J�P�wz�.���a|!�@3��"��#����?Ń3? �����(c�����@-�w6���Ke�a��:
X�q^�-�A$8g�g��� z��[a��(�������%��7�9ԗ����L��z������f�/NRi����i�-*�֮�f�ݘl��#�j�01�u�y����=�oۙl��ӥ2�c�<��f���L�.�E�gy�fT���\�^�=S2�(Ep�!&1 ��U1\��{>̥N�($��(��� �6���Ն��R��M8~���S3?ڭ9г�@K1N��k�I��v2��5�0��^A�+��~Z��N�Z�7�׾áD�>MK�x[m���Ww��۫EGނ���qE�C|�=z���'$��u��gd�8�ñB�Ֆ�����pq�!�*qT�]�]�����[�̏Xy���ˤ�J�^6��Q(�� �@1i��_'wަ�6̨��I����ә�A�6m'� �y�&ԩAtl�g�t� s�h72M{ӛ!5LNCHӜKO���fYu~):�ީT(��T(7����#��3�N*���DԹ᠚`$�����>�]z�
�Ap��� R�Tc����2� �vy��v0���,��Y���W�ʶ۪v#��Ƹ\��hU�fk�X*-J�T�E��4ւ�J�NUD\pYL>"�s�^Gb�X8����$�	`ei�]�4"�o� 0U�w-�@�}h8v%�K�|6xonl~�DE��B�Mg\�#���@�Ф�@���_�F�t��tW�#+�B�	�2Wa�_JD=�N����"N�,����.��w �{g�*�;���ͥN�"��t�S�����;2M���FZ�܍�n���O��؜�˓L���zB�Gq�C�8�-&4��r�2K�����GV�y� V�ە2�V <3L��@�>Y����:��n�3�g{���Dl�,�]x��4�5��Q+�sļ|���
d Sd!���,���P�)�O��I�3D@C�ן~,�y�루 SlKꝢ�q�u]jW7�~�+"�K}i6� iT>�tWRRi��N �>/�C`��<��cS�{쟡�t����-yQ Smځ5�&�[ksƓ��:�u��X7
�����p��_����ϭb�>Q��,�|�=�k#�/ ^
"���z|c�������S�?�Sĭ+8�u&�V��r���,0�r*�U|���*��m��J+���G���hԡ��a%>���VEBJ�O�jy��9��S]NI#(HWڐ���gg��Y�/H��0�~G���
�0�㢓$<��j���|8F<��I��c̅Df���9�Ŀ��	7��V\��nq�֔%C���_ D��'֦�g,�����[\�� )��K@.2u�T ޝa`�R��򟶥OQ�6���s��.�7�s�*	/��&>I_��t�w��QM��i7�fϜ�L��}��s����s>+Y���N�wW��<�D&�R��#C�hv��(���t��Q�~q�6�ۀ��.���[��ߘVFh&����ûoo�J�P���
�GȽ����f�o�{�}T���+����룣;O��R��D1r2Gs0�̀GvM}��+&�f�[����f���J�,/�&��Y�Ԛ�|H������jC�>�4Ξ	�щ�&ܢA�uz��ʬ��M�`�8��p�����	��0�HW�d"O��$^ՏKt��,�r���s�+�k�O[��;�O�~�����+�U�Z)����{_5�:{S��)t1?E�)�U	(�c�.��/`��Z�p�:�"�e0o�P�!m�^�1�*5���97���&�r���.R)$@�sm[�E�&` ����I���^�x�ɾR��C}�EB�@��)C���u�W��;�v>5D���zZ�@�M�����!Ђ�ܣL&-C�.�aۤ��_�x�u�p�wa�r��V����/��N�2�����d���������[fP.}F@����"q}�]U�@����f�!$Z����r�X����4cp�W��:ѫ욉<����'�N�����3��Lһg��~�&�����_�CE������~��Ï��ǔ�9�B˾>�RE[izj~M��oc��.��~C�W�)��L.�s8= �F����{�RI����:����C3�(ƃ�T�6����E��Y�`���ީI��:z@��u��T�$e��c`�^�Z�������T1����R
�V�Z�z۪h�f{M�ƃ5�y�$M*�J�2d�0v	!R��z[`���}`7�[-�O̙�*'E�˾';S����F��i	�e �ۙ��ly�f�� ������j��?�Wv����\�pAfE˝Sgu;��(�n�M߃B��8�5�$$��nq�m +پ�O8ԋ,�@�Ko��@;ak�fޥ.>�����h� FRQ��K��l١���:;xD�5���V>u3ڞ�h�*3t����qn*�ۦ�ɘ�,_^��h�7T�x���B(�a'���P܋q���o�}VeCY�=������v�ü'�ɻ����Z
��ԘA��0V�c�M��ͅ�GF��_'pFR�g����7��m ��y`�$-]��L]#����w��Q�a�3���?��0#��|	J\��]��h�,�.���Gv� ����&��nm�$�U�F�L��,C�-��P��El���r8,���7Ub78�Ѡ%R���.��d� ��^sWJ��3"��P׬{�g9*X�$�e�'�,A�ܸl�����j����<6;U�`��-�B#���b�%��d��������[t�a
#�-�8'��$	�"/
$Q�
߇Nu¿�����S�X~������zq:z��1������y�/��[�:��?��Me~�<e�����]G��\a5o�E�����}�����R�Z��Y�7rR�Z��I���gj:��7����cLB��4��-v�c��G���uUqNU�_�*.
�N)���ix$�u�o�%+��9]+h�������.�A��d����h��Ѭ�$Y�T�e������ZB78��
qv8z���5��a��%ܐ��f�Z�����R$^ #͈��!��S6�v�gl5G�����v�;:}��,Z�����
"X�A��7�1͋q��g�E�7�(��}�P��,}��.\�-�I���/K(���XNkшj2�����lE���!�g����9v�V��ħ{]���]���H��N���,�l�6 ��R@��,�J�>3d�٢�Ø�)F>i���`-G���o*T�UEf�$�@��w�_��$U����̳��L:9cR�3ѥ� ���d[!������X�˞:��Df�U"8�Y>�gU)>Vm����J΅�;�7�I��=�	�53���\�љ�q�(e50ge7�D@r�jL�����\������r��&дE�\R�T��K���xCMr�n�o�$�[��������ay,�,f:��o����3*U�R�]��;�?��?����1����ZΧ<ӫ�W����>:�'���c{'&n+�j��ك��`�w�e�����Pi��4�s!�^'TG���N��`p�V��P��R:[A��~EF8�t�c�N5+&����j�Z��Ԏ�e�R��|<w �tH��2�r���z�lɊOz��甋ڠ!�PFw�����HK�'5�-e5>��F��^:���[yud�]ʠ�k}������7j,�S:�F�]#
�*� ���\����d�D�&Np���@� �66�P{��-P�'�����i���u�1*&�Q �������:e����\f�l�Bm��RE
��1��~�Ho�\�5��d�6<��t�I�@!x������;60�Ι���~����Ǉ�~m��En�����}i��;ݣ�ûvl��(2�������\N�n]t���K\���$�{`(��M�}{����\��%-��	�tA;*y#��3Oۘ{�?V'oF��E�	E}�g����u�g�� rȮ՚=��<��y�^cJ����sgj�#	\�,���"
�@���˱KD���cI5�wt��D��234��әr��L+����E8ŏ����t��{��淿��9<�.dU� $��^���b�
5��%���f�ȱ�`����V����p�*��t����*]���DXK�w�~l���G�si,2�<��h�`즜���,���?g��J�J9��"�[O���6�?uOAr�)+=B\GYe���!6�0�'��>N��c~jKؙ�%�f��߿+_� ��ze\u���8�V:��*��hk#8Z��M�����ɢ�_�U�(m´t��0>D��i��3�3U2n��w!���[�oX�0�Dƺ8!��{�ƫd�R>,'�B��]�����=� ������آľￗ A�ʪ�d�
B�+ҋ6�a�7ce��i� |��-Xލ$S��H[����1:�v�r� �}�#�M^lHtV�3��i�Y�� ��LM\2�r��N�	��� �}�\뺖�b��L1X�m�R������p����B
����%��z5�����Nڃ
C�e�L��f�� ^��<��u��1�����[!y�k��M<?�9KFT�,�����2v�s^���6m�����~�3��2����h���ᛊ�ݫ%�4 �=B�o�p�$���-�g�5��mݣL�K[=^\�ع�b�n���!�w��n�~5+��C�ϕ��/GUd$8{��#s� ����b�}���FO�w�RfL�c	B���Aֆ{^@�i�?ې��J���_7a�8}��5�<���3�n^�ᵚ���
A��z�$~�=;y:�u2�fc/~7����}2��hdsg�k�$�^R�|w���7��[�և&�B3z֝����%++���\���b����9��c��,	&��<��C6x�֠S�5��پS��ˁ529��`�4/k�<��僚���"V�����0���'/���2�N2m�o��y �꾆HBJ��'3@o����`d�]@֡��7
\����9�S荓�z�gL��e��H�}ѕ-.���l�6��#d:p��	&t�T��c���!�|�����كE;HX�6Az�|QڌW2��e��4W��1i"O�uO��Y�Vg'�@��qRW���:s+&�A�$��T!ˑu���%y��7ꌕ��7� 2LӦ�Lʀ%��pZ�Z:n���MbXe��\@�.��J+��Eq|aU	w�_�>��t��b�	Wez�J��
�\��
�0��x��H.7�!��w}�W��i�o���C`�!�)Xo�)�:��,��&�v��}%�Dqd�A�fr�[��^C$z�6�F[+�G�x�k��P�|J����ڂP�6z�1�3����Q,�4��l�ً�v �F�3vL6{�r{4O"?�t��J$A����P�#_33�p���
�^}̀e�ue%,�t.	K��ʒJ����N���F��B���gEe{�����s$�Qۿh�d�jM��<�f���
`��G����đ[&��6׬��^������M���ٝ���xV��cr�p���bBt�<��Z9�K��ۼEO��rntx^s� K�4���DD�l3f��l �hB�[=�&�>E^ C����y�u��($�EbTL�VK+G����S��rY��A�Ƅ�:d�pU��q��Pݾ�W��΄t𩎽9���ڛ2�ɣ��E���4����Z�߈�M��E�t(�TPޤ_�4Zx��+ɐߴrN�����ˈ>�C�=3��-���>�}��ڞ��"���I
���<[㓋K�i���`�Qsz�ǿ�:|�"M�÷�W�r+�2����ҝ�M~�߇y�˖$�s���˖�gF�D�}Ez�����ຉVŬ�Ђ@��uH����q���}-+3K���`��3���be�=�5��Z~c3���G(Dt��ݬ����]��2'�؄@��(��RK� �k��#�8���
\B�dD�@����_���W�ֱ� ���� �dЋ��[��g�SMP� #th�WS@�\�9`myD�v�֚��
�L7�C�o^9�$�k��8��T�[/À��Ӓ:��;-��Pn�-rKs��e~$�ht�$�糕#c8���R�X��2}|�`_�fJ�����0�I��U^�2��	�g����c�P�œZ�M�_�tzeG]�3	=�[I�����l�rDZ�nI]k9@��W0b�Ah�wimi|�����I��sG��o��xc����oX'1!(4�,)K�M�F���cm�>��m�$�z� �P��'�]��f��JJ�Y��RtΎЖ�R4b|�lp2lL�NS7��H"����Z���n�w W��� ���շD�������R�rv��ȃp	�N�pc��s������
��z�_�UC�Z
�;�7�V�X�G�^���{���п��E�DO�J&����ye�mz������K�Z��5���9�\�;I*��m$HU��܇Db��q1Gr���:��3�����&Vmq ����*ye,o�(/Vt�el{B�� Y��;�K��50�!7�������r�:dg�ˣƯ���Vq�� ��%G��T,�V����������k{���=���;���uzh"k++�؏�Gt!菐�lrl�!
��4�~f��kK$]iiF��~���fG^��u��s�t� ���(ܣV
�[.����ˠ�v�b-�oG���>8�9U�4>���E��F��[.�3�W63��%��AN���Hn���@�.�j�����l��C�*�!ȏCN$W5���0� $�i�,�FPrP�����`�݇C#ݰ��ۖaFç��t&��E>�:�*���`�ar0��9��ը�x��E�mg��s��!]���.�{]�F�;��@�x��d������� fM����6���$$h5��.�?���%���k�AI,�6}��^���ߙL"_g����U�����`c�ŷ�b�d�޵�R��n�Z������ЇQJ1g���r0�c)���g7$oQ?1V������qn� I�V*����7�7�b4dc�Y�X���Z�i�R����H�������d�A9?U��HRtk�?'
��V1t��a��B���fB��̇�W�DC(��j���66��PL�y��il�/�ߏ(��,���~��'0�G�����1z��V�9��qG�:��J�uF܋Z��O��M�XMH�����hX�X��?}�8��X��(���L��=�����H�epd�+ZOV�--��,qZBi	L!M`߰��~D|�U%�?�o�7v)� 2i]Jb.����G����Kb�� #������2���[i�}Ul�3�<|�=���L�1��5v5ݳ`7V�'�ƍu�2��*bW��PJ� �&�g-O�
�r�U�Jxx�
@�`ŚKR.�f����;N�J��?��R�4�{X�,���1~G�6xW��*��\�q��3S�9e�[�e#��"��*֯��st�Sy��U��ٳj��6�B�Br�/])�
��)�?�˔谠r�VX�?\�=<
�3��u�$)e���NEOԎB����~2Ft�,;������c��Ӟ�P��8�IM����!h!(t\��B9M�bz<?�IW��ÐFo"��Բ�[?�D�E�@�����kM�Z�����B#&ӈ���(�>/�fP���$�J�ns�-��[S �ش���~R!�%����>ewK}$g�2�#4��h���P��^�pv`����V:�M��Ff�&� S$�E|'���g���Z|�,���>ڻ�i�9�����J� ��q�M��4�~�3o�X�:L�|\����lVpKܮ��P���-vh޺��0'$�6n�6WDt��i&7�]^:2KE�Jg;���zO)E&��en��r�%o�7�C���W곽o���
-}s��`N�M�
A���"��R�&N�ڛ�+'H�8+�u�g�������/Ĥ>��ے�m�`>��B-�E:f:�L�LF���x?�=�����?����G
K���6�Eå�&E��h `��'^��|h2���x�=�C5��m�0JH��<�ꂓ(�|��'jr�Ki��/[�,����XK4��E:R
�Ģ�����3I���%.2�����OH(t:[��C�ù퓋X��/��6��zO�>Mߓ� @�e������$��+���r��yg��k�l-�G|g���-��ĕ��d1p�����%Xa�3P��c�J3��'p�W+��������
U}�#lM��i����}���jq��n���n�S�+>����k8f��x};�s�<	Z-�(��"Ȗu�\���&HR��"f�D
΋0� �W>�	,���+i�H� d�P�/�e&��9Eh)�i|9�(;=
%MgK9�r���:#�brpY�* V��|�ݠ���ۿ s ��n _�}��.<2��\��ͣN�"��(�F���ؐU�ur�A"	��"�=��?�a+�Y��n'軯IY.)Z��e᪄({'&�JF ��`�ض�OQ�3�ه��	����薏�u�����*���剝/�<.C$5@u۸Z|J_�F���W�D�
�B��D1��+�`,(�;�wp�|�,GB�˰�U�� rg�y�d��6I��<� ��b��Kh�">���_#AƘ&�L���D���8ϋ�k\I:J�'.�ܣ(��]�� ���Ա+P�(A��/?8>��������	�[磉�`����/��Xt���[8�K�Z�P�����j���(1�Q�m�3��i�}h�n��=̿��_�X���`��PY��#1w�w��O��bj9����s�� )@s��F�e[Zs/���/���v
?͛�'D�eiH�~U����
Y��~��ڴ���LjN8q�UW�4���2�8>#�S}�\Lf�7�$gx!2��ם�$��@B��~�]=��:����_�kWŬ�� \؀��:+� `�\��{C��[�IXh'�������9��x��\�X;�:�4aR.�K=���u�f�ސ[=kN��d�!W���/š>nN�:�-�о^GD3&*;���Qs���ߔ�(��9=��'�u����L�Z�KV�k���q�+0������+��p�MY��lss�Ɋ�͠�J�����y��N��M�Q�a�Z�j�~���t �%�q �3�:(b��e.��I�H��Y�QuT�d`�����e��'��_���l�U?4q]�$i������!Di�^������ �rg�f��Am���#{I��K��f���x�!jUD��^`��v&Ĵ�����cy��G�e�#r޶_�7�d p<�T����e�=+� S���}8�3h��gR�[t���Y�M%�@������3b����\�f�|�:^4>`[����ΟlWct4�����y����[M�0�I,��wZ��V��Ώ�S!MX��� ���� Ú��:��ъnس��X0�u���O3Qd��!8G�܀�p$�u܈!E��#�Ė���7̑�!��o�\�,,ױF1�]KV�}O�{0�v�D����}�z���$ԋ2�vc��.UI���_��8ژg�W�#����f�:b�z���n͸s����歸�cUg��(Ɂ����\�j>�����(Lx�m N�4��hQ��,ui��pt�b���QY�A�N]�Ֆ;����>�_H&�H�d=��cC~P��'o�VI�}!.l��(Y����V��P#���H��nT�o��_���:���w�&�|�(0���?�8E����J����P���o���n�b�w���(�����ݻ���)�J��K7��<�jl�������ɑlJ&˲<W:~��D@��C<^�	gZ�w;&��+�t�k|J��������1�;�gq�y��&
�&���i�
�K��F t������	 �eLvD������/J��V��'eK���U����cN�`9���s܂W���B_9�g���J��R���x� i�P�\�]��Z�ߵձ�`��K�r����36Q)�"�KGl���;�#��`�a���[�n�;5>�M6Н�_l3��&��|c 6*�p�(C�'g~��n$����:��U�qb{גTW�er qR(G@�:��6Ⱦ��K�Enш)E}�ɘ)߯�>�ⷺ��ʿ�b�\�0�=FB�ڼ)����U|F������L�iB�Ꙟ�I\��q�b���X*�����5(�J��2�~�����n�2z�� ���vj�;�ݬ�%6�]�
�6��B �C��2g��r.�e�a�ԋئ4�t����L]#�<$M+e)O�p*G��b�J�.�Z�|���6���D�P{k
f*빜��_۵b�H/�x�B��-�$�ŉOٿ�AGN�1��52��H�
ʝ��X�O��ME���;^�a{z G'�~F�X�K��OD�bW���#J�BA�b����q�{� >������Ѹa��ږ��z���L�rF�w!�&K�{��_�V�kr�IdS�H�i�S�z����O��f�=�g呲1���⟶y{��;Ѽ�{�+]:��N�ھ��ƝEl���-G�E�.���||�z�uݘ�}%���`xXtZ/���<qM�ag6�L�*���^=�v"f�^d��m�29�2�A1�<�gh���Zo���9OY\�&UU�����左��hs��h-��PR��-��(�� �*/���W�?!���Z��h�F�L�B;U��S��X!��C|X��L���g�,u�E%\}����_E�+���c�`{'��5G�ѫ����аI��� �k�s;§���p��)"G
[��X�g6u�7�ˁ�;,'D�B��P�EF;ސk]��W��3�y\����(�H�a��L�C�X8y��u������U��M��$u��[\�u���x ��vD|�*
��4c0n�&5�&lv�/	����6Q�VF�x�>@�Fe|��4Ǎ��u��{U�1a��_�^��x����7����5��+�Q-0��y a�B�ʲ;xnQg9������[�V���|��u6�x�"�EC�������8�`�8��Sh��D�3�m���i�..3����^b���L=��;E��\b�M�����(b�OAѫ��]�R�Ҏa�U���!U�$1�)�I�%��a�Y�#m�׵K&�4�F3��CWH�q�EF)�a�ي�� ��9s∕M�T^����p�����_�� �?z��}�}�֦!�^�:�#b���A���y�&|���N���uzw�qkF��_n7"��%�\���g<�(|�L~J��|VE�u���$��������y�?�zhs��a�*���f�U�Ogf?�)]W����ڛ�q�c)�(c/�$�n���<�؍C�5F�s�*��Ϊ�V;�UB�$mx���0}��֝���"���
e�\v�-��2��C�N����PU)��%�#~�}�U����a��g���"��6D]�YA$������ȋ1�R�$�[�B�_rf]hR�A/��ýDQ�wi0�ɦ*����姧����B�s�%Mth����_2���w�jT�Σ!g����,�v;�O0�\\�J
|����6Y	ܲ����,�|�e80F��ݏ{�m�8b�*1��݃0O�� ��[�'W�AŴ��5�kF���^�o��~MPJ���ĺt%5�c/|�:zAs.�9�}ټ��I�g����u��B�% �8薤�sj�]@�Ӧ�-34[+Q=X݂B�w��Ey\�%{o��
���j��]�$�-�x�L��!^~ǢV�YQ�[�ƉuDB��V��?�����'w��s���-��m�6uGN����ܾ��+�\�i/V���s\�t9�z	L��ᝡ!���r xF a�pJ��n����A&嚝U�	�hڳ�#]~��VQ(g�����%�����T�
��O�P_�<�n��O���~	��-4�&7� ��x�p?�y��g A�]�=ޜ�n�0o��>z�n��p^��OouA����i��&�+l9�<I8Rn	�����Q�������x�^m��a�6!�V����!@t����+�7��4��E�/�v�5�e���z
��e��k��\������lFS"��/F�b;L��+�m)�36+ ������?�g�W=Z?�Uu��1X�������KB��;^�CUW��>͐'�=���Q?������8٦�K����*�gF�e�gIG��Vh+:y����n��w��)��rr'�}��w���X�|u������k0?�v�e��i�v��H���}Uq�Uu�)��ثK��R�%B�TE#~U�OL�ˌ�l0�l�����"F�A�{7����]@����J��FB��_a50*�֌F:�b!�}r桟Pis�C�n���+B!eTy�Jٲr��u$�Y}N�Ǟr��!p��m�$��}ǶŢ
��Yy�ЃI��qa��Rt(����%bWk����
3]_a�3s T"OR,��1�[�*�ڹ�$g���i�ޠ|M�����kޓ}���Z;��P�c�C�gL]�`��wOsIb�3��M�ঠ[�h]���Iz1V�l�S)���'�����s���b��Z�o��|Z?� ��z?+�p�'#�8h�ݛ�`��8vtng�#��3Ƞ���ݤ)C��ܑ��'����cO��m |�2Q��Kڔ�RN�����#46���c��pK zBy9 ݍ�4<�����{����3���v����Qahh4�Y��;����10�u��y�<����S~ߍ�us~w G������)W�Hȟ/0�2��逸C��i'X�� cA�����&�ﷴ*$�� GzV���?87��-�yh�B�ksJԞV6=Ғ����i,U}�����Ɏ4Q�ϕ���>0GR���SY*�Z�H,:1o��@���8��v|0���׀3���@�Go�h�a;�G/���<�@��=�Yh�c!��,)�89V�c/cpϛ����Y�)�K�+�(�R��p����: �B,�Σ�ګt�]��܌�ҙf�UQ�u��8�,aH`J�� )�>
��N��J�3 ����q[M�6Bv ��8����g�G��|�ҍVe:B^rq�w�_��p��`?h����&�ݷ�j� �Z��2Fy� ��j��M�g�iբ"e���rﯖ(^�c�~[4��sj�\�0,#Cy��V����'sXg��	:���#KB7�1Cp�u�J��w.�k
�2,0�vz��}���/6��-�T\Y��Լ�8�0��V����`���\�(9�57�Z�%��sE$Z�i��-!|�Ԛ��6��V�}��^ή��I�>v�����S��W�WI���)���ُ��Uyh��6�J����[&� �(d1V�~`3Ko�pc]6��������)�Rm�����o�[���Qq>�`b@5J��-��&!Q�\D<��b��"rV�����r���&~q���Uu�l>�[*=-=���:�\*2{��!�ƛ�h�5��L���"u��3��f-��3�q&<W)����K����7�`�����y��Y�h�/ß�	j�ޛ����U3���ܖJ^��jm�!��i�A�u�Lu��F��ޚ6�&�	�w,�B�M�i�����#I�AU�����t���e�lZ�Ec4
�����5D$wBͨ�g��� ji9 [C~h&�lU�lI���̶������#�D'��QB����T��� Q��,��C4M�祌^�Șm!���*ҳ���B{�ܭ����kN�K-�zWل�,�Z�I$�?[Č>�B`�do��O\h�E�c�{������0��D\�8�����+��ͼP��V�����2�	��.�d��Ewϸ�,_�|��_n>߀�1!�V]i<���#�2rۦ�/7CgQ�<��^h�F�)9�3��}̛;c���;���{�e0����j���6M��a�C�d�BE��mؾ�h������
�S��2���B|�9�Th9:��D=c�#rոF4��Z�;�4TW�ռ���b�4�Q�C�Pu��w{�$�S�B�&�.st����i���e��W���ê��� 5�z��~�w!{��Y�	��x[���j]T�NU��g��~�N�>7eT������lH�X�k[Jg���4��m�����h��%�y��C]�PTo�&B�L�tR6
�F\��3������� ~�o��w5��دSb�e*3��zv����J�Ӻ��;��ϡ0����]������2xs�Q��?��8��@��R�,���+۸4�={��	D����i�q�+�)5���V.�c|�q�!�r��8��2t�5v��]��ka-�6�/'[º7E ���f��n���y[g"�6�'����׀�m�"ohN�>FD�ŭ��8�\di-��@��vL`IDCUm�^z�<[���:d��$(	T��5�Ӧc+q�"�#��~�5�G��o)'?�k�'�\������j�a$�%��;����}|��s$;�����Z6K���=��/�C�_Ow�ti��S��v�OY�/e�$��G��J�iݨ���.��L��/�q:BYg^�7������b�*��.������#!��U���%������pυ�H�O��u��zN?�$��ɹhU�0�5�V/�ܟ��}�12���qz�$_�\ ��f�z`�ZP2�Y^�3����
�{�S ;:p5\FwbL��/z�,`���o"�W�U�r�W0+ȿe�e�>ʏ|Iq�Y5�o�����:f>8���,���Z��r���&�̐5�>]du燬"Ќ�0�l��P�As�>�+5��[��v�*�r�[�]fܵ�Q�B���gl�Ku>����5�C����� ؜B��B��n4T#��j?�j�oԚ��g�B>����>�tk��?��C_JMp�b���ɖ7,��%]S��'5.��o�����)s��rO����ʉxԙ��F z�s��i��70�\�/�jE������w�]E�!��?.�Z�uɞ���J�6
ï�ڙ�K*�ܦ�3�; =VY��믃���+na�J�]���#!�WD�/5�"	s�t4�.�U+��c���7���m(��n谍2���u������5� �U�5g�Oy�m{��ab	�)Iy����b��UDJ�������"�nXիҦ�W��?�R�_
8
2���6پů��.ǟB�桂c�T�5q���j97����z���H���"uKm�+Sc){���%��}�fx\AR3��G�گ̗+��/�!Hr;� R���N���%��h��d��+s�:���zI1A旗�{�& �;-�Hy�n9SRz:_6Q9�Ћ`Z��5��V��ވ���[^�d�VhI��!�ĵI��᫪ɫGtr�c�8vIF��;r�LX-'n�&�xV>����M<EX��?C�kXr-�� \:l�����2l[�䠋�\��F�m}�Cy���gy�=���i���+2�arb<M�\�䂾G��9�d�}��#(�u��N�b�(Ƌ@v[�^6]����Y���г%Z7����cG9yڕ"��<A@Ƒy/�\Ve�GY�f�>�u�]�3(tB�� 'jfw�J�~�t�"q��p��MC����L/x����������=�|7k��ʧ�&�~���
�`��HoX�n�7��^o��<�Ǹ�v-�d���?�/iTlϒ�v��G��NP��`�SQw��� ��7�A͉����G��?��L����9��`w�/�J��@��WT��{�BgЌI9���MT�F�\� �6ϝ�In�	�n^G���O���YYm� qi���;@~�=�19o�)�{5�y��T�,h#��*��ҍ��Ia�#�~�Y
���#��������jS����o#myYnYs�.n��I��3?I�����zI�K��b�ͭ=�=��᳐k�!������Ng�zB��ym�$!���4^e]��*g<w,�}ُp�I��NַO>,��ui	�N �G�צ�D��L�mX	*���o�<C�f`��Wo --��Qޡ��m�7��Ku�8&"�G�~"o�f�ܧ�	t�R��mVu�~U�?p�9�	*��I�(��>8��j���K?�,Y�ܓ&�x��̀8�R�dE���_��3��D`�*��*��+~��u*���{�չ�wU�Ŷ��*���행����z�l^$�40i�i̓W��y��R-`��4N[��&7�o(J���8tȏ������S�_2����|�a�t��᥀�Y�?+��"P�Q��l�y]�i��Q*�&��cJPx1-S��!�B�X��<����G�XA��&��E&�����1�!u4�Avx�pK����zwY��z��r��B�uzP��"w�y���m���i��CX�1�#[eEKtPrZ�mvƤ|�<�tߘ�t�8����f71S�'�rm#زN?��M�T���<<w~5{h&�Ys1Z�8>�Sw]����촧_���
џ-1�s����_�J����5)��=1\#vŸxϭ��Kj-dF�{�c�N@b��f�pXq��&�.hF!;0�a��;�E:ԗ`2�-�O�k�A{ix%�g�8Ϲ�v��@nUѸr[P[\�ù��#�T����3�UԪ�C��1]�wП����Ӄ��q����Z6�ZD}V�>�Z�Jt��G�t>�g�
�t5{�2[X�?���"��N��[w%˛y��0�n.n�mk�ԣx�kBhE�N�2�X���:K�2��o.�`��>3P���tWb�	xQ6�Ńn7��i*H	s�:D��ZB3)ٛ��3��"�t�~�]��Oͧi_�b�?�EXu[%~҉Vn��*�t�_���_�Ó�~�<��WE� ک�����`�*����V8@mƥ~����vhq	��gC43+B�Z)���# ���D� �f�Y7m�.���<��.�,)�3�-ѝ���_���93I���+��w��ދ�Ū#xD��J� _L���GO�w=��wj�D��B��t>4�Pb�п�Z�Z#v]�;$LA0�!��Q9!J�!w�𒍣���t1t���[Ʋ�AC*#���B2U��^�^��´kj��Q���&���ĽNCi���J�\t���j(Ќ���ɉ2c�]�g��*����Z�Mqc�ePb��Ug?�*NO�J��/�{#�~�ƥ����&��^�H�M���W��(����%��_k[(/�vv4��jc=����Ye�e��Fg�	�e6*����Om�.��"��I&�B���IS���vw/e��r�k��S&�6�Uu�Z�|�Rڋ#���n1j��RY����n7!�j�tW�7NX�ݎи�B�>j�v�/7���G@ڄ��~Ht��Ps���7Ի�V���!�~�8B��/�0���(+nA�A�ӯC�Q�c�,��gRV��n���.d�\q'�]�-�8�F^$r8�P��7�U�>��Uc ����R���Q�ԙk��Gz�	�n�|��b`\���"����Ң����Ĉ���G8W�u5M�;�		�Ϭ�8�U勨�.���M�KkF�?~����/^��Ao���u���]*x����z��=Ki	�x�ܧ���^��X.�l�f4�� �0��W&��ṹ�����JF��i�d+G�)�g�řpG�Y�WpBD*�5lp�3|�9����◫�n�p�@g�?��u�����|��bY�3��ɋ-r%� p*l��E�Ց3c�sX��?hP�˱�5�$�!�Yፔ��� ��4��$N�
j$��@qg#�"���&��+mͩ�����-���U8ڢ*�!���Y���⌞�fx��!����vz5�C�:���0��-<l���Nm�NW��_��WC��hG�]%���ZLCm1u���L�����uZb���5���;s-é��G����S2���{hM�%��?싖G�U��#4l1d�*!��OCV�T���R[`+P~-�V��U­@^�#^�6V����6���� e��k�`w�o����]�?>_��!�_��ŔM������� bL���ڴm����!s����;BcT���8��T��MN�u�i���5���l���2���8輹D۹�j���G�K��c��#��xd��"s�h���̜y0�O�,s��r �ȣ��#�3(�&H�q�(��{u�t�xc��Y�#6壅Iq��b�Q_�pH���c�[��t��b?L���,{�5���%�]V�y��Ce�� ���gM�	�D>�{�j��Qt��9:nL*$�X8��D̗���2�8ReB�+m�eR�h���:�I��4�l����jB s/4����G�!7F�H0��L�EC���9�N��6b�����ƘC!�����.���},�&�-%�R�N�leif�6j2I�T�� �
l���l���C�ڌ��
;�ˉ����j҆�36tYY��@����}���%�[�М�ooX��1���G�)�.���a�樽��W��\������*$,Tf	�y':�~��iƭo��̶�n��1�#�݂�������G��)6@�7��d0�n�S�tzz�����L�T�L��9��=nO�aǌ��� ف��&F=R���={x��	P/{���dr�`7܍z-I("� qT	@6�8S�v��LAF�Tk��'�8���'^N�-Y��:�m�Gr����,�m����ƺ�w�^�2��T��w��h�u?�y�Q꺝:���Q^�Jl���F$��=�Oď�g��� 5Y�%�r�S��3��m�I����*ڪr��3~-�6�	�~�E��.\V��X^߉-�.5N�9�0P�P�n�۩�y ���#�.&����_ً���A��'!�ـ���KJ����未do"0�Ј�7��
��i���5S3]�F��ª�/�z0�U'׿���%W�t���?��h�魕=�����[,DY�Xݒ��S�݂ӌF�ɥ]��!���m��=G�Z��(��Yq����M�ZM�Qk��Bo瞠������b�KND��#)�,xPr2(N*��o5�:���i��8�NU@��Osh���V����f�7���Ԭ��2{4��$���K�FN���?y� ¨Ԉ��"-���9�H��G��X�h�hݤ��Y����g����,� "A���`pN�rxߌ��.�����|�4���v�g�
�6X��6:�=�i�\`J��{�.�|x�o٠vm���"�)0�<�8� [ֺŻ�MV>�,�m�zeҭ�XPk�؅
!1�J�k�o��6�{N��$'�Tl�\�ԧ��H-K���H��P~Qiv9��gõC�F�R�֦"�wۨ�X��H{"�+2;�}������<K���qۃ��3oִ�hN:0���ө�)y9f��  �R�i>f��7�(<8>I��j(�.Tn�X)���,eSdA����j�x�� O��Ǽ�<�mQ�+��q���X^�QIܻ���Q3��H"P���ϑz<�^j��� 7�#����o��!s�o�5#07Ş �*�ω|�'d����s`2�~���2l2`2_��!8���Î��ʺ����!�f7&�?C����W6 sH�OQ,�/�����\�$�-�hW��'�vVL��хuس��2���B�^��p�6Z�:.��۹���Hob_Nl�v�>�t�P'xZ+�ꊀK�8�|i����*z	��
_(4�{8Ug�no��1:�E�F�p�+�^���ĚA���ۍm�_Fj��xA����������)�0����\~�jB�m7�����ػ�f����X�TBf��|�\��������N9��׷��V�چRAn`K�TQ�{(]����L�^�e:q��0� �NKg��0�OS�xn [��v&�)�9h�_��G���j�ap8{]hh�:������7�V�?��ܿ����2V�{���� �t��f�����3om�>�t���>\؎��@���.x; u/�1�٣ĚrX�#�hӑ���S�m�f�GE����̓Kjm�$Ao���ױgj�3�]I<%zPI�'1޿��Pk�)(?0��3}�m}���P���鮮#���o�2N�9�we;�a��q���h����D��4�s�o�B<̇^ߐ�5o��o�|)CXf!�0],�.e�~Ga���������}2XT�e0�\���Vk��z ��pU���"�	zQ'3�I�+�� R�`C�1LF0�;7�#L�Q���8���7c#+~�#�$�����F��
*�r����uv�M	����1���~~3p�Ԗ�f��'���J4�#���"�d[T�ѩ��U�
Wh��� cSxx �u5U=E��0��	&A,Y�W�ڑ"��?���f�� ~���~+�5!�TC�6BOC����gm���t�Ba��p�b��ՋF���ѷ;����<=;w����w��Q�,�����Fڞ5�0�����C�Jn�� q��� -t��N0�G�c:��4'bH��J�Г�~�|e��W���"k��`K
��	֤$rf���~o�M]\��(�!���9��8�#������u�sJ��4Bޝ�0L��1e��|���PBo���:��fG����(�������ڿ��0��"�������$O@{��&�z�}�u�*�n��M"u���[ on����������<��5�-Zr �ǐ;>�f�	����c�:/�� +�ȼQVA�����=>���쏥w"���AP�]{_��v�����m�ť�Ġ�>�V�>y�y�uީ�nq����+s��zn"r;p*(�����k��(�}$�
���e��6TVwc����LA��Ht�Ajm�Yl�q�,N9�f$���_�_�d\��a/s~&j��vS��h��y���Kp>�H��f�\>6�bD���0#�#H��iѠ�b���b8�
�;���n��l �|�j�f��� �c#�]e�s�]4�ɪ�K<�.�~6���s�d�9C�x<���"���C0Օ��J!D��e�K�v,FDǅ+}��߯�r���:��~A$�D����Pi�V��ʠ�t�(|��"K�G����B�莆Q�y���"���"C�9���'�a�7��vK�Y�ꁞ�f�P�)�y�q��2�Q�c�[]*���dÂ[=�ϣ��a���f��9nl�}}�8�W���̌<��p�p�WJ*T��l-����2k��>�lh��Z�x��
c�h�7�f
���<@Y �������u�q[X7?���i!�燑	�\��A0�d!]��f7�_G@g��5���r�p�-��y���E���߯͞󜒩�>\�_���eOb<�v3���Is��<�Ԇ01e�t^5bN&}�DIC|�O�!u��-��h	����&��eh�X�е4�u��jU����ǽ�N����.w2o=\�#���&w��e�%D+q�S7�m���aD�);t���D��&p�t��`���DȈX%0�/]��#"�	Φ��"׹o؉�X��s#v�Jo�S�+�L�U0����n����i_���"R2١���b8�o��P׽#�=l��h����^ٖ�㹔0���﩯��F�"�t�&A��nA�%L�����(�(M�X����gD>L���v�k�V���;XL�#.@��۠�c��:uBJ�Ը@:qS��?)v#vV�y�7]�h����:���}@�9q�Gn��h�$tKf%�r%��)p(�fT>�65Z�"�vt-0n�z�վ3����1�"�RZ�>B����B�(6-Q6��{ܞ�l�A�rB�Ҵ�Cc��V�#��.3H G��i�j
��܅���9�ɿ�Y���x�G,�F22�M |�!j#Ŕ~�ԄZ��;��"�g�$��V���jJ[�9�Iiֶ�/�*x���!�-�ꥡ�����Q]9Ty:ro�T^��{�7��S��2���V�օ�{ƒAe��cp �)U��+L6�l�˿?�jYe�Y���
�A�8@�7x�EOm���������n+6����w��r~`�gPA�^Nj�$�1)��P�����L�%�'�w�̐��D�Oz���Ԙ�H�1�M, \q G��7�fvܠ�V��hG��y�b&�K�4p���Ȱ�FiH��?UE��v�PܒZ�N90��K��B����A�s1A�go���V>K�fݭSt��|����
�`n0أ�|Р͙ZX5�wr�@��^�XɷT��]��������L������Vd�ȵ��o���Q��j��uGΤ�ŊdL4o������o7�~���^W����l��hEGi�zY[��ܸ���y�~r@�>*s�2{�w���EK0-�Q8��@�k�~>b&�o5�����?`��!��?�؂�la�}X,t
Fc=8��&S>�V̓U�Y�y���YZ�$&7��=��R�-�|��C�gW7~@)�?V�Y����3{�g�3���WX��`��u�݅H��~�{���uf�R&\�:�	̑<���p�_���Ì��dn����s"�Z�]�Ϟ���rNR��P�����rp�#�%/�e0N7��\L���t�l�'�Trm�^�eP ��Vn���e����^���JdJ�E��F��y��,<Y^�Pă�!���`EhC��N>63�C!�f����_<ٮ����_���&rV�I�$<H�mp.~�:�J<˔fA��6���1t�I0��`3����`�Q��f�7/@���cs�n�k�V���ZW����p
r�A�^eRU<�f�I���%C3#1l�g�	�j���ʰ�����k���ڡ9ﵩZ�2+�.x��+�0H&o�J�m�L�~�I��f97�D/���B�A��."�t��edZ[�th0�MLK��F��;�ʦ�g����		hڗ~�����>�7�\�{_�P���O.��T��Ք����mͼY�D�;�^�YEI�Q�$�����$���ڄ1GTɦ��z,v� ��G��o�Ѷܹ���T +4��nB�GfaS�z���Vm��I$�,wAU��ծ��X�M7)2U���9qi"�L�����7�G0���=EY'����E� �JC���"��n:�����~V)��K��#�p��x�Ł�jW=��'�r�-:�.�o�3�	X�-G�7��9j��5YԴӮ�߇�ob$��l��#w��O�L�a"$�U���^_*śB���V)�
���궶��:Q�5K��־���
c8A��7��Ѕ�NWl��X������1]	3�`�b����Z>*���:��0���x�dP��)3�i�`1�+�-�2���}�����j�^\J8^��[���c�y.��NzV�>z<kYb�!;�:6�a|�86��mL�Zn���}�VO&�Ŏ�)��'
�^�����p/�;#<������%N|�_�~��v�zs��,��ݷJNK�p���}W�y�1��ask����Y�O\L��LDkP�9�3-�_�Uh:H�u~�$�L�Y0���?r}P��^܋�������`%k��n�5�G��JA i� ��|�����N��e�U�UD�g�����<�	R�9�4C���S�CO��,��ic��,u{�ە1�f�[��e��R��Ifb��O�ޤ���a$-1D`�%����q�} �|"6�ތ�3Q/
 
aa�M �8� 2���n���9����{����R���T7cpǉ�m��ŋk>�$�R��x~ǗnS|�˘~bN��˘n�5#a���/�i����,/_�d�$S��؟�u��;���n���r$�ӹu���7��n�y��Fӹ&��#?<���`�e�������~4��"�rL��t��{Ъ�_i;����S3���d,����P&�ݧ�{�bv-"V�^X�H�TkIT�.! �>����O=Ek@�or��6e�t�WP���wwߜ���6;ZGٙ.�3�����*w�E�Tt$T4�ף��O[��L��j# ��J�I�`�sۦ��t�O�Uy�A�A:5���i���N�t�<!%�$�
0qΝe�����1x%I��D��v9֕؆_3���fcS4Nqaś�/O��=�
��D4��l�&��%�����QH��2&�{�.`������!�Ȱ��r�����#�]���P���x�ocS;ߍ��d��*K��Z�2�$��5�`Z�m4�L�����;_�v�O�ݕ�����	����n���mvȚ�C�˼�&wJ�̛{b�9?�O~��:�itm.�w24i2a��R�c�i/gL����MԇL��*c�'p���հ�K���X���e��x��)Wn��M�����!�荴*Tsox.`L}�V,W. cΑ��V�C\hےM��Q�%����&��]!���(�"lHĚ�Ub/�§5x �\w���΃׫�_�:��i��3������!�#㐅�Y�	eK�9?�|RQL�@7���
j����G���H-m<M8��t�g�b$T�ߓ&^>dT1	���<�L��L�a14���G��xXI͌d���C>��/�:��?]�P�==�+iYIA�,��˨�0~����DL���� 5��F���;�v�^03�Me�q(��n�2�V�I;J��yf��ڱ5�M��� *�&�40t�C�V��Ā4�� ��b�7�cl��������}�r̿��|,Lr��l�Lzsz�v�q��:�R���xw�����d��c�����pT�Yw��|#��8�y���h�Ui�+L�ӥ0`��Ra��>`E���Bhj��M�*�����-��%AK8�,nTԋ�m�c�'�Wr�����TOt�Hg�1O�R�cHgJ���^��y���/p�=_q�%	G����BND��n�\@4���ؠ�
�4D�@j4��;�F�ʆ4��u���A��
UJ�	���(
�}4"k���|r���aE��RK\-����~�ӯ\m���OI��㺝O�Dg��]�:K��`��N4-9+Ms����ydW� 3� \����cec��t����aS�7�Q�tIܶq{Q��
����Lb7��?X�
7���Vĝ���2���2�Μ4A3���'�}Q�L���s�P�2ak��y���6gc�+�	ڲ�	36�i�3��ߚ��2�aK�j��(��'-��0������U[Dcm��u��X������h�����Л!ۏ;�^m���ن������n���k�qB_��1)�Aj�0.�Yɝ�3�`�d5�������b;� ׆=ԕ4C�%�8��)f���o��_���m��=g��D?���Ə$wÙ�ZN@+�Bۅ�n
������00�jr�v}�-qoF¯���-B��_\}�2��tZd4��E� ����@��*@�{BR*�[՛�0��JO��)?R�/�|a����3c� �_���c���5#�{?�dM����={���mX��rLTX����R�[ey$͐�$�{c!�hMB7���J�������

�෺�
�.�.߾C'��Vv�v�	=L0����o6��n��@��ʼ�����h|��@�7��&���S�o��c`ei��L��n�O%*\6��������q\[>�,Rim������e�����	��FB���呸� �wbea���kH�y�s����s���0B�b���"�{]�{���%��N�HG�Q��NŽ�{������0�<��Ӫ`�┞�:�q��0�Dt��[p��r��6������*��N������
�Ӆ(�I��6�I��T���膇�8�K���4N�Ӽ�Lp�YEl��⪤����j�	>�������h!��" Q���K#g.�;�%S#�a�g1!JB^�<�#Ny��>~;��4�}�KO�"I¹x�9AL�����42v1�p<��	�}�A���癌���b1��}��aQO>�w�Ӧ��!q�#:��q�Tn��  �2���'����P3kL�yaaw�U�/ƛ�,T����r)�2}#�ќ
�cu"�jQ	�qS�� ���s�a/�=U�ͱ�L����3�Gf���Ck����]�*7֩��+;����A��(�ŬWV1 yw���1���՜)���M�����"�kI�ȃ�K^�!H8��c�����tb�;8�
�L�oy���mG���(Ǻ�s\�I�qפi
)�(��wjW�,����Q�.�Tx\S'�\�B��`�����@uj�]��a��.�(����j�t�fA��`����[�w�����W���uǉ#z�8�؁�ڻ���!��X�[���#sK(�tj�)��4�}�d��tM���8�,J�e��mQ{���dK�rK^c��� �R��PؔD88�@��8�j�Oxp���J_![����ok��~p��a���d]����_�d�lń���걝yV�G���z��,�}�$���M���ԧ�Q?V���II/^$y҄$$7zC�o�Pu|�/U�8$E�(p�����]J^,��ӗ5�M9����,L�^�urf��g`l���3	����҄�Q˴9�q���a�.Y��[�䟅�z ���{C�"�����@�ϸ!��#$���+�5ҙ4T�U���s~�J,a��3!:1��z���;��6ۋ��쵰;�7�P���{�+�R�"���<nOMH9g�NX���{!� ��^V ��Y1������э�U��Yd����j�c�Dg��P%�a;�.NQWh��V�s��%�����X.о#����={���e<ļB'N�y��~����F��%qse�n�P�M��Tqmְ��\v�8u3��;	�X�����:6��3B�GW�a?���Kn�
�M�p�R ��ۻ�l�GĦ$Y	�^�+��ɽ�)jG�;q~�;Benw�TŔޗ�1A��g��`�"��͉0"����	痏':��Ob�6��?�晦�H��.4�L�د�E=�A;X�jN�7��z���Y�mMض��9To�����vxhB�fg��С��;VEb�H#��5��o��Æ�"*��N�l"����3��2}Tw�������f�	p`����=��Q�J��h*��'�����\4� �B�T��`QY��7�gŤ��#ϱHح���/���
��	Ү�0V8<G���L�j��8��rM7�UT�u�Poɱ���U����S�_)���o��Yݴ+���(v�7��s��e�׽6�_{����,*�դ�3w����};����� �\�a��	�����W�ǂ������s��o���q�3��VY�dݧ}��ع_�M����=�B�(��XLp�U�Ċ�# C'�B�o�*O����+��S���2B�ZV��w+>�����DKaw�����
��#�#��UWFe_��4�|1�$�d1�HDdU}�=[����@c<�-�
��g���|�8q�M�tB�F�/�m2���mkH��Z}���B S��ul��������+�G�қ���&�Ҡ~���|I¢��#X�l�Av�n�%<��<�òc�ڌ��� ������Q��lB��N�KRņ%�]ݣ����	ScpL&�%��I���*�~��/�Ȅ��ҷ�T��X�������<�orqydZpQ7�~�)AN�x�ܡ�ȃ_�۴������Tp͹��^�3�#����2���ο�w���N�QG���S��/֥t�����B̶��<`b2�9�����;Ƕ�����)�#��oef��NY��tQ]!�������|i[9P.C��<�ڽo7s�?��)����NV��芢�A��g��	T�io���.nq��+	��B��Y4�c���}�D�60#7�!x匔=����ɠ{��q~m�u /��f��e,40���K9X2��r��m��W�,'j����N��\S@ˠ;ۺ�C|���5[0!�f�v�P�.��Gj���F�K'���:�ث|v��>���Px�~��O�K��'�/={G�e?i���w;{x�z��c?�t�L��A�@�������@���	�s���}�$��%�6MJ�_����S��W�u�#����۝��꾼��<�42h'�>/�4R�2*�6�<-�:	�iq���g��͝�_:��dÙ�7�Ht�Ѻ��0�e�g�N��Mi��n�"
;^�F����z�]#�/n��.F\y�a������q����3'xβ;�6��Z�v�ݫ�S[��N�2�f`Δ�#�I���V��eD���L��}N� @\~p���!�Pps W�����Z�R`�������T�9QD��({�"�C8�4LG����2��ԉݧ��d�o�]�*�e4珤�Î��x���\Q�|�|t�g���Z��}Jv"�a��]-1ߡ]��ƛ�Z˟���\P�_�w���"�\�Y�l gD��w*��Y��z7)���q��K4�"!����Ҵ�*� ��������1LL����IE���'.���S�[�tm��(���#{��7��K}Ex�5%IJ�����ӌ4��o��"�|��V�P|�o�nv.Z��E���-h��K�����s���z�d�{f�s���uh��&����Y+��5VAƝ�n:O?P_���z_#y 3��\�e�K�(�2Ƒ��ҳ�A��Ϝ���6qk����GR`J�>��3�a׻(���P7���t+?�3?��vO3s�l_�h��$ks�/9U�sd�π+~|qS3�3C��LX�a��x��w��A�ҿQ!)L�#-g����j��i+���}f���c��iZ���<��4hO�H���aG�][�6?+ba��K�9I"Oq(��a��0r��������g�_mJB�$#6��I"O�N�D����xi���i����Y���M~�� ����O��k+�8�L����󁰊o����DB�?Y�ɤ:�������F_�Q����T��=�'���y�E�!r�f���o����$=����L�2}�����e]�ހ6+i���Bv�������
Jv^�rҮD��L	�	����&�`Hw����]ִz��� r�au��d�KYz���j6�ɼc�P��򁈾Zc��IÇi�'�Ժ���ԉ2%����y�==�N�j��4!��*M�>�OR�/0��A�(�d�&���I���0#��*��p��Z�CV?yc�Y��9��i�1��xK����Х�hN���rJ���9B������p'�r�^��Ŝ������|B�,OF�,+�����(Ⱦ,gZu�����76�4�<�<a��b�	���P��V�Ҫ4��Yy��d�,�æ��TI�xW�!{rʥ�(�������9����d�������}�+�_|�"��D�7Yٌ�ǯ����WSE=��b�^B���GP�%F�iO�ɲ�cߎG0�8+)z�!G(���PM��f-���A����hk �(.���Ǹ�aVx��C �6���>���?�F����F&�lUkՖ��T�e��^��*�S\J�$�����4;�)� �Z����MX��i\ըˁ�|@�;���n�`�nW�p��0�0����XO��M̢��@2C�:�P�d��i�;H3�P�w�N9W2�$}��Ų��b1ڱ�MntxKt��Ʀ�U�Cٟњ �!턡̌
��d��AV���a�����!E�<������TnIH���}�Nx]��C�	41e�HNŠ����	
)�m�g��~�\��3_�;�_�i���7C� u�����`�oE�>���kd7���1�!M�ȁ�] S��u�jA������r��}ý��E�ԑ<��geL�+�x���y�h:!�r���1��z����zz*��@���_�ׂ�d`��ܰ#�\�ʴ
B�X��{.�{��~��.�a�V�'9kǒ�Dj�a�����0�P�e_5T�`�}?���6���-7�'�=�����[Ź60�n�@ל��;��E�s��@E �'>���#���`h
�B�^p���wu����Tb���I���)�~��V6f@�k�9K���Q���P��Yغd��k���5"��J���q���!��Or��o�
�:����7�H@��xeѿ�� �
�6��P)P��;@������x��^X�F�G�齺���8w�lޗe̮.�!�r������@=���)&�#�FP�m;�K�XB�!�S���$�t�V�?����%��̎�l&6�} ��â����J�� ���+��>���f �>��$��	���_^$�x[���32�&��k�'����D���x�6�5JF9ۡ�֣�P���h����$lo�H�����`4�3e�
g�|X?�nc:��(�;��,�X�/蹋�f����'g7ݹ��C���Bc�TH����c��
��f~#�����xct�Vѥ�]�D�{�~B��z�9~$�LQ��3n���!���Ja>�˕��U�e��N�#��iiԔ���
��8��ƌ�o+^2I�S-�ښ8����-��y��nDֱ�G"�n��&u��Xõ	'��3��p��Q���uK7p!	��(��i�B4i����+qM��ū��
�Q�F�Z�b)L����9�IB%�n���,�����j�:�ʰ��[^%17�v��|맰>H1\Ϯ7�Ol��I�F���њ%B�r��ĸ�$p"�T��ڒZ�S�@;���o�; ���1�=�"}���[���
�Vro�M�9�����%ۄ��G�uj�3�s Jc�E�rLw3���'�x��;W�}_\�pӑ��{��kƀ�HD��1����9F�H��݌���Θ؁�,W��z��Ie*^Z�2��B���H	�t�l��\�8>N�<�aٟc���C�a�Tu�T-X�q���$%�0o_��U�� �44әؾ1Sn�_�.��uL+
�O��m�1Z{��;P�4zhx�ny�I�V�J��=￸��&&i�S	I���lzy���\T@��ca΂�@X�I[�Tj6vG?ٕT����+��4���d��X���=G/*e)RD d�5����<��w& @ ]}" ��)�_��Y$�FH�r?8���a���ė5U�om">�J��h���'Y���}[X�����-��&��U��ɲe`:�����bS�H���4�m$���C���0�yp$�I��"<Y�+��>��OY��%�V΋MK�3ٱk�>��-D��r���z����I5=�~<M�Dac�����c�m����.��u�c�No�-�`��߱�6�	�@�F1+��·?MT���s�J�1��Wmh��-(/@�+��'�~O��Q�}��	�����2I6����Y�<T��^����8Ɣ(����`�h,��\X��U�o+;��@G�Nb���`����߬ЉX5�M�l%
	{><4q~ψ�����:�;<�6"�Ʈ���9�p'��g���dKj�F�)�m�I?�����V�v��(�_
�c۟Gzu�;fq��uq�EY��Ę�F��Aig��;%�B�����{����Ms����%�{I�덟�c����6�ĐAv��-���0qH��Y0�����J�L�=����}��Z>��4��L�]ɛI�I����X��}�Irvq|\  8n��?�Q��-0Ȫ�s���o|�h-a��w7����a0n�ȓ̖�=|^E^���\���v��>U0\ް1-��CB�b��=N�.���!���s�e�-Ȳ��v�Ƞ��)B��d�B��fi`3��w{��jJj)n�|��~�tj�5�� �W��v��t �hc#�tn��K`�'����q4�MFh�K&�(���3�~6?îй�ڢ�����򔏑��?g��1��t�q�t0�0�o���c��cD�գ�,�5�@���)F)������:.����I#��I�t�W#��\�H(	e�f�ä��������4uO��J_=�����U�xF��+�´6�>͛B���}�RLfޛ#DQ�������ռ��^-7nx(���]dv���̃�Y�֩TR������K���>�XŇ�Fn�҃�!�H�d�(�Ӣt�F�����
���l�$Md��t\���1fl�  �o�Q9��G�Ѝ������hm�.$��hF�sq(1S����bq�x�rbHv*���c1��Y����C�\G��o��X��ڣ�U̲*C��m��'5��-n,}	?����pQ^�H�}p��8�*h�S0��;| M����^���t��R����Ŷ�|�=͖@��K�d U:���X��s)d�
�1�� �f��$D���G�]_���SG�6~6��G��#��������
%���s�
�_�a·F��
o=�v5za\Q���y�:j029w�)S4��!��Q�zd�>Al�A�T�v¨zfT��f��@��W7�}<~V!�3)��s���,,�f�o��H�������^���SYQ��R�R���P;HG ����wN��Y�>����ؽ�����m���&��Q�k�5�S��5����oQ��;{��9�� ����4A搓%��$����y�A���b�^0�Q�;K�n�Z�鬉0,��maZ�rA%��σ{Z6HmF%/�7<fNi��@���iُ�VM����˩ʦ��^f�M�`Eܿ�s��a�k��l0[�\��U�>��{C�
�p+m�Y��}�s��Go}�P��e��ۍ�t�"@��j�����_�p��qg3>Q����rB��Z@H.ɑ��-g|��?i�#��W�5"�;w�ե"�خ,�(ރ:���=hvN�>��b�[�Bc}@Qb�^�;�p�V��#���9�5�H{�Wb��,�8T���>�E�����ئ��\��k�g7�?��].GO��h��񱻳o�m�=~Lf>:�r�f�Pnk�=�W{�o���K�ڷ�oz����k�X�ք�"7y��ru�A���?����[��7��O{���W�V������R�{2Pl�A`۞�;�n�9�t�Z=�s'1�;+�p*5͞����!˗0�}*X���6�|�	�44���
[j�GS��]#�����]����a��s�7�5_،]݇��F�9�'��_z�^X@k����B�7r_��e��,G�hb↞�� >Gy
�&� :*�EZ�qA���
a��\�`��/B�>�	j�~��\p��v�����c���WgY�����y@�>m�6����Kz��M�y2Ә������t�r<�st�� Z�����&.�m��%��B�^KҒ�f��߄�l>�D�����K~=^��B-9<�$~�$��N%݉�Ϣx��Ra��C�;��M���d�OX�z�7&N��y�a��d����+�OϠ�BuPto���f�H'	�g�Yg������F�^��렿n�v�e������*r���]��`i���`7z~M��p���&e��J� �z�$b���SGi������'^���r
�iǲY-������Z���I	���ni����X4�B!,zo���܉�@�	�խ�!��N>c�^_�9�
4K^C��<ix݈�[�V ����p�̢>�D�dr%��u|�f���q�e�°6l��a����Y��-�j,U�X(s:+I�r�B��E�Y��g�?��kSR��a��N���p��i�@��,�x��,S��R���F��i�D�\��
o8��S;^H��j��,$�O-ʽ�a�- E��Z�v���L���0�\<�1�\�u(P9*����haD_؁���w��'�$.�m�.q���5aGd*p����4&��p�Ba����o��)���YP�[_h�by>��3��a\�� m�d#L
~�):tgk5��B�0=�����O��lS�SAO��e�p�Éj)u��-�Y3x��c�
�!n����ɂ9lګ�R۱�j�_�?!����7�Tf%@X��[�A���R� |5����gF	��c�X��1�Z�ܸ�roOU��Y�tQ�m���b)Ἔ�����"ܑ��z#5��v���7��S�W�� �!Sd/ݱ��_!T��xFd9`��e�[��u�ӗ�6f몭?QNE����,M�;T�]��7�ybVr}�Vq��Ka� ����E��vt�+o�a5;��H���M����F>X=�w��Z�<���ł�0|x(�?�Ͽzs�����q�ܛz�E�] W'�j�#8Q'�Og�q��7ټ�t�� ��މ�ص8�^mUU���	̻�~��ۇN�/P˿���>]����=���u����Z��kri ��C����(վװc{ƛj�׫�O`Aw��'Ymǭ��B�b�:�\:�z9�F���u|0D��\��Je�dK���D�v���g(܄Dw�I#�y��[���_|�'@��=����S+�����S�^�i�z2̱�
#�'hw���ř(�qXL`Bw��J=}ǻ�� Hwĝ���b��Q�f�C�_ש��n(2�g��~wԉ�y��n4p�K��SgF�[��1R9�W��k�ͫ��	rñe/�0�bV	�x�p�		�Z���}��ʏ�7D�<&����3�$fYZu%�<[�������]�!(�3�B�mC`k_�_�6\'-#<T1?�Ip_؀k��&��=��d��W��-��*�:��t����g��FJ��c�~�F$�����Y��W�6P	Pp^ݥ�c�3J@eǿ@3x|�w����ru��M��<�U�s=H�z_�>3��a��W�$!�#'56`�Gr����{M�T�O+Q�	�Ȣ{lA�����s��;sD+�R-���<�#�a�U����##9BMQ�%p<p�rG���{݈ o��'�������¬�:eQ,��72��8�=$Rg�d
�=�f_}�a�Yk�/�j�z�kev�߿+O 5�RV�n߱7{U�b��Nt��������ۚ�]�Z=bv�t�Y#c�Y����[V���� }����V	Y�<x�t��KkYc )�}�GP��nM'���;��>J{]{|��|K�N�̌~&��ِI�,<�i�&*b��H`�B�hn�W�$��Q�P<_	�=�q?JU��Ɉ��'�-��:0�ĘҰJ�I��}�Q.�c	�8�l���Ln&2���yN��OԞ?ߋ�-����>σ�V�@!}	�N`��١�n���$�{Yk�ȍ��	/\8���pL����h����E`;���V�5�%�F%�;#��m`���]jk4v��!��:�A�ot�*����a��;�G��0Y�x��4��bj�7 O ��Ck���-��]"��x�W��&��W��@]C�Y��1j�o9}FN�`R�ۀvr�N/��2H1�f��,����F�Z���}�
3�N��q��%q��j�P���'�����I���ع%����Kg|^"sA.���M�A]r�yY<{a�Rj� ��Y�'����Qp}a{f�v��.�R�xx�>��V��K��A���c.�u��u$VSӕZ�x^��2�;�h�����C*fF)F��Υ��h�R;D�17O��&��3�m4��x6fI0��̈�|Z<�����:j����:d���_
Q?���ӽz��4,o��а�a۩�wX �8:�^c*:����_�����u�	t}� nx﹊L(�����&�-��q7�
���Љw0�oo�oD����J��r�nށ��v�-�́�7����ͳޟ�[i�Ia�!��iָՈcoX!������2��o��GȈ�e���/Q��t��7�Ǖ�]���?�9�� *����c�J��I?-����:�R-Ġ-����6;�@��*m�V�"���������W�}�De��W�[���f3Ǚ�T�����p��86J�;Ⱥx<S:��xu���~2ySC7/��X��,�d��P�g�$�'�M�l/�`�B_�S.�r,��B��c��`��/V�����a�s�W�i&O¬�=CL����|Vf�7���q���j��q4y�P�{�Į}�cf���	`^jn����$%�<Œ�?8�=�j
.H�K��#�LE���"��U"9�)�h���V�A�դ��ܫ���oJj
��`R:���@�%�T�73D��� �e��=}C#
pg:\����3��|��p�������)'�q�TG~����@%�"���(��i�k}��(5��h�	^T���T]�?y$v���B׏bԧL������5_�e�@
�ӂ#츆:��ɑ����`�оns����r&^ J����a�#�v�� ��iD �XkK���a-%�0��Q� ���/qY���+kС�$��#d�ԚW�r�и��ll �~��� V4<+q�ߌc�L�HϚ�������9�������I������ɢ�N�~ϲdj�[���Ø���[4�V��ܦ�mά��6�_���>Rꍽ���޷zW��mc�#��U����}�����qڃ�ʯ�P/M�Wd�GV�<P'�^l�OumD���0L4�I�|���WY'�>ö0GX �!�h����D���!�z� �u��N��e�ZE����&&�V{[5�k������o�2��R���Hb���N,�{��r4����>G��V!���o�8�4�HA�jb���hy�ϭp.��:��y9�D!g�:{�Ϟ�ۍd���pE�nX7ح��f�B�K9�4U>O����
Z�vZ@���`A��p�K�j� �-d�u���A^�L/�-�>��M�+��r�#�*F#���<��QH+jF�ɋy�Q:�o�
㇭C�0é���]C�F8���5E�gX_K�wv9`uW��^�޲�4�S+$�1_?�_��gJ$�̬��#��m���[�-�8����,��"�����	����͊d�"y��}�x� A�=3���ݝKfai�b
tc��t��Z��_�Kj�9Q��q�FƩp�mp��rB�>��jK��N4.�.w�����K�ٰ��|�T���Ɍ-����cYG~�!rx����ȃ2�:�tU�(=��Y��;�?��jC~���k*!�=�W'n����wt��u��!&���/�����;޷�M���4��p��e���z�,S��M96^_���q�9Z[�?�������u�0g�MB%��u�tPt����\,=��zQ�?�2UO��"��J�)zf���x��"�����T�:��h��x�k8���2�Hm�s�I�3�G����ĹYj�";�q}����\���^z�(2eK�I5�߲Uإ@�z�R��S�������*���(�2�@�+���N�����[� hҚ�\�+��ěWذl��Q+�$A���!ᇌY��{c�N��:��FD(��f�S	�W�h�rE�A@�.-=I�aV��x�.7�*�ey���KQ-!��)_��9B��%�G-������ir�j�l�`�М�k��g��U�<�ρ��cz'�q�|:�g ���1�v�6-���L�ε��q�Ff����z>.��W)v'dg���
`תּ��ȐZ�%��'�'�a�i�ȞE �|���ټ��]j��F_�r�ܢ�]�\�O��J}<�C�������9�r�
���rc]��w�����%��>	RL���_St��������������7{g_B�R��v�Z�P��kǹ���֥,�gXx���a}F'��d�Oc�e�
�c6n|/-JW�͔�b�S�*`3
��8+A����	�4��,��� ͎	Fl��P����B�Z��l���WK�?>���zi� UrY��.�����d�`$^^;b1ң ��6�q�@C�7t>h�s�٪�i�mNT��3��hW嬩�R7HD���9�r�M�ߒ��'�������*�u�k��!8������U.hOd�9R�IO�~@���^�*U�9K<�{� �7%��D�m���[��Ъ�F<�
N�7���8Ŧpfv�����%�p�b�|ۏW�|jh��j֐a���:�Zw� tT��}�[f�(�є.
���w/� �WN6"�d#A�P�����_M�[Q0@��YթI����Z&(���uN�]A�{�g�/�W1��u��{	�0�C~]u:�
���!��͏~�n�"�H�B�6T�F�-W'���K�v�(ʀVˮ��0�.Mn�7]��~0��Ē��8��]5�y�ا�jS2��փ��mbt�Rd��vE�4���L�5���V�,z��<��i��ukL��*�6�I��V^����H�~
��f�Ǡռ9P=�"n�-���������Ц/�w�'��*��%�( � �����ΙJ�����T�;e�=�w��W���J��i�q�
��	Z�e����$�iR5��LY�SA����.���OO�P�h�.��Jp�_��CKW�1��z��N��)��$n��çK���Gj�ZA�G�]3C�ikp�[����Ȱ�#?��WJ��`?v�R�yO�Qa.[���#`�@�5R�D����}%%A��m�q!��l��{!n5ؼ����\{1����'Gy�ə�?��Ǳq.�\�ֵh�Nq�P)�l{�X[��p:ȥԴ��qft^W�2�8�c%Kj�,�2�~�E��*��-z��'s�C�보����g�N��u�سz�'ڢ>��G�ga�H�?�.aR������liJ-���<�S�?�����l��C�ۙ��~�@-u� � Mǆ�6)����9!
�V7�LŞ|�C�A����������E��s�n��?80�-�;��7����[X�y�W�ֆ�Wlh�n�S�p}a����k�Y0j�^xL�4���\4gϊ�����A�?����
|�{.���s�<�؝(��+��C;����T�m�bE��z*[w�ԋ�j(�l�Ac1�#��"-Gy=$ٮ%^E��a��Q�8�\�в�������	<({�<dއ�1.�߉Ul�y+
�)���kK�����e����1�������s���{	�K�����uH����$�FH��oa��QCL\z4 П��uq��}(nD�)�W��zm�S"�gg�G�������e� ��ѻuA*�x��R�+U/�O۽ɠ�"d�眶�g&���q*��'�GA�:K��%�*���\�����^�o'�F����I��1!\M(�O����#��R8;Ts9K�QXeg�� L��yU#��`p�y��*��~��Ý���zS���be��5-�6,����Ƒ^(y�I�1 �l���ߣ�������s3m��/{��4FxT.��¯1��̜ϡiȓ�W�����!�V�L��l��2�Muj����ْ'ǒFG�xe�%
"Y��r4h.�U4o��t8���7�VK�<�i\������eQ�z�o(#bUk�3�o���Hu�(���r���#��#c��^�+��}�lv��b/��'�Aw��X(��	�z<�.#H��.��8l�-�¿��!V
�)�"��g��5��4���ُ�+O���f�����{p�TT8�c,���cIQ��U��/f=O�unٽo�X�\�?���/!�����,�7@��n��Ȁdu����[�+�s���$�Anp��|��Q>��ῂw)��x�ۜ��.�@k6�η��9Q)��ӧ�B��9�HP��y��/؍�8W�9�n7@Q�1^�L�p�˹x�a,����c���L�J�8��JL�� ���0ؿ��<�qo�K(�X�ì��b���t��\?y5mH(n���K�;\L���ac��jںy_�:�������˳̽EmO}�\�����NQ��`u.��#6��i,D.��35%K��l���7�!�h_:����O?�,���5Nh�`�`|A�G�:<�	X���u�v��Ϝ�<"�����F�W��Ԩ����Gd�F`�	�ܽCE�&�Zj'?ҔtQ�dZ�e轌�� F[bt�߲쬫F֤��X+YX���B�a��0��Z*@�#K3��q�?ɋh*6��KP0��
J@�A�� -+�f�����lB�Cl�l� :�S��[vzP�5��ɋ[�������n�
a�l˼��=S�s��-/<����۳�:G� X<F�����4N�
xx���O�B���ՙβ�el�b'/u�u��8��M$�		��l��:�w���������F��@�W��t������A^ث=��η����Uy5���jލ�Ĝ]we�ˎ�d� �Ȁ��w#�UI\�b�ʤ�ˣX; ������9���cxWl��N: ��� ��5��K��P���6���{?��߭�lP��\t��<�췱*� 9�d* ��Y~�9U� �X~ZQd@������s������ec�[�����鏙O��k~}Q�]O5#���L�R���m�Z&b���VZdg�~�B��!�g�8���c���$a�τ�d��qk�l��F�dO-�{_��o�aO�K�6D����Ҁ��/8O
E�]
�K�i2oX�9�t�:A�2]>�Zl�*_��r�����ޤ���-p �D:cY�i���l�=��Z�w��|�.������cԃ�[�:��L"�"&���W揜���@Bf�FQ�.��Ě
������p�[���3Y��mfQ�������a�e/JC�G@X=�;異�x�껶�bY�~��=��$R=���b��g/P>�mC�������N�x`]X�G��T=j�	�?��5m�k��J|����u��3���>uғF����1��<]����]�ї�ǻ���q�����tE�Mm����Ⱥ��iyimX�M:��7g�%l�s��s�Y��o=�v4@�L��~����� 1��*��3���3O��%A�%*�Q�UR�� ��%��`^���7w���(��=��Bt��m}�unR�!��˅�����M]]�)��������	�����c�v �I,�F2jQQ�O���m3jկ���>���q�*D!�Z�K�@�K����.q��x\܃�˘c��ur�Fi�+=���
 �G竪ͧ�o�狞��B������ܼ\����K(�A�'��It��t�'�l�8w�;�x���6Ø��"+�Y�0����@t��I�x�@@[?VW]�z��Uf4y�a�J�C|| ��)Y�ݤ��-N�E�3v?
D�h޲wS�I&n��D����v���eI�!��^+�,�Fۍ�Q��a<Vx����U�g����{��W�bZ^{=��6v�/��/�+DU��8�����x�O��O8�f����/R�4$�O~�K���)�P��a];)!-����15�J�#6�S6�Z�QzG�E�t���/�cY6OKxw�
��.[�I�B�rƘc��}��{�/��:�8��7X�i��p��~�b�ӵ�1�;�]F!LͿ��ʌ=��J������f@�jgLFG�����'$���_����Y�e/�,��"@{5Ee M�TGxͥ�d|���[yIk�/��uW¥�J1�<QY����3��\:W�-�\/����n�ȹ����&��/��R���Zu�X,�s$�eL�@�Ei|0J�(�YCd��-v���56s-i�ּ�����k����%����?-m��?�Z����ZVpo@XO���	y���������e��M|BF���r��Ɵ��8H�Ɯ\��>ՙ{e>~	��h���._[��;�J;��#K���p ���|4]~ ��I%ܚ�4S��馓/���K��"O`\�SS���*;+!8�#��p���6�
z�FS�)=v i�`��a�L����(�G?���=���%,$���'YR��B��;��>g���5�KZ{��>�U����2�P ��"����SV�mR(�gπ�$v�����weQ��کG4���
$1[_e�kȂ���ߜ�I��_4��_��Q�{|��7kp��^�وC��Vܒ�]�J�/��Ȋ��'�v��o_����Sj�O�k��Dg6����[B��6�jMƥ��Y֍W�٢a��J���C��n��ii�z�+��d(.�'>�Ǟ����{��0Ǩe����nD�h�MƐ�Zdj۔U��ր�"yS�kr�u�N���M�]��e���SP�x@6�!��M���+G��Y�(��t��l��:��[��0�i$��7_@���Rۉ��NK߀���#Ж���2��֘�2���b�=��4�����s�'��P�n��jj<�C���}!�2s�E(��	�LǷB�"Lo�6=��\GG�A�-������q�H& {�ؘ�8e��v�[˜��H���綎S@���3� ]_v��Y�U�x��'cӊ�8�'����;���,�ۣ��@B��$Vq�"#"�%ΖS�)��pz��oA�Z��)��H)��a��%�h�����d~�\���c���9q9�����RbM��d�M�Iz�HM�:{��^%�W�f�IbXcK������=�z"�B��´��z��5���I=54��[/��.�ޫН��
S�K�B�Ru���d(�W��mB?��-7OD���~&U��u!��p��xJ��g�La[D)�o_dG�눣G{����*;���RP}R`Қ�7�����"Wuh3�2S�8�@Y��g�����T���x��뷜�z��`O0����o�I���k;�^��֯�U˅׏�<���&-�:����`��
:ϱ��Q��b"3�c7�N!e��K5b�o^)&n�n;�������3X_�\81��^�=l�����)P֣M���٥f\�Um\�iZ��켢�j��Nw�	_�+�ɮi@� J��ۯ���׎R�Av?y��Rf��xMXj���Q\#+i4�r_5�F�:�Od��is����)�۶^�]̜�Q��w�Ү��(�r���X�%9׭e����_K�R
!L��2�1���P 4���8�w"�GB�$+��my;��[�	{��E���A����&�K�M����;��[��W���ed���@{7�=Y0��:v�Y!L-���ݭ[<��Ƶ�����ӽ��ؘ���ľ�ի��p�IM�0e�)Ӽ&?[F��FIw��]ּ���.�R���Ӎ¬>a�03�r��`D`�G!�?A���Vp��ܢW��D���ܢGpL���	Y5�a$Ȗf3�󰞈��6���%���!f�	�y�kG�po�6i�2��c������/�d�f���5߬��V������A�k��H��Z@k%�"ÉA���p���"����]ki����ґ|�NH�}�5�.ZD�f#@)����DIA�X���|��v�\��	&��!�d�;����^�^���@�3�
�>bmnq^�:�`�?��$_�M�X���r%�pZ��1f���q�݉�۽J ��8T�(x��Ӎ�p1�"}���p�N�d������meCsK�1u�*�<��-���6�5,'���Xe��ŁLW̫�A�0Z���V�D�\��
�dc��Χ��Z�����?ނ^dy�|��b��z� 0�����Q����TjH�f�R�B��de�o�PM����2�!�֨w���(�%��0r�@�.���$p仢��>�9jՊ������ՅGT
����,q�U�����PM�G8Al����)�b�r�e�}�@ӎ,S���p=�C8�Y�u�W*u2"�Ҷ�n^�v�'��.uVz�B��zN6q�Frg��2&rvB�_
������O�������/�W|W$�M� �'�������9oX8){��<-�h}�#�����[^�B�~H��s*. ��(Ǫw�A5TU�D|�'�������jԟ�ӆ���߇��!��c(�Ή�"Yq�W�����<A��K71�y��V�d��H�.������:�֢�N�9�:����p�Mj��X(�e�@j�hon�p��c�+/�d��>�'������̷���]'=𻃠z�OW�R؂��yAi�G��r_�cJ�z�M��_���mF3Q����,B	ݔ�Vn_0��x�x����M��� ��@P� X̶fm���7�7�e|Ǒ�k���\�|�U+��^�٥�a9H�/b���Nąm�C�ȹM���8�׶��|��7໫b�@�y2���ǺN��`��fD�#�'r"��`��KLi�0�b�{->�\�T�-��{e����[�[����0 ��S�ʢ��_æ����A��b�2���\������qA��+�{te2b��s�I�Ӣ떉Ztw1P��	Z���$�jݬu	9����t�b�hj��T�����%QW�F\����Ŀ܎�5ӏB4WN��D�{(����u4e�<��a7�_�ѡW嶃��D�0��d�/�KjC�_uOW�˛�S}��$���zS]�4R�,<�*"N�gTw�ø�f3�F�ju�	-J!��zy�c����
U?�j_��fF;�˪U���I�
�b_��D�l�#�[-�����9����&���xb�xT��⍔[�kK-��&Ґa�ۖ�+�2J�3<��Ax��{1\���py����F*�����}����+��z���$����4F妃8�"	��h�p�\��h���=��$�&���MPv,*C���z~�@�m����D��}��V���]�rZVߑ8����Zv��E��dD>�S�v�P(cYX��Q^�� �uQ������&ϳ��`�q&�^V_hP#{���lB�	kk7�,����:�gԙ�cA,��;�Q���=������ �c���=��9(b�5"�z����8�(���lZP�Cհ1'b/�?�����t�&�%Bw�ύ	�:��Z��?]sd��� 6h0�z#d�WgC�L�O�G�}E�EOJ�܍6�fl�Nvo�2{D�<�,h!m-�Wl��>3��4fp���{X�0�T��X��J��^���d�0�N1�㿢�W�Y[�~8��o6�|�j���\�|����砗�ɇ�/̥�������ꦘi�gm,$�rf�"��W7_,�H���p����GF�z���^p�vx��^6=o��B骔(��k��qBq>�C��iEJ1�N� �D/���ßN�2�2�F��'���J��$���W���h݃1[�$!�{W�Β�2~K1�`�u��cn�[��	lfѽ�Mޞ��q���L��x���w���h��ׯ��(�/��X#���������h]��;���������
�?�O~�{n���O�U>��Zv���3i��M��H�oG�����n%�nKO�%�Ep'(s><!�|�'�?e�IRz89(Fw/�S4'�Lo$;������X��$�����Ҝ�H�XelL9�o{�ʶ�.��Wy?� �l��OFd��Z8�E��F;�3�R�Uq�͐��� +y�+�h�����9%��1s����v�LT7L��o��'�w�����@��zTas��1��]��wý�s���z�ŝ���ͩaW'B��L����)\�--�ҥ>�e�[�@,�2��1#��� ��ʊ�K�����0߾�_�Yu2��tT-Y��k�+?�͗��5����԰���,���'�!�IX���A�5稰<��Hclm�m`��u��.y�Ѡ��RH�e۟����V��U2�9m���e������q44���#�D1_�2��K���CAXL���E���<+|[R�.@)k!"hoU�\���t-44��s	3�j�Qsݳ��ʻ��83�2�(6qOe��H���z��RY!�V�𮌮��k���w؅��OJ��dn�ص볈�s�9� v��QPQ$�HK�>���g�' �����K�0�BT����ݸp ����8<�F�s�
��_Ne9�q~_W±����O�oi��;�%/��.2���UTt$�����,b��_ٖ��TȈ�&�����p�86!P���k
;aVܠ��n��a.z�8�S�t�|&�چ�@y<�\�wT��5-���d�glu%�]��E�VS��Ovz�D�)�:�����nH&�)}�	���7�hF�a��-�2�TF�Li����'�eK��{v�a��n9��G��ġ1]����:5^��Un�:��H�S��@����J��V ���0���l\;$�E"<���|����{X�Q�3��5k>\N���Y)h!�z[ڏ�X�D�~�s���iE�N�E��^�flU��N��Zy��s�z�	���te����&��_�|�����@���,P�ċ[�ƟgU�Sܺ/��"��|Q��>j���J
V5'g�U�V뵧:�����8�Wj���:�	߷J#��6�,ݘ�hL��1���7�C�5г�A��-٨�[V���h3��4�8W�'�Z��h����� ә��T�xU�W��p�}b��n2��(E�P5 ?��2{\�Sw�,X�a�E���y����D2f���8y^�MP��ʎ�*CC�_����X���c� �~��ܕr�	�dxLc ^]�Њ)�d���ga�b�!Ή���#���`H(]d߱a�.��c�|z�G'L�a��AE�d.M�����XqI~iXA��x���U�(%;�@�bh��z7c��#�&���׸v�\�;{F�4>ɱ׼?X`���ۍ�կ��W{��U]}�Fs���nq���eYTOk!ĸ����ˍ�Xs��_���϶���~ڮu"�:`s��yN����5���.� ������괾s,�e�9<i��+�>���x�G�����86H%:�`T �O����,7��(��k���pG�%HqI~k��	�9�A�/"C˝ĦI�r���,�pƘft�a�h�W�\t4(�Zf�>�VD_J8
�]����}E�i��sԵ|�I5�\�������ϡ���+�wۂ�h���+s�G�;�ﬞ`.ή�
�9V���Z��S�����A`Է�<�~��;e6�;(A���`5���^�R��t��I*����6���� �^�C�Q�sC�r�Rj˒a��D��Y�H�v�� �VӨB��:K�/�f����f�қ�HW�B�L���t�SLJN�co�
b_ER�}�){��Ss.��E{��/�bA��?���gq�%�޾���:�+߉0��ߙڎ�Q������T�"o]W�Bx ��O��e�>�*sL%�o3Mz�8��yJ�L�y����%�	Kq%K�K\2߱��q�W�	g(a��&�NC��\<˭0��[f)���0���Eo�JK�4�1��k8�y_���ŇNHu�g%��u���6��6D�O��)u�W&�Ȁ-a5L}�=�>'��^�\�����28�f�2bQYQtKo4������y��[}	�V�q�CRH�5XF�����h���$Ʌ��f��1���*�$��e�U<��V�p����!�ȝ=a�~l(�x�} ��;UY��eB�DPUR4?�����sy�:���o���ʽS���we2�K��$��j��b���j/м��|A�����Y�-t�EX:����a� )n�,$�0��	�CM�v�S�)f	Ñ)���A���AԂ,L�I�-w�@� �j�I�%Zt����_����#�q��kB!��G��IJBO��=�N��zd�XYq���{�*�BS�6���������{; �R�ʌ��]w+Yg��	�V�#wK���b� D�Y��]f�e��O�i�i���\����&��_]��.��w�0w��&����TD�E���0[�/�ج�Y�!XV���x��P��lˮכ#�KHNg�o�[�	��2�h�8��]���J-�Ǭ&sC����N�R@ �WF~��#
�% UC"1����z��^AXHz]Tf@^h4=ACuR��Mk�����>�{�¼��!4��5�X�{'�(z�O�ؼ��-j�19�$��wŀݤ��eY�-�?�Q>\�d���x`����%~�玛�n
3"1�]+u��T�5��ה�y&�A]�CM�~�{����La͉�����~W�v5�	@�r�7t	�Ƨ77R�������Pd��S&��<Ǝ�����Y��s"�����:nRJ�Iބ#Q o��f�^�Z4�o�F!�QD0���ᯐ4+��e!�QT#m��z�#��ΌY���k�ҍ�iQ��RI8�&���/��3R�=|�g�=��les-����.����H>I��A��d�g�}ː���
O����@L>HU�$�!ڹ�)��ۅ�%(9���OʯI	�q�z��\ �Hc8�/˿9����R�Pu6F�1���c����W��>Ȟ�-]�f2���L�Lu +@Q!����k5v��b�_�΄�!�7��t��� ��UZf����.��en�ࢴ�r�����^������k� ��J�c��Ľ<�\��i���r�*0"Z)�Ğ;�������0�㲂��T�zw�1���詶 ���Q�)L̬=����r��}�6E��WR��������-�UXS ~�(RV�u�e�V��-�>Oȗ��$����rry�X?�Fu����I�l;�a1��v<H�/7=7�a��~K��TP����\c�"���#{<���B[��R���0{Ύ�W�~�.)�e�`*��~�j�g�6Om���eEw��Ӗ���LU���^ʭcB����R�8)E�y�&���lg�X򐿨�}Y-��{%]L�4p�#͵�A�Z���yw�M�㻔
D�a�l7�Tz�s��qyA����ǽ�P�_�) x7\���G�2���܃W���0�L	$����s�I��N�o�� �T��Gk|��1|�<�2��`�,�٣V�0Y�K��ݔ$���J�"SL� �!�Gg�\C��>�?���H�
T(z� �"G�1[I,GĮ��鈬'BB�Չ�z���Ճ3�s�}�H�c��<*�Yg�����鑽��*L�"=ɢqK�m7�S�<����2њ���C��3�L�n<e�@��>k��=H�ǫ9��]y�k�`�g9��C>Q�_�� `����B�r=��5�����hl��≯���U�S�Ԩ���,�����X��y9��[�~҆6יWM��?����].d��/��2;���G�4Nz❊� ,�ѫ/g�i�c�q�J��_���liS{L�YƲ�Y��0��&�<��P�E{��8�6r��	�
O���)@��Xp#3TJҘSy�]��ފ����MU����K��`�3�yr ���GLʤ,���[k�w���x���*
3����!N��#W��.���4��V(U*���4K[!%��2��`-
d�D8�ҩ�'Ϫ�����!���B2 ��G��\
+�x�(�W+۟�8�|�^.����@L(�%������M�@
��D�*�~Sɝi
6O����r3��A�$M�uy�������EK Pğ0(�u ]}UG��9�^Av2f<�C=$����=��3�iv9qa%�Pg������wcA�J�D�Mb�(��*�S��?��x�/V�xۥSV$�I@���UԱG	�&i��|aS?j�c��$Kr|:��\g�E�j`�\@�.��n�#�Q<�gy��ռ��߻�t��F���l�>�!e a0��:̅2F_z��M���5�l���U��)G�`�
~ɒ,������fѵ�����ͮ86]����o=��I�L��4^�[��J}�6Id��C4ȿy*�2��w+�s��Rp��-��ڠ���YaG�U��.1b7��8""��	Ք�����\J��G)Y�`!9;����#�h����{��Aū����b��Nb(��1KO�����V�G�>�g�	���yG�Ŵ�5KV��f�0���os����q:A+���׀/kO���j�N_X�b�D>7�v�s������M�v�O�)��f��t�F��*��M��o���Iy7�j���@�ި�:�pW�~��ie����b�0$��~��z��M����0����y���yM���-B�<A<���w�p�'oÏ1�"�Ɍ�Y�q����kO}C$�k2��n�NC�Ѯ2��qf���i���k��7 ��X��Hb~�y�����\<��� �Z�k���u
X���51A�#�}g�x��V�_�5��x�Q��@�)c�ј��M���C��z�aZ��S�x���>�֨�P�����/Fـ�n��W]j���s�&�����TZB[��,�A�4�AYН���odZ�o�҄ț���{)�8�ʬ�6�)�X�3ou\�[W���ˌ'��5!t� v쥻�����F�u�׭��E��`	��/p4��fil�Y�K^&C\�ɟ�wŰ�r�e�`�ń�Y�����}���=��@��A�ŦY��=l\�bR͂�/��>�=� �՗&}@~t��[���d�3BW�Q�xـ�!	,F��W�CSO��,�X��k���[��F�%w���̒����K�)xau�B�y���0������ONf/�� 7Rć�ݑ�4��s#G��� n��B2�L3ɓz�dr3�:�:n�b.�Sr���)Z i����L��t�ŷ�s�r��@�#F����+�)�akS|r@����
�3��*p��vY ��f���H?�����˕+6�S:�m�2!օK��6g!���H��E���\ز!gd� 0�b�SGsA�k���
X����۫z!��S��a�8���:uqN���B�æ���hJ��Z�h�(�'�@g>���h��^&��m@L��k�	��3��q�xo�%	$QjX^�6?�co���fut���s�n�>h�d[������4n�����F��?�R}�j,p�&��)66�#�X�����\�e���U-ǂoW����>�A0֖2�n��[���Pe"&$���b����|qx2��{�I�޺A����˔�M������]#VFF�j3�cG'�[W�����L�$�#������3���G�՛[����ޗw���0D�70t�s�B��{̔�+i-�q�nh�z^>tN��qS_6�Q�֖Ljw���@�o,y���v�	�?�/Ŷ�@�<W5�����X��[�;���gFʜҜ�[�@�Yf �n �� 

Wp(�=ԝwOEQ���SLD��5����'S��V?��ِ��	� k)6��4`.y7Iͯ�;m?��bo��Aq�؏&D�-"ҎE#�=X��E�M�{�[V��[�Lj�ҭ����<�"��/���(��i�C��:�7�@+��ѹ���`�9�C Z���� �6C�Q�a4sZ�L:�A���L��A��k�Η������zӪ�κu6!��
�N��S3�x�计�]XUh��n��H�����.��t���|d�1C�w͐^�nמ��C��84cV��������4�\�Z�n�9�?a��Ք"M�k\qwnOI:�Z6&$`=�Lm����1����WcE��s�M(J�41�bI**>7u��9�kMR⧼`�$
��i��R2��Yնnv̹RLT��tQ����"��&��
�q�.�A�NÕvj��f����GE�,���JQ�R ����������m�E�[�'��sR�^̱�"�c*Z�*�Tp|$���,	[�<LiD?�8�	�t墷e<�#����=���[��������F�1��춧SO�:�r}����Ms��Q���u�~�uS��
inz�f�I��n�3q�t[A�YS�k}A)������/��E��> Ӷ�X�9�3��� ���ݖ�}�=Bԗv-Z��ϱă�jN4�N�E$�y.�S��'M:��u"��H2�V6�^
�b�_�Rg���h�����+�sWΔo �%T 6E�l�sM�-�s��z����{"�n����fN���FeE�M�+b���N�=��7�Z�kB�^al�ȗ2[�C�� -<X$��G�$�1-w߁��� �ތC�N�gV�?#މ#�3�Wp,�~��:1�+�N��DR2�Wqz�b㒔�Q����`�L�=���:�j��qmyEԗ���(up .�R��x�[Iƺ	�p1���DLu��U�v����{����d��f��pyxͅA��
`�JXy	%)�M��-7z)��l�cR��\3�u���oӬ����Q�F�_��t��5Ut�W*��P
��QP~N��|T�K=p>e���*�n;�'��,�]5{T00��yQl��w��-�k�����-a�=�����Q�E����Wk�eX%�S\��K�x�d}�	���~jV>���܆��� `N:�qC"����H��a��u��V1
�5y�5ר�@�o�r��?ڣK<-���cp*˗�K��u?dh��	Ʀ	)yi�,�m�*���X�Z
dH|��e�{=���#�+�ǟ�	�����"�џY�l"��$vd���&A-kA�j�q�eN�y���Kn*Vۨ.Y(���='��}g�[~pH!C��9$B8�ʢUB<�QubW'Ҕ`!�I��`�_��f���g�?[���5%�7��gr�}�:k� ����oH�mp�k[R��[ 7��\�A�'/�&t�)�"E<8��0*��r&<&\��x,�m�Y�<,����]�����<�4��)�C��R�U*�k�#B3B���d�=�hX0�&�Ost4�4Ol�/��@0DL$`��r���>�.=��8�E�1'�м�X�5��g�a�Y2Md�S�/M�`<�pX�bVqg���v�����B3�o�(�R�-�p	�f9����B�������grܸ�a3�eZ���� �(�a�|�������.�](E5)��5`�4��bO4q=SJ���`
� ^� O��yv�࡜b'd���Sg��н��O�Mr��������9�0Y�d�n�Uی�]&�7�s9�$�rS{1��R���t�8J�9lOa������Nm�[�%	<s���Q���
 x�-�||��Vw�R���{o�P�U��H'zQ��0<���$|0ö�K#p�UH�]�A��ELRH�?ܗ���M�J���-U�sӿ|��]��]�^��%I��N�Z��Npof���k�,(���,��6�`�a"���Y�>���+۲���Ύ+�ؚ)��g�ع���P��s�}�X|Q��m�[d��M����B�wx�b*c�f�Z�D4�8�=��	���˰�_�C�z7rܬ�X�&7�m�FX��a�OÇ��xD����b���2�j ߄��'{L��
N������=�	�ŰvH�e�I��Ӡ��UeIe5jz��Nchˏ/�SV�]_ ��C�$��7U�������b=�SU0j�5��z�@	zX���S7q,��搋�����K���F�W�_}�1�E;q���VW̺�wMY��H��/yD1z ?�-/�]��fv^H�ɍ���2��[�p�}fw(��U#>���l+�HN:��\���A l�O��G֡��3�q�V{eW�1���)A��j~i��V�,��&J�ׇK[O1���9���ݥ�
}*�4e����8���?� �	���w<3A ��`�u��;:
$���8��#��k\�h`CI24x�$�W͟?xvv�I����s�l*#�
�� M�­\��2
s#)��0�T�n�;Z8|��Α�6S �R!��ô6�>����2��� ��d$�%�5^�'�����X��z�	��X�xdu�AR��}���{�X�7Q��A����SV@#����ڋc�;�G���	"�v�/W�Xv�μ}yֈ�e�!�Q�l��mh�#�]>��/~Ҩ��a��� ����l�f���N����0��\�H?s��$k^��M%5Y���u���Z&b�a��D�K�2�̕'J��h�O%��bU�Ӫ�8��SP�72[�X�������(|�JMP�h���	��!^9��Z��%�l,f�z��p�́�nd�|�S��p�p���k�ը�����%`�R^������į���5��\���	�7r�*Ba�)��C��1��n4��?N�s:�]�:¬�(�"��b�D����,���J!��t� ʍ���_u�/p�
�g"��ˣNu�������Q��>CJ�h�d���o
��Y���)- WҲ�+���5���Wn#Ru?Ь��x W.)#��0������D�23#����9k�G|�?�R�t6��3�m��3��+9��ңs2UL��>)���<*��2� m#��2HI��e���) ���� (�/��	S�c����:��C��	�P�![���<<L�֝~O@G���pS��yL�o�R
nB#s��'_-_�}�"/��Y��)Y�r̯�Z�Jކ�ޡh�F����MӺ=������o���ǜn(�U�pM����zs���*��d�p��o�Ѥ7��Y�lnI��̻�ǘM��R����K�7���i�  ���J����I,�=�#�@�:?j�^}�m��3�g���$�|j�X\j��
G��!�%>Q����=��w�t�%&'�n�s;s�>��,d�8��4g�s>[�ي�~�M��Pn��w�+�ؗ��m}��ir_��U�:?-j�$�)�v���\�Ln�؅)^U(�|���:�EP��P���Y,x�7^�2�VN���gq2=�z%��K��x�󽘑b���Z)�LA	Iv6u�����tfJ��:G�p�4��� g�ؓ���/6� ��%	��N~�N�UT�+tv�ө��i��B�Sd��m�"U�?����%Vg��Xz��4��+��I��L���L���C*3�ƣvg�j�(,k�tZM�ȲsJ1����"�7��#-�J�4q\y�Um�.���T_v�(�$�(9�KF\=3E`A��	��$��{kV�ҙ^>�i
������h0���r�pco-6��??���>Tb��XD0���7���YQ
{Q��p:nq%ryJK�� ���adq�Ֆxq�QǦ}�f��m9f��>�{9(֘k�����h\��q�������ĦGg�̣z�3y�iu�6�,�j�lC�#�A���)�����y�$<�Q�������k,1�r�]E��?ޯC�cw���}��7w��u̯��Y�f�*�����ި�y]�J|�ׁ��-��v�����W6e�M�4Y/?�D�����&�N��\��Bx�s]J���zX&ð���7��y�*�	����I~h}��o�Ͳ��'Xty�:X�IH.�.^�N�Z���jw�������}6�үhug�ʖ?��SYk&�!+V����_]v�(�.���y]?����V��g��r����9@$�!�t��B��o�E�k�/S���\ ���Q�vr)��1z���l=$�e�n���3:�[�qS�����3a$r�W��Q��� �lk��lp�}��k�Qhؚ	��@�7��q,����/A}*?��ޡ�k�O�� �H.��Ј���q�����t�_y��+��N}�Y�L�
)m}a�p�����x>s�l��n�����Sb��>�r4������׳���᠊K��G���J$b��r]� �.��J5��W���o��9*���ܼ�Y��
���)��.wQ��X"�$�֤�p�~�XZs����k�o�UZ;B]t���Bc͈o�N2L{J� �<��%�r)������"V��.��P��i�c��۸=#�������{U$���\P������p>�%�U&J�)�P������0ý�2�l�s�0-�X*ԧ���}�8ǟd�R�wz�0B�E:P�&�a<��e���Ս<Z�����MђGs��AcѢh�)�������bT���$�K�I�P���G���Y=�}дc؍e��ۺ��dܝ��H|1JKB7�
$jc���Q(�G�˄B	V�]xϿ����� ��h�ӱ����˗ЍB�%8&1��X�)>M}�7�Y�I�1D+��Lj-l����N k��oå�c[vFo\��u��!��2f٭d�L:��,{���ʊ��7�v<�%�N��`�%@�A�h��"c1N9�B��Y�`��R����
Qܶ�}P���ސC�:|��ֺ�\
�;�?ZV�p��1<&��d��C�S����od ���5>���f5GT�(~'|Ӂ΄bR�����Β������	�����3��1�h|�+,��иI���[���x����t��z@��+��׮,�|g�-���E�MeI��}�_Գ�J���c�6hO�����Ny��h,��	4+�L��4��(א���+k�r+debQ%�� ���}��I�El"�4�5����*J����������������1��n��_�V�Aӓ���S���B�:|�s����\!:�墌���X}�1�=8�������ߘ�E�t����`��8Z��c��`���X�u�R2:1�ǝɳ�)�r����Ͷ�Urײ�>�SG��$���W3�^ˎڣ��V,�ў#hT�o	�_j�`��O�����m��=�&6R��/ª�������6�B؀jf�8jë �	����Ӑ�Iy\����"�+s�K0�+>����ˮ#�K��i���ۨ�Ѓ��� 4N���k��Ü�#���U��"�2S8(./������cX�
L�ƅ��ɺ
 @C$�p��WE� =�MMj!�]��m����VU�����d�l5����͗�ܡv��s>��q��t�h��]6E[l�����F������J*G*ړ�mv��������JM�yocX&�r�큧�� �+���W�rDϒ�nv6;Xje��\ղ�C��h7s�=P�/�;�o}�G���Z���!��G��[&���{
|�Kx�_
�� ���
��qbXb�F��4'�v�yt��NG�:�>ι����?!�4u��:�Q>�TB]������,ˋc�{>��d��q��\���d{>2���9a`�y�"��>�ՠ&�x^]x������w	B`�	.�%��$����ɶERq�:@i��Hzk{�(�'J"��]�JѸ%~4�7yQ�s/��pՊ�m�+K���� �\k?<�7�\�9�~s��e��~[:�f��׫�z*�Uqxq�X�����h�ǟ�(HPS��)11����;�Z</v&
��AK�5@Xͫ�ځ@�ݺi�:���~t4��9Ѝ@�4���]�U0s�XsBDR��뿀=w9"D���!Btضp�?E�Rj��C y���{����j+�ru��m���v�~��?F'��#�l�Dͻf����p'��Q�Q�2��z3����8NLdn9
dH�*;�`KZF�F�q�*�h[�A�X=�n`���j��_h�ϩu��+rm}|���M�a̕���)(�X�~�l�ӨdՅ���1��܏�}�;��0�����:^�����`����2��e�]���
E������f˪�W���z;t$���i&V8j�)x.Yob��!���=�X�){�9BB^a>6����B��rx���&�s����՚.�Hj�u`���tîfu�n��Ӵֶ�p`}M�[��st_`�q�%@�9%���a�}P�P((>��K{����
I	�c�W.'0�q�Ag@Dg-��'Ǒ�a��k<����L{��n����	���M��sY�q�����A�J�*$jN�t�Sxd�t��q�{�_k������Ҡq>o���/����[`O*�G�\b&�������+!�M�h8��'��Y�m��a����\�ou�D4�l��#����rdK��'Z?��#BCt�adWS�{ͣ����S�
l��l�,}^R����R����
t/�)�,�Q���W����][�����$y��~���:5�
A���an�)js�d�o�Э&7�%�DR��m�A��}$�*����rz}�d	$:��^�Kp�=2�����8�E�)�@�q�Ds#�S.�%O��ON����)�Q�����{2���6���S��������w�/؈x!�*P�0,���G8U1���m˯M)�9}��v�L�G\ס&v�誺*zу`Q+m=�8d���G_"e�G���K��K���3+�0����I�V� �ʄ(��-���8���b������޹��/�9��s��h��djfQ0ġ�~�0Gg&��.�����9b;|o�G��M߅�@��-�a,�w3������`jS�b�����H,���D�mu\��؇�Og�7�o�.��>\���x�x�+���2�0|��%�;�**�'�O{�Xv�*=݁�S�V�?�Gׅ��<��C��Q�Q�;.��u
Д?��`�. ���<�56����G �56�rR��Y��S�\͇�Y�����}Aa�}H �N�S	����5��I2;ϡ�UY�ާU���\�������0�"Mq�{�,ze5�&��z��I�A���?H�'_��k�aG��f��y���������"���~]�k4�K6Z�S�oa����}BA2kO�T��*�(�pe�����Ez�j���	>���� ň���j-D��]���=_!,��8�s"8�o�����;��E)�S��֣R���۳gӵpJ����3�Mڹ���+y�/�ʡ�� �� v��l�`G�[�-�[�v?r�w(�͕)f	9�6�Ѷl���sLu�pm�En�f�MC&��E����'��CX�n�yr ܒ�X ��{��� �P2�� �\C�̮ȷbw�;���ac���v?�IQb0+��2�/=��8�v�0j�0�$���_�Ê���Dڹ��M�(�(�I�#<g5��ĕ��<�4S�/�n)��/B�u�ƗM�>�]�x��ٗ^�˚Q�+��A��붃��B��7һ;��y��K�rG�8\kme&�e����ǵ
��{���}/OԆ� %����+�����6�{ov0F]���w^�j�=��>M}:�|��R{��I��Ȩd�4��9� ��:�Y1 Y��e �������&��PCx�q=_n��+>n�������L�Rm�W�akB1�����9�#�¦�"/���.�7�\+�y0j|����'�	��cP  ]�z�9� ����ž���TgT��|�����e����C�s��Q��N�e�H��l;���-��V�`usR��}�M/�����S'�>��=�p(��=>=�K'�߉N�B�@,�r�\D�^C�T�};rL;'q�����K���C<lX���� ���[�uU�a˕�l�B��Q}�l�`؞��-/z"�B�_$��Z7�;�P6�S������-S�\e�`!l�goV���9�Y]36x��=բ�e���<�>O�ǀ�ں?�=�Q��H� |i� 0�+�����>S�$����"�����Q�N��30"��9Az4��1�C������k&�߯�F���v l�'B_Q�{0s��w\BT��W��4>q��_����9�O:p;����FcC�6P�/]������廓�3�p��� *�0<��)i?���u=q)�&��^��| �mzU�w!��b��#��Z���"0<�'�T;$X0���WmO���%3��r,旇�H�Cw�E�Nl��Ilr�a����#�m��EJ4z�e! ����0�Uh.��c4���%ݠ�O���j�K��9�t�4�b����c�����Ō��λ�RC�l�{�|��,L�y����k8�w˂fE�Bc��/�e5`�FrTz�h�u~ôR-U�Jedh��p�E���v�6Z�� /�E���5*�ؓ��J���`Ï�u9ߖWL_I��Y2�/��*,������l��f^�?~b�c��σ�P5����Z��K�n�#v�@�;P��~��D�����>q�,� a���`^�j�*�6x�G�t�ITC'M�0���PG���ߎ�:u1L&�q�[5=�� ¨��6=􊴫����lH�
$�,$�i���u
y&`?�zT�F�ͅxw�rK���\�o`��7_�7�W^�}���ʉ@*��#�d�Q�:ܾJ	Ɔeq�γ4����f�5�U4 2}������6������n�}?c=$��O��I��˼P<����E�R�XO�����M�:�szV$�����ol�Q�6��m瓓�yg�8e%���īK��he|�J��|n��b��N	gy%@�7��ٶ�,j��nO�/���9��Nɞ�|gY|\�L��|�5�CU�zմ��@B4_�A**0��>�E%�K� _ȑ|�l�{ tF��#lRVz�80S �E���P�`�}���� 	���IN�჈��c����&�Jm�"0��	9�5�'[:�{D�$�L�����D���5�ϐ�����/w�.l��	�$��������Α.0*�50뭎"�#�AH]PV]+ �C�����.��B�$��-��څ��@�}�y�a�]b)OAY(�����s"̧�u�}��!�a�}���8?��9r�,�<��"������[��ͪ���hǩy&ĦH8G:�1=02����u�e��M���wD��+{0,�iqP���5�Lai�-�-Nw��ۯ3=��$�oA�	�:��f�J�B��0������$���ʶ�A.������b����9����8��K�9?���T��(��d��0$�$��V���"��}ap4�Hv���O���H�!ԅ�b��d_%���ͨQ�ךu�zN��qh|��]J\~���0��dp��o&��'6<_�^�J$e"QO"�?�7��l���D�SFg�����@�5��}�I�+�P�:=���l�j�K{XG@�uPC�ۖZo�}��yT^����r���?X!�ţ���ys�CY�t���^��`>�v��M�C+Л��c��e�_xv�nZ���*#%���W}u��Z�L�f��'=�֠Ā�=eu��q!=��>��Ta�j-�uc�lA��]�k�g'����K��o9J������Q�صt��d׎e�ܻnPf6sǦ���G0i��d�Q���C32[�]�k��`�SY��vi�fEh���rW�$�y@nQ�C��\M��@����K�G���|�F�=��v o]G���ݢ\���ݗd��2��#:q9�1����gZi;�q�P+6�k���,��B�������Ez���t!���4���g��%�uo:�I�I�n�K�����ޮ����r�BR�#�~,���cg���:P�R��G�/� �$.�A���aB��:-��4��h��4���� P���:�����<+揰�YR�O2�o�L@���]��d�"]�I1���S�sIp�y\�v�"I��9t5�^��8�Epٕ��ㆌ���;�g�z�b�z�W
�%�zƹI+�A"��s�>�(��X���ڒZu
Ծo��h,n-�v��K�O)7]�2���q�����i�>r�����!!?;J�>���Zp�ަB3C�EѰ�h�h"&�b�Ȱ�X����~�?6���bS���w��������Ac M����V%�_Moa� ��}�p����7������@2'A�5��ēcV9�kw�ԏ��lP���+���vbB��4�jFQ$V�	E��8�v]�m�����dn�Š:nX�ItX���k:K|�%�^�K
��Ă�ĭ�}���Ծ��׳�g���?�f�^�6�'|�o@"��v�(�շ-:a�x	ތ]m[xͻ��"lc���T�0��R�~�o�-Ox�W�<���*M�iE�I�i<n�r]���_w�1_��lph8.������y�ģ�N�H@h$�뫼8��8��/<���p/�tG����������B��: k���/� �A#�[��*1*ws^�I���`]41�Y�Wu;�s�Gd!洽����V�y�>�~A�;��L�E~?}�R�7i�&@�B�y,�`��o���b7{����ط$��sC��NwE)o����=r;��̣���V^���G����@��z����M;C'"uC�W�B/����Q��|o��L�N��x�U.�-6��?��2�<&�,�9�OS�Y��y�������c(/ph7�%B6dY"�s���K*�(\{�cfX�a���[���\z�~S�4;~6�!�v�!'���{�B\\��C5jp�� q����z�2{}�Ͱ[��Z���^�#MO�q�gg��`�'� ]�<���9蠜�i�Hɧ���DV�����HD�8��c2K�L&Sz��M[�H�Ȕ�2�q嬊�]]-Ŕ�y�B�\�S'Y�,��c�}��f1Ӗ��֔\�'�����̅��["D�~4�����s3d+�cF��G�RIAl��pB����l��0y3�ү���|��z`���k����4Pd���x��_��Ǘm�v�-z��u�U��-N�{�8�"�C@��:@w���g�Ї@�7rN�ʸA@ݖ��M͓ov�:*C �;�E�7��^���� ���F�TGN��&M��2r2�p�6��ƯԊ�$<A3a|�LZ􏪜G�5 ��P�{�J�6i��T'Q3�V'UT�{��������s�ԥ���(�l�R�,��,�t��몡&-[1&\عX7��)����Ќ��C�8��ϵwUk��>R�#5D��R�8,U�H���ƴXZbOv� �95�G���Z3�X����X:��E>��s%�HȢ��ΐ췞��i�E�-6P��	�'�R�Ѓ�8&���)m�p�CCy?�"e� 1�/��Yh嗓-è?$�q����?�B)*�(w������"�&�#؏�\��#ǙesO\!��?�A��̌�'�}���˲�s�;5".2�5�y�ͩ�
�"�j����V�_�Bc�C�<��vJm7\^�I�7!Ƞ�N������U`WjL�xăhK����d
B�6�0l}�oQJ3�лjhHx��)����G>/�J���*�W@+�P�'c��TV����9�
ؐ�l���Fֳ�@ۦ�e�I��Io6\�&�ץ��8j�v���ccl:9���Q��l�s��4̨�9@��?�I�2�2$�a���j�G�ͅ���$�fVpˉ�#HϬEN�$I"��8�G�/�M���(K�:=~A	0KD(�bH���X]�m���o�Q.��>�T' I�t���H�/x��W96w�|W(�!6���J;X���KSA�����"�0�>��[�D��i����J���� ?1��L��2��PT	�c���1T��n��ÎB����;������?��E��Ø����6?��-m���O���nU'98�Vl�F���^��a���o9w�vqW�n�*%gJ#_.h/��rd�F�ȸV�ܡE�1΍�p��d{M�;�$]�v�Ψ�Iq}xX�lEO
��i[p%Ԋ���92sV�3�rx�FT��F�B���,W���L׽����h@��L���>!��az؉����@K�{ϸ&0�6���Ghn��U�	�J��)k��\J^F���i�F�����
�B�I�[Bly� c?�m8~�.���i�"Hh�Z�O(��mg�8��X�c���o�K��mM���6E<����0$��̆�R����~��㜓M�K�}_n��P�������8"�����N|�&�oȯ�؛yʔS��y�KN�� �<a�M�^�6���Ѥ&�^׋�>4��N���$Ҍ��(q�*m-r\�(W��<�!�U�4�(-���=Z����������@�>"k��`�]e�W���NW�ڱ��+�eXW:��� �[�Ї����ߕ]C*��7SZ��	����Yz���؃ύ��t���R�$���9���{mLeu&���qyrk�+��;���25����3�l����g�������:1ۖ��`/���M	��{�v{|�[N�] �Ü.iX	�%~�KZ�{ܼq�#�zwJ��&|-���ם���L?Ю^�6��C�=���̔�v��bI�V K���X���wEz��p z�Q$��A,tǠ�z9t����n|�?̅�_ �ۼ2M�#K4�9qۡ�v��oΥ�=�m��>�\����N}X	|ʹ���#�u�2Sx��L�V_����������ߟ�:Ӟ ���(�1[$_-�ك��� |���������ۂ�=�i��oR��f�R�ք�O�9�B��H�ɮjK�Q�xD'ؿ�#>��h9^�lw�'��v%��s�@wm@�E��SkH�F��_����A+Z&G�0x]E�NL���cLe��n��kF҉��f�J���@1�UO�?�Y�?�!�K,6Cjs�c@3��Ϋ<�����0�1_�m�G��~�mj~D�.m��f��r(�NᗪNA.D`��.�o�Q���Z���aP�wrq9�A�4i�������Q+����g��_�ҭ���(�D��!O�AwE{���XOC\+8�\�[�]?���ԑ\#��<�z�}�F�`s��s5e�s6�re���ah���K��*���Ʃe�Ug��2��k��.�E�D��
g�<�ZW�H8N�S�At�5���ʫa5z�p@����&P��UH#3.��G.*���=WUs����݇S_�2#4����U��(�@��jJ���K��h�d(\N����Y'?�t�2*����z��E������4��9χ�ͦ��zfq3�;0EB|�
���6Q���nӉb@��}p[4b1�u�1?ĩ&�eS�?>�ɏf�h#�*p�� oq�t�a�8���lC�r�g�Tɹ���8��B:�W�%����*��Aݓ5��^��Z�;�f�����
�q�����B(�yʩ��sqP �V$L@i��Tò�(I4T�&��S��Hgp3�;�E�	/]�/9AXFT��Q��&}r�S�,�����É���#g��`�u��;��_ӡ��������bt�8�9�.�}��W�5� ���_G������+	�-��b��D;�b8:^���W]��$����F�	�W�1]Pۡ�%��0\��>�->A}�ݪ9h�F�RyyBܿ�ac������_K��f�7��_Z�3��� υ's�Rʐ{Q���T!����O��v��`��Ч����R6.�	B� uKCS@p�\	(Naῷ���ɰ�c�w?�!`��/]*�꼕�]�3��w1�c�W�U����7O���.x��U3�ey�Qk?�,��P��Y NaZ����x�qb��-��XI^��{��A�+�F�d���Z��i�u?���%3�܃��x�=�?sbމl8��}j�˾�0��&����nw;���DJ��34MԻ�����߄!�0L��^JӄN��~l�u��,Zl%��H��/�����]��%!�hR���G��}�&|����n�E�U�GeOg��M��ƙb��D�h�fT��y���և�y`��k��@GF�U:��E~���ۉ?��2Ԉ��$����/M��g�<�B�ϔ��s�)��Q_(�
���y�.9��f��C�C���d��ϑj��u$&���믴z����WEq���$�j�����L,��Px�؜��7���b�.+��:bƉ`�}�a����]z[�����a�K���/�tJ�=����aU�`����t$�)R��\r-Y�B��UO���4nz�~m�ٴ�tol�ʧt
� c~D�Tw:��r@ǷA�>Ę�V���i@�M�*"4�w��I�t���c�~}kx�Ůg�	�L�g��WE��r�M�S_�A�8�\�&\��wg�y�f}Y��=�h����$����H� V��_����T�m����F��u[5�y��~��ª��"Kn��$v_Fs8�˙~ޮ�b'R`xP���t��R�����4���Cl�4<>x���	��&�t	��	R2x�(Q�њ�#D�Dv� �B��*C�?6zr@����j���&�]�o������]��O9V��q�o^V��hE��`��)�G����uQ�m��}\?:��R�|FD�)�?Z$ه�T'"�hxT�zdVb�0n<X�
!ĩxWEW\�٦�rH����`�<{�,�r���`��ߏ�V�g�� �mi��r��e|/��� m�
�Zy�l�a�n:z��n���]5^��p��iƁj�Α�	�r8r�����T��F�G��Ӥ����j�ϥ*v���.pu�G��:��TY%#T&��wM���[��R�N�O@w׷� @API���_�^'��k�9�JW.�d����T9k��WZ�W�
���	 ��� 3�0 ���i�5����ȫ��{�/1NCf,�
V� j��q�iz=��_�$:]�t�%QH/�h�+�ٰ��gI�){���r���I��)�l���"Z��A��T4��DRtTZ�*ܚ�w�q�|{�K��Ji_\tȈ�v���۽�cҌ�*^64�E�v�	 �:��sj6�tF��hP�Ƨ��no_Ɵ��|�}A�ݚ��3S��ny�˃j>G��͉O�
����Ͽ����"��~!�B���j��lf.s��kFD�"�0,�(]��|d=�<!�&��z�zqK�'�(����Q���������h�Lɳi�	��r�M��z���yaB�Vx�Ӌ���s!W>�:A����
F���b���;V'�.ϼ\q3'<'L�Œ�)g��)+>��_��qZ�
�'NV��k\��jڇ�B�J6z��n���Va����d9)05��v� �%��>����?�ckP����8�>��#/���S�S��˯1>Z�����y�]�v�AWjP�~��\�1�t�x�?��w��~���$�>�V�K5=�/t��=��=������L�K��2 �;z� �B�9�� �iE�Ivc�&o�K/z�(I�w�;�C��@��UZ�S�ioT��%|� y�2�����-W�1���m�q���d��Ab������?}){�QV���eɪK#���Q����&ކ͝J�-�f���=e�����t������'U�"��^���*��]+��A~���\fMn��k�j��t�����\��nS�@%�	��|��z|�W3�޷�ό���?n�J$^�G�a��Iv�������4�F����䕇���n��P��5"ZT/�8�;)"���������44[#��>�+�ԥmNs9Fv�)��b�sԂ���e��tx�M��m�<����]����_{��D�kb#I�"r���˃_�c���%x7P�x�}'�֓~��[D��C
d��./R��$�f���!��e�:�P߲�Vx�����d�Er�5�â?;c���k�q����$-%��'u\��<o����@�e���Ai ����i3� r˙W�'E��ПmF���)�^\����l��΀U�-,^��6j����g�Xnû�d�����\�ܥ��7N�A({ĚW@[Y�,�`���e|�T�Q���]f$� �*u3b�/���j�4�EH�;8�%��ӹs1�b�>�5'{�6�����V�&�������Y��Bͨ6���&�FW�z���W�b��5Ү0��&��1dE��Mv�S���p�U�X��W1����07�k'�����6�tN��c�3�Y��o_
�Nr���:��6\[�K�b�������lg�4�ХU=�N.1?���ڲf3�x�� Mר���1��O�{�P�e}� ò���^�i�f���.T����&��Y�I隫
gI�yo�����v-��X�%o�R�c�����7
�M�N�ZO���k}�ϐϣ�ݛZ���ڄN닶A��,�і��,�$F���/�������[�E�O����q%)p�\4x�]l�,r��!Gp�Yz�����z5�Y��|U��<��#��t�K���7�z. N>���~�_T�8	0�s�;_�	�x����ȥܽk���G�R̖���b�-�Iw�!ZP��]��?��s:\�?�,���6��xw�z�]�/-�2�1�$�Jj�J��	,yeϷ� 7��j*/$����=L۷Ra��"�Y�SR�Oƚ����B��	1_��q�tC��`��e"j[���Y�F�֊<����6���S%���'7�6�b���Y �u�,���fW\k'D(�rx�^�Fi@�kZĖr`�L41'�_=0�ȵ�b2�}�N�6*I�����eu�<�b�=�y�|F���%Cl���a)�Z��<�A8A��d��#+"�/]�E�X���JE_��0v���+$E�[�"�@t��I�w{���/��3Z`N��7/^g���L�+!O+O:���3�-ٜ��k�����Ȑ4�����D����8��?������}���Y�?���Zڠ�n��ҍ�����#���aM�o�^G�CHS^�#��z��S�hͲ�荃(�K�ԇb�UA5�֧[9��}��@��J�D*�Y�\��0��]��^@׎������>��.?/ E��tũ2��@zW���XRH�x]�7�A?�F�%g!W6[��@�e��������Ǘ�:<�}_J3��7�#�b�q �伥i�_~v�H�#	P�WQ��l-�� ЊLU�C�8���8|�{N� �� ��K8X���S���\YO��t�D0���4@P����C���ౢ������3�����]"�����B`k����p��'�H�)a����;㎝�:��- �N\�~պ�������eJ(��Y�AԔk
Z�l^XF���x�Vț�H૰�C��R#��-T�����Pf ����͆��#�|�н��m��8��i���ا	��������=F����k��C~��PR̉'cM<Z��H5�s���$^��4�j��߲f"�]�E��@�0\�(�sպJ�ʅ�v֩2�l'���ZR�&"�'rZY��o�N=j
����^ܱg����$(����oWޖ���60��bæ��=�}jC�Iچ��r�͸�j�L��F*�� 5�Ne��@�P�{�f]���KKLnw� ]&+��m{ھ���Tf��'׆+�W�J���OO��_e}��1J�R�Ñ[e��jp{0Wc�SS�A;���9��Nr�b�zN��:�$�?:Td�s��{��٨��+�M���a;,�r�2P���¹~d�$)[G�:f,���Y�����4z�EH��H�=C��Fɬd�@
�l��	Q���RMn1y�Ͳ})�dX��ʈ��y�yPY�OI{2��$��������9�#V5��r��!{�9�����y��R�2�L/��y��?�a6<4���е���P%�L
��D�zT���8�^��_�`����~���a.E��$G.k��<��&Bk��_)���YFw���+$�}	��i���{@'�J��t��Gq����Yc=vǰ����y�]'"=��)�Zϫ�����R4	������u�ETvXu��-��k�u_ٌ}E�8���)����6�36I���B�2��u;�w��6)ё3�HQx-4��jy!�������K�S2:=��?֜�ޫ�$���4^�N�9��(
���T�p��*��E�Λ? *S�ݭ�p+eq��%>��,�<��������S?������I��Χ�1�LA�*�\g#�1e�}��7/��Yr���6���r�\r���X�u�$��/<CE�H;�F�f3��*4���K�z���s24��<9�ߩ��#�����J�՜���O3ܳ��"��8>���ʒn�6�AN�����Dֳ7����4%�e$�?�Ĕ�@�@̚�P	�v�ϩ��AJv����F�3 Q9m'Aw�77��8�>[`ӌ��~{{~�˟�m��>=a�"I����q|)��)�A�Ñ�9Q�N?�YQDlat�z*Zb���Ľ��bh��?7�:t�)�&���)(�s���t��0bj0�dˆ�NiסҰ ���	���x�'�uO7"C(_�$:�6�9J��Qt�j�Ɔ�n�
��r,Q�M%��[��J�3�}��6����GY�ɇ��6.Q#�mԷn��4���xN��P�r��?A��MDkGddS"ˢ��=��54�Y���r�#!�~��z(v-1�GD�NE,�6�+s�U�m�%$o�'�,#ڡ�9a��ʽS��꼓 e=c��� w)�5�	���+Jل��b�� ����� R;�v��TO�[�h�l��?��RjFX>k�3���_� *.k�*'k�)}��x�9B{��	Գw�u�e�v��a�.u�ıP�o3 �/��j��'uM������+a�w'�`eq�0�By��7�2q ���g3�%��l6��ԣ�921�����S%�buT7|A�}�d\�z��I&�Σ���s7п�Z��zi�,���������Om��u�D��u�L_vR	�v�V�8E�+�-lN�V�,�-��T,x�G��#���D*�,��>�_.�g�J��.�/��j�{]"JȚN?G��X�
S��Z%{ǽ��Ѡzo҉�ԹʻE�N�`��VZ{�И3i��=C�d �-!z'���<�c�v��5 ����(iXO�w�O�������(�!\�5���T�-h�6�շ�"g�|H���w���c���M)Ul�W�2�=��Zn�af���U���	�6���tHS5��'��ZL�W1���~U^�t��fS�F{�;ag,�f�y�%T>�r�`Fh��Aj��!�)v=���� �L�������8�<��dXg�7e<f���7J�`�����7�����%&�q(PT���N����w?**H�?^Ԓa)���-�z ��FN��=�� ]�K=
]ZX�$�c�`y8N��,���f׋mG E���*1!��晴�y��pu���[6�J�~6���#�" �F�M��d�_z<?��u��a�l�0�(�X�+�r��j���^�*��]�lz`����?E1�ǁU��Vsit��'��h܍����F_��a�6^����W7&�\ 6Q�B�<G��qg��R�ibP�&k
���:�y2׳�g��_3,�,���쾲 2z��<�e��|sD6V)�[=��~��&�������)�ݻ u���̚W�@��������(��S���ް���C��~��c��{�2��9.���jhQGdFz��7]�S�۲B�l8�q�W'��,�.��:!1fj.2��cp�p�_f�T~��?U�XQu�O���� �vY���%R?���@��ıj�W�Ue)E�ڷR{�	7	F���@'W����Q�ϼ�F:�]x��p�.�	?�ߥPݔ����M��޵%p4&݋�X��ԞF��,]��]��'���̒����٧�1D�0��:�c�L7V�����.4�����<�. 5�G<Nhq$&��29���f�ObB�}9�׽��e|��w�+��n�2Qo���'��|�{L~�������y�@>��*���m�N�ƍ&�fw������OWX�����pY�3�l�h!�q�#Ҙ�j#g�Ҫ?ւvq�H\�4�WY4I/8С�q�w���O�=*��JW_���9g;��I�n�&NF4�=Q�����X����6#s���^���b�X�-��x.�I��X����{���܄m{�w1v��ɾ�N��7b��gț?��B֝~�n&��^)@6Ύ,�ĉT��J� oq�g����"�ƹ�U�������R'�Ih<f��!�{�M�>��=1�41ق�)vaB_y�%��_�gx*P�Gm2ڦ�lüR�j^��g�X��#���ϯ�{V�H�n<܎�S���V:��ف"+��s�+�M!��e#��!�h6/�bk�W�﫿e��Tڗ�M>���}�\�}���\�͚�c�oo�&y�r����ۭ��ɪvs?���w�5yk�$�����;9Lzc���t��}��T��TF.à�R�3Va*��L]�;Т@b��  ���r��T��ŉƛ=cP�'`F�|_�o
�D��~�-g���,dr��C��~m+_�74�����jƀ0�n�'3��z��J4�q���1� ��%�i�׮"c�����������&�����'�@�>�e�\+x�>d��Bd�j#\���밨�����B�Gӈ��p�zfk���߸L�h5��� ��d�G3E���F��Olԡ�\A�o�O���$GbWA0D ��c�M�� �.���K0��G�R�f��{��D�qXM��҆��i8�(�F����琜0/̟��ɽ��1�́G"oF�y0:R=(����{iJ�ӷ�ې��z�ĺۆ��QR:~)ԃW���#4F7ɜ���7�W!�hq��"��؏
.�r�"d��*]33�tp���!ewK�r��#G��j'�\]˦6�q#dKՠ�N6��}�R\O�2���Ϭ`lsv'�% �8�ߧu���;��Z�����ܨU:�AjR�zg�B-��y�:���0|[}&R�Δ����Cx��2i�A���|\j
,[b�ؗĺ4���I�,��
���M5�t,1^�5r�?��Yk� ��B����b�Xck���K�R���Ӏ��v3AH
��{�xـx4���.}>�D��&"��-,���T~�\�'�_���Lzx#]�20;N�E�����H��|��=�i�2����.�Wv�o����b����)5���\�^i໎d��Y �ԉ�S=���`tGұ.�'@�F=J7�cF[E�5��g�w�!��<����^����J�$Z� �]����������J��S:'�F�����7\Ǯ�B��M��*L�dm�v�-��ne��� ��^�οx��d6k��a|�;�"��LC�u��䳻��#Lfʞ{G ��ey%��PSz7$����%�4R�kNd�/� լ��u����5�����/�y�4�[LV�=��wc��0�����>aǦc���j���-�7�rF�_�+%�y�mu)L�>�2kHrk�9q���ج�"��ä��D�e��1�`cp0:�W՛��������2,�D����zp�����j��ɦ���I�]�Bf@�7c�U�/�̓%Hi�jޏج���n'���{n���ӜzIZ(�*OP||�}�>�xY�4����,��7R-��G��ж�]��� ��b�@j�m�u̟Y��1�z��=��|�������
!�A���.����9�=�D��@O\��W�z�6�Wa/�{J��Lzr�����*ל�7n�J�hF$�'�8�3�[�w�nW��-�q���N�K�1�
k��ь����'Ks^���~F�{h����p��JDA��4���v���{9�a��
��q�[���d��Y�eҫ"���϶Q�$��_.!�5^&W���F�-|*j�E�R;�+�M�Ź�P�l:F�R�a�*@⤞�/�Ok��q��W�H�����ı�֭Ӯ�CzKud�UȢ�>\U�k��	�����A�s3�:�;dv�jJ1��3:��z	*�`�g�ÙP��Cx��gzSc�,	\�71��
&��@��9����Y"��~C[��8�/����(�+sxx�L���U
B�߿)ְ����G�#�\�)1n��s:������A�={�|��e�zY�?ƕ��.�-fH��NY�z��S����;��&YG9�U�0�
U7Ap	Hs�i��H�jX�7i�Ծ��?C�`?��Dt��UV�=N ���6���N5"�)e躔u.��
H���+��N�6��B��4��8X�6&-:�>�Qb+E8 �s�g�%�!Sy0��A��~j{�IF�8�C(�Z���	��F:�ʏ��뮁sL��<&�������s� ġ�Ti׸8��G��BE�!J�IN�ІC;*b�5Z��;G�[dbB��$�B��ʹ�rG
%�5δv�f������_�^Ǉ�ӥp9�=�vx�j�39bEn�)&X�Q�{�AЭ��wZ�i�v�e�!��Ec�v�-}B: i-�BF����-���7G ��=m�|��1���)9#h�vD��o]i�۴ۂs�9f��iRͯ�Z���^԰�%���M�|dm�N��Q��^5�U��"W�Jf�4�y���
s?����%S��5 v J���0ؐli�e�
�Dr�R})�纽r��\pdFq)4m�X=��kZ ��\�Ol�{�p�C'�:T��J��������#ȋ�͗R����I	Mck��f�	#��Z㚂�E��l�]��~�L�Pd��3���oi�;g&+� �VY����d2+�-,�|; �9e�ɴ�8�t�̝�ʞ#�@�	��nv�*�gL��x��<u��3�
F0�(̯M�ʕʼT�Mg�|n��������3��?NM}�w"'���o(E���i�Idp���&'ޓ>\��P�&
�^�y���D`��6f��*�H��G�5���[0� u�ϕ���ٕN�z7ӮB��<Q%o&����A�H�|J�K;�)�"�i߇�7���'�Mr�Ü�@����x`�x��U�*�d�sk)��P��6Ft���2|�3K-��X��꽽�e��L��U�($q�5�����L��wTcF�PvЖ�]�'L8����aCi��<��c��1�ZFts�i��lu0 a�=��^�.#�����I��$�m�P��H�EM)�Ts�4a�C�7�P*i A��Z�T<k0|V���|�?. O5 hZ{��9������#Y%o�I1k���7o������*OW1��eq�R��E��~(A������l�Hi�Uδ���5��B�̀��<�.���0?��m���FAc�4���ϳ�w��L����Y�����nGp�ݸ<�K��G�T(�,�C�]�6'�tMu��:�}1m���D��<�"5?sD�M�W������G�G�)i��C���Sz��yQR>�� �秺 ��i�4�掠_��V��n���/{��J:��9�/��;1ۗ��F�[r$[Y`	D�l���G�N2���^B���{���ݷ͛~��(W�v�|��[�<>#�x��Ӹ#���G�ƿ��#���(�vE���~_kMFZ�?�H��Юz�	��M��V-�����1����q~f���T\�޵�J��i�n>�&��ym�X�,)�)^�^柶%jh]���N�>�7�*Z�h�O��l�B��t��-���O9r��	B7ǽ��QǕ�x���K�r6��;&���[)�7�I��p�8�W, �Ն�,\�-6����)� ����Y���k��z��ӑ�8��lc��N�^���k���)G�|M�_�|�!���L��t�n���2o�����z�Ĩg�p�q�L@��D���j�bTLJ��Ⱦ���5P}N���`�s�5��[H(�l�ٴ���V\�~s|�d�O���!�����Ƭ�B�LT+�f��z��=u:�����O�� )�CQlc�P�U�H�FG�2;J $�a<�1�x���}r�0<���ze�5ȯ�.�ݾu���ϸ�ι8�F�z�7�;�S>?E�mJm�7mN�XR�`+��vEm���L�������r�1���/��w`�A�7.5�|�����)~�تa�����I�=�����m�`4��'P<uf��jX:��<
wU5�
X@�E�?��MÃ�4�/J8[@���;~�R��sD��VF�TOW��G��IU}!3�f�y
�-�Y˂Y��ϱ2�,0��e�&�4�qfN��Q������呂�s�4�+\�f V�����U�!��F���I�#3{H�U� n���	���)��|��25��wk��Ox�Y_��.8]�z0�����B!t��yÏY!���4��}
�8-)P�{;��j �ۮ�����6{�I�����������ڼ;�ũA�Akr.&�� ����F�Ѵ�L�;Km��Iڢ�d�QfE��1�ٲ��^�v���f��fh��2�& QHҩ+=ͽhAt70���c�vrV>6M���{r�W-Z�4Ng>tOWlE~Pa~�f�y�x�.��_h��%�'�)�bʜ����k�BY�]�G�T�XEu� �չO��]nY�|5�y;o��*Ԅ 8�9��ֽ�����˕��ϟ�yLIܧ���ڦ���K��y^�}ٮF���	�_�s��w�@�v�؍�ŋ|3�\�n^��>=�-<l(�h܎[W�B�ڜ1o����?�Y;4�U:4v
ŒY�#�3�ҕtmp�1��������j������Y��-T�G
���#���k$(QE������M��d�+���������~�#ML�
�5��"�ep�X�r��m���2��xR�\:��#�\� �8�o��^��"6�h��$��{�j�|Ys^��'��b�ھ�M}����V���Hqy�Q��~a�Gt�[<�;�����Py�X���%�+/x��#Y���_v�G��t6%�X�D�Z������,�{�����1K��,��$�����q`C�Av�S]�h�َUP!JVn��,h3hi��m�i{K��vPE���w����&WWÈhF�����Tc�uV)�rN�5�fX�Ȁ���7�+o��91� 0�=ǧx�^N�~��l�����.�%��]�Y���}?@��V�Õng�Ԋ6�$���z�k����R�5����wj_,���C4��gƞ�Y\�U6y��Ik�u>��n�S����Zwh�u��@��������+�����H$����c΋	`�|����lՉ�ud��=qe����V �Ѥt��t�7����E�)E�=��'�	�}�&�|����Ri���R�RD�!�����4���<p�	��MT���7l&�ta5_�UEg�*�h.�J��)�׃�]�m�)=��т�^DQ�%rUݫW+҂�P+J	�D]��NA�E ���C�F���4p��ڮr�xf�P��x('MxWQ�ӹ�����d���U�m�(��'�:D�y�^L!`�p�"�b|�x
��}IMXa �IJ1���<�[��g���
kc�F�ktr�{k����F�?�I^$Db��7��C��]�=M)��Z׳M��o/���C���v`��J �5����#F�3X7
9�pG.���B�02w���+�ք'��Ѝ	�,�ڧ�=}˕�H��=ig��N����;�c�������m����b/�[=u\�0�M��.E���am���2I��ы�~��@6�l���3��O�a8�`䦱%��Fs�<�#�[�C�; Զ��o>�.�h�a�kAʿ����D�E_�`Z��E�TJ�s��8�����[��o�ľ98l��W-���ec�Igr�<5���x�cA˝�¸n� ��3�p(�iֱ}7�󩈓�WG8SP6�ks�����K՚-�9ԟ��3+; ��g���P�����gú!f��|�t
R���_Z�8zi��H�J���"O����h&�Q��ړu�m8[/+S�% 3}.�rx�\n�F��:LO`�ЦG|v*)���8��#^�h�y�0~�s�Ű�n������:�#W�dۣd]�����T�s�����U����n��F��(#\M�JK����C�Z�2ԉcΥ�Q�q��9�	lJ�͢Uo�	�.��}����Y��.��W�|����+��Q)��Q��G��8�ֽ��m(�P���W-0��v��};0�T�d.���r���X<�L����}��P'R+8<P��kO7D�Ye�D�8�"4~MC�[~�tL���e�~_mU�� ��A�8��\a�p��W���73g��߶E��J�5�;�U4�\��9Z�G��8/,U	�ihx�_���9^�֪���!mx!ׅpiҖ������.ª�S�/�,HZ'i����y.�%����o�O�VQ|W��N���"�N��P
��߈$.uN�Ӆ�����j֙?{�����v&"ؖ%���M��g%���*h�,p.�>�Ǳ�!�䝳C6K��BKi�6\�n[R�z����)on����EE�i�=��2��;��2Ϭ4m�2!�-;8��Kk�-��Ë���O�J�@�#(U���@·Y�Y��ٺ��(�\��Z�H,�i�����K���ē��V��,�����t��C4��7��0�H��x����y�!���w����h�r�G��`�}�Ǭ5� zRiJ0��~d�^|�Hw������&����@��Qgd�i�Yy�Q��٠$�)��9wL���.�z���",r�݈ly.ͬ�F��"lT�@�?����>(-��{Vk�����I!�5":(ދ�o���>�]hr��Ul������9pT��O��ss����z�b�i��O��<�D�I[A<��?;�� �����h��2��m븳�Z�j��?!�,�ڬ� �5�:"0�Y-3:5Km*���MU��}�bN�9���3�:�|��JQ�n�"����&%B�f�|{"nla��7,g@� ��`񰷴h�?�G������aEף�n0�� '�:�F�������ЎJl�.>�=�`�I�Yo�Ub-��%^{mp�ɴx��ǀ�V��,)�&&Bf.	�(
"�}�d�f	���u��b)����@� ��z�78���}�[/J�� I�^!��s��
�hg�����Q&'�kw(Q��~U;��[IՁ�5P�'��JjdY�T�tM��สQ;�y(nU��>���#H�u�4p�����F�^��(H~��Ӗ3ɋdOO�����}Xģ�N�5_���
�1���H߂�涂�N��DM���4�pd ��r��z��63SG�!#�?��72H^V�������Z/Y�)G���5�08���K��wp꥕�$~�<Zm�>����ǐ�K����MJ�u�����-�e��k}*8�d<g!ӈh�!j��(4�kl���-E�6����Q�B��Ѹ�B�������jb�i6V�JV����@o�s���[��6���*4����#�QƦ%R�?�c���J�:���iL���cJnbsp$�٨@쿀���{�8 X���z�,P�E��5�1-P�����V��#��t��k(�#���{]{�`]E!�y� �dH&�^>l���W>�w+�O��}�C�P�y��r��~�p��w���;0v�����s6��sU���7pL41��������Hz�ِJ���*0<;KH��=�ֵ�m����xT�mU@����tQ�w���GVw�uH��P^`c�p���QǼ���{ԅ�W�"?�x����S�s�E�jۂ��h����hko�| ���=i*����ǆ���lo� ˂ί�z� �\�݌��:�/|?�K����_Hp��U�����A�o��Y�%�� �GNY���}뇻�!]�x���Ƿ�(9���?���|�)׀NX>$$c�i�u��'��r�0���>'xP) �J�a�l�"�y�"��4���㌞*��T�1��7Zg��8��!4E�7��,��a� o# H����0݈����qP�0��dh����|�N@��x,��&J�Ua������hmZXs(ދi�C��>^��}�&>�s��<�>����VlUC8�,�Ҳ��'[�a���>�C��E��<�`��t�D�Ar�)71;����uR����V��O��v��;�7��������@n&�������N/�A^6x@*U�e�l�I�ZCr[Np�)��~^K�zQk�(á������Kl��?Q�е������+�G��爀��Ke�nV���LC֤Clʩ�܊_ÏD�����ￗ�5�U���y�W���#7ټK�}�]���ҭOO�v�kÙ��^7�a7/oJw�1'��0���O4B{:Žm-jw�/_�IKmc}D;��BW�V	|�n��v��W8��y��7�)Z�"�"��:�<�t���=����V��84��cRE�{ ���B��%Ah0�]����@ڛ����ewYT�O~>�a�i�Yx��O� ?�U��z�K2EJb�Q�P%���մ�vK���1}_��̵�j$�3~�V�����W��q����L�\�d)���0��q� �G���a~vT�m��.�8�n[�H�h�A��"r�~�d� !7)
!��kf�%���LI���L������グVw�v�����w�Zmt�gk\h _F�X�:!(��7,M 0#��;'4o�p魱�v�QE�!z)IHΛ�e��99X�Џ��%L�/fL��� n�R��
�Q�XdJfnM'DXg������F���-��f�=!́��##02���Ô7� ��O��<w������rPOp�#.%�Ǝة$�������ވlJ��M=Y����XE��מ�xo�	����z&��9��簎��7%d�L޿>�U��g��vR�>'�?�g.�w�:��-;���f5/j�3��+�ҶYR���������i)*�'V�aO�s��ņ�^�&ov�j]ՓF��Zp@�TJ�/CF/k�/%1H��WCr���kx3��C
a�����@ys�\hzÈ9�N�T �����-M�������\��O%�8^ǻ��:�m�ں3����'�?jo��L8>=[L�����������ܭ|%�C�Cwv;����X��������b��P!�Z���7�QR�LJ�}��`wh�����X2�6z���:W��y�UX6�ʟ�NA�xe����т�\v�<���Y��!�]�m��R�Ǚ%��dG �,�M2S0R8�q$�p�`�r+�A�P���0v׾կC��pSNj�o�ݿm���,��h,�)�k{��MRC2�qz8j���{�?@��t$������l �]�M,3�M��~`����K
�VM�7������1Zz�m8ќ�8(�d<}0x���%3�(��j��Kbpr(��8�@��=_��0͉��z>('i �W�<�G��� �|^�����^����Ӗ$�|��TBę��D��{E2]���:	����O?p�M�N)ވd�Rh���"<���O�=�q��}���\����@�x�ЗC]}A)J60;��DL>��!vK5~���%�q����9j
D�[���!~y���8$3n�G3vS�;�}|�a��AG���@6��+Ӆ-<��`n~�l�|8	��J��c}S9{�cN?l��t,�˯n����ou���C��P}��(�����=��L+\��D�Cs<�#�O1̹lL�]��XDb���	�-B�2P:%��Ѵ�!i'�uW��+���}�KQ���z����`T%�-���1ͣ���ӿJ� ��Z��$�yx,<�O��"R��/��e�$��2���jU�:x�+֗.��,���z��\{9*�jۥ*j�9�mS�+�pP�e��[���Rٿ�-���m�����'pL>�tʙ$��S���-��N�H,�gAu{��":�i�����~	���4��c�)4ccD݌�=knC�����jm�^zi��1�XD,R�6ҁ��0���!�8� ��F#�ۚ����p���bo�<�vޚZh�ǁE��t�L�Hc�~��m<˽�{aIS����5P�Ǚ�9Y�5�A����Q��T�����g�Vҏ,c��C�چ^���<��
WR_8��[#�����LAF�K��W?�q�d�횚Ή�}�e�����ʆ�V�LԀ|�2��m��0>�ם�5ox8��|S�o��'��g��r��đ1�*F�U�6M��=��� ���N2mQ�;��#[Ҕ���ƕ�@]�:����r�+&Ɍ�0��a!�h��h
�y|�y���7$[ᥨi2�ޑ�K�+B㗀굢7o{�.���B��l����&bp�f�UαT�� � ��A�ZA�]m��_0��j��kK�L�
��~5��M"�ʟ'���@(���<q�t]��h�:� ��N�k�D�l�daт�=tZ�%�fU�ݹ���&X0�+n�K�<b̹o[[	:)�]|�9�q�q��od��z��_�Q��ە�����,�:U���,����c#u��/��,�X~�W��M	�Pf��
�K*�ZAb���U�5}�ƵM�^���x��#�����&��~����[�[�vD����a�L���W�)�]� {�uт�� �R��E�q�bN�@ݩ��rg�r<�1�w�n4��P�.ֆE�\}F�|�>1��BM��1瘕�p��#�";x�-lZF$�T����v�H��*I���9����ϒ��U{�y���!D4߾Uo	�2�w4�>G;Ϝ�Ԍ� M�=ۇ��ҦGVA��,�����%0
ZPV���Q����~��V��6���1V���)�0e�-XN���*���x�Hs��P�ȳ�\����Vy��T!�Q'��]/��r좸��O&�}�|F�{qㄴ�P���ե�BMר,b��5�)N�3Ќ6>wg*�c�D�i������s�Z�Ln/�y�������AJ���|�lG�`���~JOI�Y��߈W�u�S�X��������=EQ<�).$�ZCV��Gq����3?�vx1���!����/�ޯ�􃎏*��s��.��F��_��*c��l��r�{�E�V��"�7�GR*?]��'�u�1��͂?V�����5@v�}���>���;�X$'-۹����<�1�(�7���wc���#��b�+�<�gC�z�?y��8��l���7�_`��saǋ������	�ߟ�^W<�4&R�^�
���ܺ��E{�����s~�--���t�ʖѡ?�� �/����	���{1�n3�b�4�h}5�����*�
����d�WX� �R$1�I�w���A2q���m��FQ7�{ �G���$n�c��HJ�e0��A����ky3���)���`�|�1< ��Cp��u\w+�]���-M�A��_�)5N.)��%��T�@A��[����������t��ߔ����-��۵�(�)͟��nI�����w��d�Vq�
��n�6qu¯�W�:upѕ���R ~�c�QH��'4yc
�{���v��g�TK��Q�/��d����t
��*]�����Յc��Q�5
��K�W�X��w��r�m�WH���ſ���:�Ñ�j��Kl����JS�pK�p�,���=Y�ۇE���zE˽���%"�#8��j�$Ɏ5�&�����k�<Ն��i[��G�����!�0s^�u?j��C�2����ZMG%#��Ѝ�P���s6����� �?0*���^�g![�@������~'_r)KV[����×w�ۜ�P�ul'MC?�u�N�;Jꥑ񊹓Qj�X�����$c��Ŏ�a��d���:���g����NŬ9��7�=!|�%��^h�4�m]�p�����	O��h���o���-r�9�іzda:��`��S�����$�Ϡ�����J�>幭7� 9TA
$rT	���}~�KXn&���e�.�<?�z��Q#�g�9����p���mͥ�
C����A9�2���Ǉ���ϻ�,i�ѡ ���>v��64�-z;�?��ۭ+�X�WL
��h�˅��u�=��[��Qԅp�eW�����-��U��{�-�����:� xa�S�+|0E�v`6��((c-�=�Qd.���9�#ON��7�>�^ q�"J	C�I4t��9����E�-�&3hVI�	��A��enKo��y};����/l 42�'�vse�%m:��W�/�G1J&�y�c� �^6O���cؓ�(7�-�,�WG�k�%C�[{aD�wFk+o�L2?��4��/?C��%7��z!�P#���ٱ�0�V?�������2݊c�V���RtN��W��2ɏ��{37/�Ĩ���A9���jLděS�M$宗o�_ȵɉ���8��y���*Xw������Oz��|��V�M�(W���6�eTE7��EWʤ��6������]�h �ƿ1��JǖJ��&��U�Ӌ:��qG�g[Y;�3��5U��/�Si]����O�U�L�n��ʪ�]/��por����*+��M{�=>���^@@�q��Rr�S�ޝ6��*ѹ#�1�]yh�9U#��r�kT3,ES�k3��%y�>
Ћ���l&ͼ3��x�31��s�3n� \c��~h�3�q��v?�W,�<A�7{�8��HN�6҆
PP�CV�*K!
dB-�#@E�N%:m������B�/2�	�R	C���K��z1��$��O�s�w˄c)[d��Ԇ��ۘ�[��Q�;��L��ETD���-_�u��N��&�C!�)ˡ�1�g�����C�P	Co�X�ҩt$
�2�b��ER�ޤg���sx�.��6�8`����$�ր�������������S�³�ґD��W5d7��)�_�F�������eզGx�*�� 0_�3�I
J��!�0���R��m�|�b�9/9T��6Z�������z�>��g:Qw�I���ZH��5�ݻ9�Z2�Ss�i�)�9B\��Á�	`�t1����>l�g�Ε�BGLP�@�\WV2XP�e �I�q�P�)�϶�T��̈k�L�L��Pp;/��
��XTEyϮ`�$g�^h�Gy\���J�N��=�]������f�#��tU����wf�L.@�r%WM�oX���E���W	P��ˣ�c���(M��D:�<2�D��z�#U\!��Y�� t��05ؑ�e�h��Ei:E�R��F��ŕ?U�碓PBߚ�xEDf�I /%;�f�����Q䐝Te��Tf�M
�mp�!��(�[�������.v�g��T񮰃ޮt�u
�eEb�ŵ�.q��pk���k��I`s෇Ud߿q�%���x�FK��t�����8af��#w��"C_�V=nd�kH�@��֗#���]'���I�vˬ� *F���,�����P�փ�N�;L7#c�c�w$eIF�#K��h@�K�s���r��.޷+�X
j)��oG�V3}�op ��}rf�jx���v�jO8��n:m��0q�7�&������_�bMrLEb[�	RH.�4�ܐS�̔�7V�F�����ܕ7}'Ǩ�#=�8���j���~.csi&��V#�_	�4H�v ozvܻV�!hd���p�-9�4���;R��Đ]��%'�g~��6fp��WY�oJ�q�Q�uM~YJѿTN��𤡒����pz�9	L o��I����+QN��aމ�b=��f}��ԏ�iގ��xli�)�R�=��Otv��&�<�:0�F��:�t�[ND���4����*��N
9(V+��XӶ���֪hJ��b,ﱴ��^~n	K>y�����~���V������A�o�*q�_!���]�Y�[~�.�uG/��
�;�k7� �׉��R4u;��}�i˩��Si�}
t\���8uy�/ȣ���ЖO��#����;�ʼ+����� w�êt���g���1��%x^w�E�n��G�t�XQ��M�k����mPD�ˬ��Z�%��W��|S�q�wv �����E^c�Be{,���D�1c��z���d���bxa�5��Mij=U<`��_U	�#��5
HE�w@#�Gٮ� ��a��2O���jq8���4�f��C�j�-7ɪA��+�ީ�8�j����'�.�	�$�=�!1I�e���[�%(_�?a�o��ω���!$ɭ��&�����1`�bNw��~e��5��K|&���W��G��SBV{3F����d`/�O�B���n����!2�|�[l�Mk���>�k`���_�N��L�~EU��dK���v���X���ㆰ�r��o�頓�$z0���&2
!��-Ō��U@\+��|Z�Fo����I��[�Ab�x�0c�s��"�{�Ec�#83�,���[���b�=K.����.T��?�e
�n��bhݤ⟞�m���m�`p�X����B8�qx�\$���*��|SzG,�<�.������﷾%G��vY�M��O�{}S���g�LE���$NS�Y�|�ÇG�]��g�����  ����/O�e�הH�xh�|./im�"�h���������Y��G#�&m�%Op������E=�eS�|� ��v~l#Pk@�	���f��Pȱ����ǝQ^�zc��ox[�������=��g�o���� CŚ|��D8�Q��eD�ڐ��g(6|'����Ğ�&�7'iQ�h���DQ��$���M�F�	щd�>�^�@�������9��>���*�W��6����o���������βx<���-|���\^�#�q~�ɭ�t���wrG�(�ªQտ� �3T��ͩ�U_^��i{�W�� ��E��W������*|�l������K�a8j���5,�;��h1���1	�K`fɔ=?�~�"96b���PAԘ�Q�WϜ֯���0A�ˁfG�F���CO�_�؀r0�M���]�UEo#�찉��J���w� �kvQq�šO�,��A�}�ZE%��u�ʬ����b-[v���S�*��71���0���F¢��U��o�� ����3�:���#��rpJ�1�L�W�Xh��`��"�b��.��60q4��Lq���?ah�B�r>jR����X�p1nU�X �b���$�ļ�0ho�4X����ɰ���T(�(<�6�_��@��0Sn�ޒ�K�$~��\���4��MJ�uZS�l;l�����b.��F�!�AP΄@�ѭ�^��/�Yq�nZI�aF�a�[�L�	�F1��)��]w�B�7.�Up�P�L��I8H�o�M;
�\�z�$��b����U}���� Z�\���RS��֪u�e����uV:�t$��9P����d0_�<=��5y
���F��B��ؽ�'@�zwt�|B�i{|EBu����j|�d.�1$���o���4���3��d��`�C�0��\7Ct��Kq	Pt��â�7 ?/�D�������q�Q����d�Y��۬"���V�l�����i+�\�kЊu�NM� HY��J��^HI�`��	��#�Ǆ����<��E�H�;�\BD9 [��!T�}�EhO�j���Ey�����U���_xhؗ��h�+�X*�C��w��-,���nS���^���	v�P��H�ץ?��ۆ�Ѽ
ع�����=���������~���߿�)�xY�~���-T��j������bŪ�(צ�ğM� ��T�����˙e _/�.��U�G1C�
���s�����Hgw�'��v*���(�ۄ�B�#4�5�i�ƉC�_�؟��n�Y�`����r@�S���)��>�$��fN��Y=�*u\�_��_��Q�j ��y9��� ��j�A��5X��{�)��S0w��o�e�@�t�j�a���L�a �d����$�Y����	�T���P�q��"�^�V%��
��jr��t �kJ^��n_W�ƨ]���`�n"�R��� ��X1�s�N�]i�<�.���Syu���9��k�<�����.v�%�6�����yU@o
���k&H��@�:\���u��c��o��)����˱�E�z�W����)�TX54�vSo�~:�������i ��HJ.]{��"	܇�l��6`t����\�)����󈳎��u;[տ�2�8o|�*��%qN��{����I�x3٩�{���E;I3�6�8��@"N=�H�g�LxJ����ZWR�Ы�U#�hސ@0���	�+m�[����
��������9p.)H�#LѐY���%*\T�������B�e��ow&������	V�WM��m��.��1��;�Q�W��w|X�d�a��-)�o�nhʤ��a�ʰ�����)n�s ���!��{��K |�ը"��N��[Њ>����K�`�G����Q�_5���*�r��ӥ�D�|�H����`o�I���rԷ���S萡����%Ȑj|Vf���ilLt�-'�nv�J�R:�fѹ������mδ�%����ŷʌ�;e�iQ7����P��J�m7`�Ŗ��y=�g�)�6���)� e&&��tXe��f���^͍��@�u� �T�m+�t2aB��i����4���H�7[�ǖG���m��P�	�����iwGPkV>�ЊX��!���U��L��R�r	N�E�UI2�]��ܳz���ܯ�=�1�7��mq�gٺ�51ㆾIaQ������}��d������ �k�&��Jc�:/�1�|=�q��F�O�۳��p�f���0>`"����Ӱqw�sK��L��}|�m�
����)SV"�cl��P5J!m41:ٚ���)r�X"4i�D��G�c[C[��y2G�ۦ��U����;#��iMh��ɶCV�T��>�;Z ��T�}�;�?�E/��-��6����v���!]�+˄ͳ��E/ī,Y,e�� �Y���_�1��HV'.��ON�m(Ao- �W���sV8F�t�[��`>=��j햤l����HL�[��D���:��6�(��Rھ�U.;)~�l�����I�"��{{+g~�5�Y�9\���@�&�GJ�v#�=3��*��/q��=�U�P�����`t"���7H?�$O>P����W@�3&A�e)#��ǌm�'�����GT�h����iO�W�Pw�ʵ1��ߢ��y+5�7ϴa��Mi[�zYaъ0 �՝�����Uː
EU�M��E1���d.Â4x!1󜪐���S��C����c�l�Kd'�Bޅ�Uk>���:��7G��S:��u0��mcx�)73d���:���e�J8�B�b�:a���*1��$J�5B�<1Ϭ��/�_N:)�W�_1ЎFҲ���&c���ê�>5��?a�$o�j���DI�����Y�u�N��D���@u<ﳉvֆD	r-85RQNw��u�4�h.:f�Zz��-غ�#��d��5Ӟ;�(Xɬ
��F$�լ�0��� ���z??'Sྔ��<�)3��0�s���Z��k}�6�m>(��*��ƴh�R�@$\\���شK���u�J�-&�@-��i�����˚��R8z�i�ZA ]W�'�>tD/���#�+��������Ȩ6��1J�����H?�E��h0h�亜Ҙ��Ƒ+�G��{^��͆d���c<�162��vw��ʮ���W���6����*�lx�������X^��p��ҭ��^���?���t&�Yu°$hh
OaOIP�+mh��J������EW6��ߺ�����u�n-�b���%Њ/��`�l�����E��GA� ,���m"	�?��q:���+���#�w��٭3\����A�8���
5F���2�^&�l���ͽ3v�Y�Ē���٥��bL�4��}��&l��g�p�����m[b�������pS�4.,�pɖ�s��d;$|�A�E�$d�h�A����Г]@��U�ӭ��i�	���Xkn �'ĽV	�Г��i�pB��d����[�j�QYq�DľLߛ�/a�8��^�Ӳ�5���#T�u+H�9��p���k�������
A�cG��(�*�Ƭ��K�ü�I�Xk%��c���I�	����O��߬�G4�\����?3��W*"���/w�|���*]O�}��n3�'�Gcq,�-[�R��wq�OtZ��RgPcl���� ���k{�+31�h7�,<=��bj�U�|��p�@c���Al%��oPi
3صd���I~s[F�a+�������MIF|���u>�X����6/�dƈX�`�����\CV�T���\�ծ�7��A�C�&��g�gl�°fPQ$ӣ�F��=)���$}���7���Ҙ����2��g��?7Mm��~�[����e����<�����a�����,%����%>6[f��=�$�R��Q��1ĻcU�j��!A�:�X�-$�簔�?]��ES�����Ђ��D�~HCJ4.���Z�t��`��U~_4&�s��YDc���MV7���P��: �4����e��������L?v�?�������G���0Y�W)�O��|h�� W��@F˃���M��%�P�x,���[���f+ V����� Y@��n ���4��-�N�͹rUb�>���N����14�t����ZCc���x`�+*�"M���w�¦�;WQ�i�#i�5�6��Hӈ�XM~��&�f>S�C�Z�T@�ƚ�z`�yDbaU;�]0qQ�]C�=k�� 3��-z#�%#JZZt?���ئ���.sB��9?���4�=w09�o��y?O��Ϋ��Q���)����8�(6�p-�'J����:>�*�;/l�������^�XGlA��e�4v�Uұt�>jv�W���&�,���P�����-���Y2d[��-���V��&�leΑ	Z�V�B�}n�A_�Tz��t�X���M��ݢҬ2ͭ�\m`ɍC	zs�O�����	�r��L��p?�!زV�w�(�I�����՘����8�ZݱI/�X���y䟔:����ʾ$'<
��9��^L<�O�A��C��ی��*J���T5P��%Wz�Q�T��_jtv�>	x%�����	y�9��|!�ia)J���3|�#�o���sN���aQ0\���&��QZ��� 09,)��o{�S�q��?v4������_녀�B�ה'\��$YWQ����@9��k;�� �����gE��n�K\W'+�7S��<����z���Cu�U/����ׄ��J�.� ����~��nhe�~G��G�8�I	M)�t-Dvt*[F)|�����HF��Go`�Ѥ
]�q�2r S��v�L��|�j�αLz��Y���m���g��Y�S4y�S;�G(���*.�b��R{��;��6�ƀŜ|є� ��N��2�o�h��Ե�J���Iܜ:RP&M�X���=?��5��0�܌�����0d�nm��<��J7^2�!>ѐ|�0)Ǽ]������s���yq��[�����B�QD�^���{��:�Ic]^��pb{�	��D�&�K؇v*�L1-F��Ҽo���q#�S.t ��@oy��
ۖ��!��6�~�\�ݣ�p��ٛĈ�o�`����LZ^��)WD��:X�v�|a5�SY(�B'�����������p�;h�l `�ZI��T��<��6��ˆ_��L#MV�4�D`B^a�`��;����W�S�t+-��[}�v �z]a��$T�05���΋Md0"6���9?�Av��mjS�8�(��� �F�D��~�m����y��6o��+w����o������s �cZ�R�HFذ��J֪�߈���q���A�e�p�K4������U%�!�Ou�nC@��JS�N�Dzf���&��M7���/4mo/��]:_�=�����q�i����^��Stb
�d���9��!�Z��:	5E��L��ZDj��u�uD�����Lk9T�*�Z�4�{ْ�/�j�Ցf�{�W��n}šX`�
kU�
-���mubH�0�P��@�hǹ�_����!-���\�u��?W t����I�P$+��K?��Z��C��H8�Hʆ&~p�&?� <#zH�� ߙ�'��h��# �۸P:ْ- K�?�.e���!���9h+f>y�n��d��5�V�&{�ۮ�ϑ���n��
�򓒯 �j
0���Dk�*m���d�"Q�]��BZ��m��8!�C!5gO�_s�{��؋n(������5�f��-���y��$ '��k6h&�0C�n��Ԁ���s�c�@%OU�0`�?k(��?�����J ��9���9��|ȱ�}�2,Z�jl���.�Hd�`�p�_�Z6h���C�h�=���Qa��Mc���-�4�RP覫����w��Z%'�ά�?0n�5�̋sI||� D� �|6��=�~W*ŝ\�� ��"Q92e<��Eir�Z|�u���� �v5�O�~�����%	M/!=%u���;g<8�l�4v�覶���C���!C�4� �[���JJ��l�!�����H�fFd?���,��b�-�l-�v m��6���ȁ�J��o\%@�������z'��?;/HF��z�@ߐ#�y��ztI�1��5z�����{v�c0���c�)`Ś����$@�����.#I�(H|VM�k݊�UV�ޖ��K�U룪_M���@�i�0>A<�ϔօ���B�Y-�>��;G(/
y�?���D�iRq<W2
���
ʦ(Z��u;V�0a� ��w�Z?�j"_����y��Ș�_���8������$�<�*&<�1�N7.�ar���)�jtq����8�e+����
�g9%�dN�:����Ĭͣů�b���B�1� �W-Re�좲Ē���Kۂ��t�V�u[RUK"m^]&a��_=�;lh[���m��(���!L��ړ�<x��/�
�q�R4�+
W#�kO��lS�j‥�w6�
|h5x�n5�Ss�H���&��Y�11͐�=O�4M�ۯ�k�����������U*��9#�u��lFm(�����a� ᠕�`�{Z*��8��9��|��Z|S�e��۲��VLu�Z�ܵ?i��ay�rK��o2u~�j�5S=�F����3�D�B�
��n(�5`3+����u�ڔ5rY���^ϠK��eQ:N~!�����jV@q)��#��}J��>�{���o�W����ru)�O�G%�7�R�&r�P��;����/d~
�[q�`�q|�����v����Z�h��ɎX�u�F]���t�=�a	j�o46�ȉ�)��k�N���qqa3$?#�8�~���1墡$��0
��@��i��|�D%�Su����`���b�6 ��I;�c����T77N���)(�R(��!�5�sџp']��oޢ��W��"h��e��R��Tc��t���gW0�]{�ϔ�N�y����8�CD�l\��B�ӵ=s-�2�T;o.	�l���B�!8�h_��Cڿ��5R�Ȗ�9[�s爀Im�^>8~��Z�p��$��\H}��q�b���w��5D�r��S��S���^ f�r��/�� �X�d��6i��T.��^Ч�R�zz�Ed�J� .�d�e�s�;3n��x��{�ݏL��Ұ,ǿb�N�c 9b}T�B)��%�V�pl�S�C��h�h'ݓ�R��#푹��v��E����H�X���j<v�KA�v�p��D2q���;?�1���F�'�H��7͡=[=AdU;,F�:cWb��RUD��~_�}"l�}�9�'�=��cH.�fvv;kh���.a����<!��A�ǿvh���Ꮼ�\ke{aZr���J=�u7��ƪ��L�)
�Z�| ����H֤�����V1��̥8v�n� �0�9!���p��>�5��e������5fEG�7��wQ��=�zQ��d{Jz�,ڬ��!�\�a�GF�|4LJ���E����s����J�r�}��B��X�.^x�=mGF8��F�40��<7����+�"�p�UHT�8�J�2)���b��吿L��Q��J1���<7��ĝkq{p�5DHb��0�a��@(�f (!�1��9�{Nu���|s�;��B�$h{�a�N��敱��GgjD+R�m�����9�ߵ��~4R�L��O<btd��w��XjRb���	)��gӛ����:�pm��=�;ig j�U�=��(�X�@\���4�l��]%l�����pw��&"�=ҧ�`�9����+j 9��E�c��5�ɗheksm�&�����;]_���l���߱����铛Y�;[��Ξ֞����7̄����oZ�u����x�`��U'�f�Z���ugQ�m1�*r)/�H��$�����_��J�+D��ʶ�V�V�^�!W�2 ���{$&ɦ�w�(���l��[A�$4�^�#��:�e�`��=��{���u�l�K����s�T)� _Åp!�e�8�)%���~H-ǔ���3�:{�% �<�}a��Z���N#:㤶�P0|Tq���eM�8ŀ�@2�9tv�E��u����o���u�)��I��1C&cV�yd���o#UX���F��l�_�N�M���e�����r��(#,�SP⥷����_�F�C����M�P�nk
������O\��A'���&��/9���A�g��x����p�ʷ�̫2��^'.�;1���ݬ�Q���4��<#�5{;Am���)}���RЈ�-�����H��7��7XY7���ʑ�� H^�U��O/���W�N�E��=�y6�sT��2@�>�j{���O�7��!vr���nڵ|���yۻ�s㻿݅�d���L 8�MP�u���-�S@�[nɵ�Z�t�? #+͐�؀��|^�)}Y���;��a��D���KǓ���/~�@�K�-/�q��B�eڀ.{ݍ�[#/�	b'����v;qj�JE8��p�-3Jc�V��������s�_�`����2�����ߥ�X���s�������E\~�fѲ���Յ�eo�t#�?{},���-�F3�.x�g�U���V|�n0Gڇ�-�XVB�f��#��S�6��1ֱb�]/���?m�f̮c�a��AN�h+��w�.Gʒɖ�s5h�E0Z�_��/��?qǢ��qf����{L
6�b*L��,ƕ�R�C�ϥT[,I�g�ܨ�m�`�B�������� ��g��mY��bq��d+�x��R�V|��k ��n�q����� ���A%ϲW�90d�F0=��.U .�����H��H���j*	eb�кB	s�G����F�"�DVg
0� �F�35���.]�
���55O��踼���z�����AĎ�����K<;�3�e����0�u�E��X����\��4�1-D�yׄ�/z�c��%��|7C�y&��n��u^.tG���Q^d���-���5'�[]8gK���L�y��N�Y>���V�Tw��ݣ����#���9B��[*���L~ǢK�Zαr��XO�t���@����iكk���N�c`�+�EI�����ؑ�Ү�餽�^i�AU�%��E�R舾��&��4���v�L���,���B�M	�g(;�
rQ���ٍ�Շ���ۈA<��2k���c��*i`t=�KxA}de�n��ɪr��
���ĕz�,?ct��'4�$e%���:�C-�  ݲ��.��x�.{����p��Pl�:�ia| Ӆ�|�|G�����=F]��
���KU��@<o����8��N:MM��&�������#_Б	���{,��L�bÑ,'���s����E��[nO)��Pc�!\^�G�!�1mE�'�]r���`oa^��249�m���T��YF�ʓD�Dn�x�y�[��#l=g���*��ϩ��B��[f�(1˭�r�{I��+/(�(VR#Ok���B�/���2��60�(y��q��,%�e��&��x��f��}�{����]��=e=�y�W]\-�b�Į��E!�p�����B����	i�.��vP���~�18%��,#R�D�h	iƖ��ݾ�,�ey����<�l���ޤ ���F�BY�E�'�&a��_������z��X�>�aP0%U]�`�z��zu{w��տ�ƀ7�yfX�2EM�p��Rٱ����Mxd�'}�3mn/��W?���j}.��Ye+_]D����Hl�z�1�ζ�Pb��&�d!�fM��ٺ�V�o��[2�a�I�8��Kj�T��̓F7G�(�mmrWc�J7�ܡ�w������!A��LhѬk�qٺ�)��l\��?�&�Fj���k/�c�:;2�*t��?u�ؘ⭵�Hl����(�v6���{�Sg�P��$�g6�>�����a��jݑ��l�a>9i�Jq�ťh�/&��6�q�B���=Ւ&)�}�ſ�7��X��{i�6$���!ʵl��J�j}��ՆA)�ʮr!6-��_�-��}����Ҕ��O�<�E����T���<%xs��4��5���a[.s5�|�J���C�DA�-���݇q�,����-DN�fGwh������<1#�kSO����b��h_���M5@�;kkg�G���R`W1�`ñ�
$Ԏ����IL��l�nˁ�	EXr~W�;��K�!r%�}�BmK�8VP�N�1�٩�Z&B�LK���dB� A��~8ِw.�:��6���������w��b�h`�|N3��n����{W�X�7�ŖWx7�x2}�x>��P5���5��	��O1�� ����|%z*WUF�}%ːu�'h2`� hT�]�c�O&�a�ͷi�IG��:���P����Cb���H��x�"Ve�#|������i����:�p�Adq�������
d�ռ)�9k'�<�
̡2�;ъ�t[��L��!��e�Ɩ�@��vK��-u���!�k�Jc?�OE*!Eg�D��;�$p(�e�R��*p� I��~����)o-�4����ODji�mz�R�x)6���0�� fM���C��W�#��s�_�s��^��ÔQ�i����v?��6�Sd�^��� ���'���`_�IUbv2�;�����d4�!� ���mߚB�)!��|^��ظ>E���U?(zX�gasy�"�"s�xP��']��t�й���bqF�=��!�?7_x�X�f��[0��N�9���`2��~$�"���S���6w���k �����ɹ���Ԧ���'8R��z�(<֍�Xi�?��w�E�l�ũz��ɺ�ȥ7�Ym��ˈ�W��<'�
��P�M��S�o%��4��+���ͤ�>��Y�^��|>"o5�2aP!�;��R'�l�����%���įDjJ� ��?
w�C'"�B�}/�K]���4��_ݼƿ�|h�{��pQ�|ب�����Id��H	~r��k����:��ݘ�L�E���E�@B{�E�TJ�8�	l��WS&[�wb��(�)�7���1����^eR5Q�D�!2�����E2���S�^zù��6�s��q��|�J�J���犚�e�L~�W�F���%�U�I��T�}"��k�n��\7>N|���,|e>� ������/@3~(~�u �T�A7�{v������@�^,oW��<��jP��}��(e����!�^�Y9gW�l¹�$F��'Nt��`�ɽ��KE��6#�4�@�p��ꈴ\�^]U���� ��yv��63�B����`C�}����q��F��ff�`/ʽ��;Ԙ)"N6�N�.��p� �<2�z�iI.�f��T��J	�Ύ=�U�`!gc�f����.��<��4���R�x�+�ɒ�>�H��<��:.+%򉜳-S48��n&�OB�o-�^���Y���:ˡ�D����Ie�ުM`�EZ9��wa΍L�������Df�y� R�Ё{���}�I%1���w��dgD��cI˫6�� *��劸0�)���%�}�Bq�N���{^QsKh���+?�
Bɞ�+���3����5rQ���^m��B\%�ǖ��,}�T�O��6����m�N��%��n{.1��!Z���Iq%Q���R�0 w$Q͆�E�|�a�/���H��KL���h[X����`���Hu0 �����L,�!h9��x�[�
;�,���&�>��O���	�<�*љҋl�N3�W\�ذ���kwb�\%����wuL~���z�1���~=�2T�mV���Go��7YY�J;ؗ�=��#r@��-�����2���MNq�Vά8��?^V�*ʿZPJÃ�	��[<�Y�w��ڋ@�!����8�KX嘏���^yb�_���,�O��>�f~�F2�-��4���	�D,A�D	�������1���uY���䊸�����d�<2g+�m7�F�s��Ӑc��͹~Ѣ�"R��b�u��yX�hQ���̆/n�Q�t�P��5�^R!Y�T
(��^��)
R�c�i��zh�V}v���`i�Gu�.���9���i�w0i� ����T�@+��7��o�"��,l��Т�Gv��~�YE�O�"H��A�����̝������H������);�{�^��^t��ZN ����q��	�GmԄh�L~�ɽ��������"v��wyg<�Ɨ8�ԥg� 9{�}㌃���E�#�J��-�1-jq�n1�L�(O�����.��4���9BY����M��J�;}�D��~9�y\��*o�"o�2�g�Z7�na+�����wՅ�������;�u���*@|*��+�>4���8XS`^u�G1ݵ�'�q���ѫ�Ó�9����$lv0_���	�K�{ۂ��+�a�v[�⵰�!�y�w��rO���ݰ��gKn���|ԭ���毐X2�w��z���E�R�3�"KE���R�b���n;^���S'�>4�����S�47+��gR�^Budi'�f�P�%��1T%����%+!�������t��c_�`^.�(��i���=��N����a%�w���C�h�Y)9��)Ŵ�1����"�B�T�T����<�%���Ў�$�7�L�h%�-'U�74��u�u��������J�l�,����CLJ��Ŷ�V�9�G����?�W!���o��.+���9��v����N��o�Ȕ_��̫1�ʥisR�V��#$,c����C������m+��e��x�M��EjZ��t���_4�h������F�,����J���*�e����"S7ԏ��,�h��!&�Z7�ߘ��B.^0z����"&�Z�v9CY��Q�7x���8sk�Ǖi�yw�E<~Yx�����w��Z`�wI�A��iz�sl:H����kAi�Ps����8Nl�l0RBJc%�ҩtss,��L::lc��:�0++�*�Ru�5õE;��h�d�x�ٛ��Mޔ� I_�N�2!�dq��1�yWI$�5�p.~�O���ʴp�4��2�>3��rcV�G���Pb���y��~�Y�ޫiD|g�Ȳ�F#��R�ɈK�vil�61�X;�3�D&�.<\����1oAQhԚv���</�y����J,�����E���KM·ab�z�neN�*-9�Z�S���҃J��8���l%�h6��G�@�/l/���p< ���/����㽋M��H#V�QwWG�J�)"\�Q{�E�鮕���X�I:�g��t&O��16�B��2O��~��N�Ч���*��HX!!�gG�$��$~����(�p�Wjߵm���_ժ�����f$��nKen�Fk&89i�@��"��l+�β}���;�Mۨ�?A��*�����1�*�On!�=������a��I�$|¤߯o�?�d�X]#8��_�[�r6�^��p۟R�M+\��É_�6����,S�Ei�l��Ԩ�nI��wE
��]jC��&����ݮ��x�n���F�Z<'u@��y�Xv��~�p'9h4zgЈ�H�E�!Pxw7^z���MN
� #����(��4,�7�4o`r������=�@�cٱ5T�ֳ�(eJ!~	���)��u���R�BY��&�=���C�i���_p������d�[��i��&��i
���yy�D��6r�,���{�C��%��R��q�lkXu�gL6A��wp�$��e[[q]J��n�\�j�e��"�<3�#�j�O�9i����6��-o�
P4�H�n|g����,�=��$1���^� ���EkJe<#s�s�e>���9's����@~~;�zz�%�nyvS��R>�Y����WiE���"�s�@�TV�p����l�
�U)��.:��9<]X���q|��������kw�_���:c�q֑6A�4��#�c�X%���#�V.]1�U�s�Ʈ����W�ݩ�����I>����@D
�\����g���p��H8��|K�c:e�FG��ø�P��dS�$���n��|�dV$JvX��(��Ym�T��է5~��cF������'�爏�����^&.�4=]F�rP��fᙾ�Bȫ&�H���[
���51�h�#3�f{Z�B-�LP���N�|%���IE}'1������#��	?�DHGM.�웑q4�N�\^O���'�mU��k�g�$�R�@��}��0�p-~���w��iSuvE1&��ۭ�fV��1���,�+�3���O��>;)�������Zl�X#�A�K�A���2��MMo�I��x�����1�x=�,���-��d����-���_�	u��Ys��,�IЗi,	�QqƼ	y������AQ/�R�6T'��B�S%In��(�H�	0�����_�:ݎ<�}�cL��AР+V�w
b�]�)AL���%�t/K���R3�:M����9�`����~��!|�j� rPu���&�?*"�_{��槡��8,
�M=;E�g�U�����=o����Q��Yn>�Gkm-�9�^Wo�%�q�߸��G��-,b;PKdCS[�Ȼ��c�� SXF���*� ۸�������#2��C�	�v;)��&V}�Hx�������ܸ�e����	|+M����x1ex�b�X�j�l�ƻ۫u^y��v����iB��}���Q �"?���z�:^�Aٌ�3q�' 3���=��Ȱ>�[����q��n?�n���}����zhi�-iH���C�Q��4�⧥Z���+b�������o����Y2�^������0���J[C`m�gs�%�����L��`@�!*�ܗ���2^C�2;+��c�(�@kBY-X� ��[oJ�C!W77���Z�j���:Y�{���:����b���`��Pab�cZ��PS>��Rq����B�$
*.�H3�T���${nw�����ǆ�f��LZ*,35�R�̂y��_�B(L=�n��ɵ�ws
lF�eH�0��@q�25�&FKN��`�įa�"9���� {Z.����z���ݍ'|�%�w��F=={���u�x`�x�t�9���5ޙ3���P����@��X���J����� ,\�'���>���1�����E��-z��K�q[Ka S�hR1~�Q��?v>�t�����,͕L �իV�/.,3��}fsC��ѥiwV�d7{�E������ы��&B�X��
�)����7h��t���QErqi-��i�ƃ�3�>k6+��%; �ۖD� X��^� ���R�5`�ޞ�>�� b~��r&|$��O��j�y����:@��"
_]1ax&*�엊��%,�z��ԫlav�Mc#���6c��ȵ��|0,�����V9
�9��Q��O<G��c�M�#�^��A��qXp�r.�������@�G˹�6�vg^Yp(�>`e�$�'D�96#:�]��Xm��_�J���-��&攪IP�3�*1ꨥ�Ҁ�.����z���#=10��3��82#�|�z ᮙ� ��'
%����[�1��,�0/O�2m)����qG��T7\�q���L;ӷRw�nL��&���O�V?ڷbL��χ2�/'���X���V�@xd1��E�C�Y1� ��
\���lu:��vݥ����V��dn�?���������,�����ȷ{3�6g�o�-�R08��}9|L��-���_I���o��)�#A��J^�%i����������kӷ����*	Io���?��ԣ��&ݾ��x^�Z�Ո���,��	�l�7ZC>��v�p��U�09UmH�;�E1G�:~S����l�}8m2�����D�$��\�j@BJ��}��{#�[p�jE(��Pou��E��EIO����^���d������T3ڞ�)���rJ�C).�����j���f����'y�޳� ��Dޔ��Je�3ME�YS�Rm����� A�V�E��Ò@{Zש�&%�8q��r&�v�D9h����+v>�,)}l��o�
�(�C�\ED�q�)~�P�?jh4�&�z�E,�j�;p�C&cH��cI�m>�:j�ܲYG_bt�&��p�
��M6�>����Ϭ�g֜���;���iF6
���hc��>34>*�3���]&v��W�Xsܓ��R1��q�����)�MG�Y�e��->��p���I|ҟ����2��:	{����%~�}L���Ժj�C_����M�U43Qz�JA�0U�WQ�?��moq,�)5PT�,�����b�^ϭ��+fO,�e� ����'l��͚W؟����B&'x���M'[=�2�qw�$Ԇ�� 
��R|��V�{��i��L=���k�0_���q��i��a�7���$6��QV̘�\I\�d�!drݍ���o���G`X`>�A =���K��B��}恘��J��s�?�JM����	˭�-5�(���S�������y�BaW+�|�u��D�I����7�b#t�/�4 ���19�p+>������m�F>/7�b,�2�� 4��q=�Ö�����D#}G/Ey�
��߮R~\� �iֶd�Z�ܴs��Z\-e��R�B������|���]y� �V�I��i ��:�Ve7�Y����N���硪}�w�#�|�n�x��K��BB��=�Ar��9���ғ{���Z����}儉s�g���an�[�H�9f�� �9(j���n�#�G�}�P�b:��4d�����ף�Kp������W_�H�95/�yXl��WG�,_��h�,�����Ug���
�ed�h��x�hܖ�a��$-�$:���6�kY>O�c��Nt�=�g$3��Ǳl�52�7u��Qr�B���f�0*dh�9�[�v���t� �?Nz��=�=[�bN�;&Eu{}��Kf�H��,FDƣ��\�% ��j�{�����հF�ȶf�cs!?��3mv�[��A=ֲ��ʖ�߳��h��u����*X�ᬫ�}�=���`����)�ptXc�2�t ���6O�J��}Y����	���)�`�w�"�w�����~1��E�Q��[�Kvz���I��$�Ex���R�k1�*�I�C.~���	�p���K���x!,~�\=��{�9�����Nwr�#�%�%��C/|#W�f��m�5�36�̟y³�Ѝg:��R$�u�6y�=ݑ�[)#�`J_`y��ѹ�
���c��;�iÁ#�DO��?u��.A(Y7U55lӿ��+����
�\}�%#B��rыr���m����8a䣬��Ǫ舶Vgtc���ෳ��T�/|fX����2K����}���JJR` ̇G��q�х��NW�vP�f�/���ȭ�e���/�jmcNe�|Pg@�]%f�ω ��5n�0��>�����5���(�-��3Ί1�$%O���
[*{���j�����A%�j���W���8���z� d=�ar��t8��~-z��ԡ��y���#�����e+�1ҧ<�TM��qZy!xE\�uZ���/y�/B�Y��ظx!�DJ���Rl𸩟ZzO��}*(��J֨7�;�ʊrim~P7;~ V�&�hF�䰾��ue)�� -U����a�a����7��4OV"�� T�z?@DL! ��!�J�����*���68��'�O3����'Y6�a戓�������ܟ�7�~��2�2�F�a�37��8m�7	I��5����R�t������i ��\^"�]f�L��T��s�A/*	L�?����h��� >��������	m4���D>M]����{M�L!4c؊jx�Ԇ�>�CQb�����S�hM��9QWS��kh�D���'��E^=Aq�og�O;�4�'������" �)W���fY�M��/B[s|D��u�L��҈���N�CŦ�Ma���R��\���ewQ����,�HF�}1�(�M�D{#)o��j��x1''�Hf,�����zFV˒��;�� ��d�ot�/y�G�T5�X��ZP��M�v�\1BR?�[.�b�|a������)n�,$��s�l<n~����ڰ
)n�bɮ#�Ǥ���jKH��g\W*�%mR�d�x�det���zSz䕨���Iݭ7�9����.
�����e�
$�BF`MA�g�0Ը��I[�t���-	��ϼ�&_�����H�h�8t�,n�i?X� ���2��ks�hc��IAK��2s*/�%k�Ɇ���2�q�9փtr�y���uZ�@s����p��__CSp�Fl(m={�ߑ�v���$�k�f�_���E�9��>r����}RSĒ6��: �>�u��m�.�O�V�2�Ԝ3�<a=�#oܝ��~�!K�&��Ҵ27m��]1�^�8��U*���l��1]kD���a:�ո�!`saLO��S3�Q[:���ny�O�l�u:����>��ҵOrc�w�	w�[qaC�L@�j��i�����1�K��|��{bh�u� ��%��Չ��M�ߤ�k.���]|���+ �8a�º�@|%�G�x<r��;���$�:�	�DfO5N���e�:�U��VȊ����4d�~_��~�����eO�9�����D`���7_���s!Í�j�@.t|�<�b�	&n7��1yQ��]�X��ПT��0���	�����és�;ݿ?�,<���[���!�d�kf�ʪ�J�'܋��O�L=Zt"\ר�������ބM7\�ՁY ͘�h$=��x��nH�P�u��{���}��)�~��r��>���xLj(��JE���x�`��ܬ��x%!�ޚ��1�P��u�+~��{�@7G�@�	ߺ0\|�x�sx��y#�H�x�^�y�|�쇠o�+j~#���ĎR�T�"��p�uP�� I}�Hx� +���+���ZFm��6��퀬�qp|~�zߦ�0�1^��a6&�B�z�	7�����s���x:�tS]Gi)�Z�����߻3<pA�*SF���Q鶣#�?��]�}�m�y����X�����'F/(�@���FiP��^O'اnϙ:���.,2èF|! F��I��˅����Ap#;���"V�0O0ާC&5J�}9�= ��f	;����R�J�78ٕ2���
-�@za�� K���4Q�V�Ev�.�0���p���kd���O��b��'3E7og9/hEn��z-p��m�,���E �_�(��@BE]!7�����7a6�ZZ�mU�b;G�("
'Mm�`%�K����w/�W5��:�Ok����f�Fi�!Ά�����W�����i�C�\�'�"/�f�����O:�O� ��}�^���/�9SFG��L��N&��<q�1��<dt��Z��r0�?�%���-�����j��hsӝ�A��w�Bнf`�:���Z��ɲ硵�k?L0g�����i����sQ�M�A�-�H�] �K��3���R��`ɇ5gr�t p�K�H��p9r?�|�g�c='8��;Ƹ �Bo1a��w�5�]��\��3�a��\e��m�솴G�wBRA:(�ԢG���*�U���ȭ5G�\$ٔ)���=d��_�,����l��
��W���*�W�p�018]Me�d�ڌ��f��;����-�4��f�d)���T�^R�U������@y���P�`t^����5O���|c�����ڼ���<�q!�w�1m|���CƳu>M���~Fdeg���5rYmB�"��o��
�#����ߌ͐�,y�f<��9���w�'J�*4xہj�g@����?��v�i�g�5�=�0�A(V�¡w�L��
O�-x�~����fu5��٠{6��9㛃ĺ�*d�j��ݙ���T�������X��������^$4���w]U/v��)����=�ćr}D�,Hn*��ee�9�n�O�٤�;x��y�R��dr��Sb�-�X�U�G��?͙<uK,��G?A�ӕ�5(SrkH����(O&m�+vzO�m��.���ʄ48���t<�>����UF���*����u�߾�/��ҬZ�~��v]���o46��J@����UN�|�9��wM]�\3���M�3����FP�`G�;�8�ߚx��]:�S�&������ � O $υ����.n�4NÔ?�w�'A�m�"7018rS��*`�Ԗӝ�-�g�޹!.|�A7�R��$tb����}n�������);�S:<ڔ������svFR������Cgi�o���;��sC�1��˘�o~*�6Z��J�z��c�l�Б�<�o����"��K	�m;ի�t���xV"�,��XV+<��o{T_�j���S�1�e%S}�(:%��n���r�P0ޒB��%�6����h#R[�?��E��"�Y�!����Ω���TǢ��}7�1�(��:��F�ד5��+|���$f�-5��Yt��*3�m�6����i"%O�6Mw�j{Q�u�]'�>���G�k�?g0x��U�'���kCwx�f�v�i��m�,�&��8��k�<Ge�t�(-�n��Ku(�2���R���_	E49�q9�Oa�>ߖ����K�Фy���5�S|e���F�8��蠯�˙�0���D2��I��d��4�����`l_���2�T=|:��ѣ��vXYS�����k�]�!Br��R�K؇k("�R���Uھ�y��?#b�^<��R2�=�$�;A�}�����
�iԜ�i(p�/ 5˧;i�D!6��,=�p�5�0�t%���m���rfkp�[`�'�L&c�"7�C`v�׊=kj������2��"E��/��e3Kw�T�_�^)X7*O�>�K*�7��F���~�:ߑ��HM<�j��"�S�IU�I����!�	���4\�lu���h3糘EJ��,)�T]�]V�/�kF[��`�=��>N�
����Wu�~�<r���m�c�$)m���.~�=�w5M[�G
�ޛ1�n:��ܜ�f�/�Ɂ:=MHE����8���VeWj�@�,�!�#���
�lv�ښ{�j?�UN���ӡ� S�A������{ql�Ϧz�*J'�l5$#9P�1˩���/R!hW�b�t�!�����A�*���-��Ћ7�K8C��7I����(�&�!�~�R�.^��sc&���}�m�w4���~B�0̎�<[�H#IQxRH%�H>N�U0��a�j��W���e�?�"�5�����F̗�a�t����asB�
��B1S+�]�7���{�FnIڧ��b��ĉ��I��[���k�$R��\�<n��q�꼌Z��O���I��w/?�����)A�8�]�;�4��''3r�j.V�MB?�2@˩��ԓ��� C�)��(u9��Ufbm�_�֭qD,� ���d74>�C�n6���HXǼ�V�uԍ�y3D�nrbڭ��ne}8p	kK)����bs��&�bQ��E ���)Ԝ�ے�k����{����C��Q�C��F꘴پ���j��+��O����~����͘zR+��9�W2�-�Qj]�l٠4р���WeI3��X�p�Z� ��6�f�d�:��hJ�)q�m��"$�j��h@��_�F�y,�O���0�6|/�'dU#�?� �V�Y~���_Xw�n��uKS��7�;R`�&�M]������A���ŧ0�:yw��gv��^�����T�\��Zl����^�$�cq�0��K8���\�ަ����͢{Ѿʁ���,�kZ�y1`LO0�d>�y�vs�T�Q4���|#|�}���6#��m�n5�~���!{��3����}��E#X�p�UU1�&\1��b�	eO=��V�=��]5�?L��Hwe(� D;�ǥ�̬�3x�(���Ȳ�q)߶�Ͳ�o�徠�U �"��Ofw��Qƺf2hx�,�`������Y	�ybqEe�*��r�9�31l�uP��Ì��P��͗K7DI&=7<���l_�Гm8�o�Y�#ֆ�:�s�?M}����\E�(�ZVO�髟76�+�Q�|r��l����e��2������c��h#����i��k/[����Lc��c�N!�x_�!}��#<�u�<�Ϲ�F�RA�H;�%��`�����y��\l&�N��k6��6z�����ti��v=n����< 5t��eW�_a�4�I܂o�Jo���ܒ��'�f��f����Gȋqی;�]�7;U�m�t%�h�;�(���ou��"��.�	�q��[��bR�J��+���u�����*�|��˳M�0��|U����eH@u٩��w��U�W:E��G��h���K��d�s��rT/EZƢL9J�T��.Nھ��]�����~�p�˖�"P�o[��o�g�t�qಯw�I��ė����j�*���/>�\��D�'|cuX,��vs�[��
M[�h�]ڝX�Ř#������H�%bk�򌦈m�qO ����.��9�v{Ny8#�0\�AU�������o���V"�$��ߙw�[a���R�v�E3��<Hu�`>�����x���װ�����3�#����M��"�Zi���{�G�K5��l(=nu��hz�Q�<�5%�[�=Ou��ҫÇ����X�)���?;�h�0�:J�D���$�� h������.Ӭ�q���A;��=���W8Y���š�{"7�ڏ��F�Y�b	D����G{�wj1@�~�L�C��eU�����:~�0$��%Y��WAK�`Ɛ`H�0���2�g�|e��%o���
F�V�"�^f���:��Ľ�%Bs���9��%B���H��9eno�Y?����0vo߼B�uشǲ���?����0a��c/�d�;�����>�M�-ܜ&>+ d1N�-��hS���D�H`�8�֨]�?0�������."t��Gх����Y�Mu%[��o��U
��|t���iJ�v	���w~���s���}� D�Z�����f(3'�3o0����ΌC��kBoW���	_e�"�.R�q},ջP�"� &��w2{5��Ci�4���~��Z��?L��;�XU�A �\������;�ّ�ha2������ִ\��!���HPţ���-��c����y�f�m��8���V�J���c��w�^�q�dM��E��J�'�H�q_b-ӹ1�&�F���t�"�����2�S�,�@���g�r�����+]<�
�p�<2������+w�u��K"
��sUZX�������+'TB�[�/���[/"��-�����Z���~�$�b�C#���<&uHQG�4���J�"bn�t���u�DGP��E�eSs39���4��i����:�^�������P@i�eL`��ܑ�޵��-��]���0S`�6b��Z2k����s=4�<���uV�'UZ��.� {�;
H��W�mg�!��
���$1P?gZ,��}!6�1�Rak����Q;D6����A��,�4���/Tsk�;�]�幺��M���(t'����1M,��$��� �B��E�=%�aM����8�������҃L|S�i������u�O���w� V]�9r���Z�热D��lT\���>��_r���	+9���3���T4�}��N��c���cA�Z��g��E�DE1g��ؤ(��70� �w�k�"7O.B| .�����Ɵ\dMs H�Е¶�����,�by�O�`�� �h�~h�zG@�R�aX �A*ۯ���P���B����q��\2��g����QUi(�	��9j��
�r���������A��d�%x���Y���Cq��Ϗ�*<�۽(-�U���f�:4�u���
r��G�(�n����.�/�Ux�~�,F��&�5�[���EP�[�	���T�a������6G@O�K>�V��ڧ��v�:�Z�����qk;������.?�-o�c��do&��"�QPY��Gý��>��(P�ih�W�& �u�~CB�U�%i��}�a^1U�^ֈ�>
V2��B�h '�-�u��ISRL��n�ϕ�k��f4��V�\DC��w��M|4�H�����'^4�G��/����.#�J��9/�4�fݔ'{l��َ	�� ۂL�Rq�z3�x4<�����a�xh�����2cAph�YK<��C�0��{t�>��s�k#=�0�5x�CP�#?�o{s�SyI�ř�N��`O�K$#�/8a�!�M?X���{&/Ě<Ҡ43�WR�� �lR���Pw����ݺ���0�5uat�$p��V��)e��E�����j$�xpI6`�a��Z2q*��] �o������P++Ey9.U�S��"���[����h�O���M��� >�@�1�z�I:@�9θ�A/r-��(�� ӏw#�zk@��?Fx��1<ӜSg>�aH�nJl���TIX�Nc3$/�"b��'��VÛ��(q���I����׾��P�j��Kzİ�U,���׶0���$_ĖW�����Y�ĳ�m"V���F�H�l-=b='\���e$Z�l���{�j��,��λ}sk���6As��Cy?�X-Kͤ�1۳��2>F�MN��� ���}�������Ȣ8xqQ��=&�2�tJ�=ϣ�&��9��aЫI�&��n�V{�%��P��ʝ�$�6�d&*��i×ęM�#.�g�3��%�J�O*��"h�ؕtLc� pdk�r�*{+��5��.�����k�������b�%R��A�S�N�>׉{#8�fNJ�r�%^�c�8��w\��<���T�W�B �h	��|�T�^�Z���)�����|���P�PE)�^T��0�8��z���:F��%[f�|c�k����w2!���8pH� Pz����K1��x8u�R5Z� �@���X�G�̕Xy��$=�2(�M0B�1����.�@��������=׌�!�����m$�
b3]�r��e�'ܡ��o �mū:S�A����FM@�ɮwX7]c5-��ҏ9%&}��e�b�K����.����x٨��M-�fE~�]TP�L�*����$��ffi3Ӓs���
E�6H}n�Q<ϵOeh���sފ���f���}dL�� ^�*F�Kڂ�{��2���ػM�ee�?�>�~��$'�t�ԯg~�e �P����7"oAcM��H�L+�q=o���� �oWҵ٫�F��W�vD2�M:*�V_��N��.i�|���Kw��$
g��0Ug�-���-�/������7��҉2�Ÿ�5<ꊏ"_Em��x#���Jp�ؾY}8���F���a�|y�|T�?\�P� �cX���2�,F4q!M�>�" A��i��hOi�x�0�Wz����T��|�-�߹)�5˨h5�e��az?��t����@'w�'�|�SLa��i>ތ�I�)X��%nJ	V�#���U����(.n���|�<�N�+������c���Dɞ�R)e{��{�5#m��Օ�Y�gV9�����}iк��ݓZ���]��QW߳�`q�nۗ6�tp��D�ڱy��\R���˄��Z�'!��^�:Ad�<�,�O2�XMB�fj����1H�������������uo�֏O�	����lU�^�y�ńO���Hᡏ�5�_q�o�!:�l��bĕ�nM�^4��@{R�	�"L�'�N�����[�W��ٶ��+Dɗ�sQġ)�@T\��׃P��RN�>ЍN�5wX2i�٧��𶈤�M?�ڡ=��l�x��I�ÿ:?���Ù���j��u%�F@e�D�.�jh��=��҉�M&N�����'zi��(�����a�QcoȘD
�4�,#��sA�f9��<���Xq$�)���|e.j�c�o�)��a�1��E� ��m����~e"���7�,��	Q���eS�3��/Z~?�����;j���n�µ��k�P���!��J�u�oE�ll����#x����N�}X���v��jb�vT�ȉ�/�>�n��w1��r�V��ⅱ�"\{v٬�L�9+aI�4�����l�������}4ӌk>P�!w%�Šb��`L�w5AL�}��6��IP��6%�W�#��7�p��hI�����އ/Bs�p�w�����%	�R�V�I6Fr�>���?ДY���OeM
��p\�[�K�~u�	�4�y�!�[�L2�� ����d	n𵂙}������2,�Q�C�����m��1D�9�-w���jO%�l��?Ќ�޷��m��}����l��(ye����j��[��~v0�K�.�ÜH��Lq��V�����(� �|�y���9+a"��߭���fp�5���D$���F:�x�M�pxqa�����e��j�.T�G�� â��}��d ��P>�:%
ڱ��K~PM�
��qO�)��.2�,�¢����?<�S��"��G�B�)��
a�2�B���e����M�Ӄ�����i���Nc���9������Y�FZU�	n%�uL�iOBG�^�6�y:�yC�N�L9i�\l���l�ڡ��xCUB��4(͑E|���`�ٮ:N������J�f(z�CP� �x\�66�/X��Ys��Է�Һ�}�	�i��f�we8J��F��b�Rw�)�2�Ay!��ѽ��j߿#�`�G�������/�R9�@}�
Z�2�3g���_���õ�00���5�xj�.fR,�R�8I�[*��.\[�C^����|�Fn	0�bHFm�b<��m����5
�x��)!׽��6���w�Z}7w���?�RS�9��A�\g2�*YV���` ��Ij�\>I�I�Y�>����ETH��Ļ�S����-ɝb�{a��T�Q%�If]��m,��A�W��2����j�_���?#Lݣ��Uh=kG]W����$�D�:2`}`�2O� �m9���WV�d��ϝ^J��)B�i���!�ä/yl?vXu��k�!�n6'�at�I�u��z!0��?��R�i���aV��}�^(3��~����֋��i;�`�e�)�۠����)鴯���H�ަ+�|yC^V٭Z�u?:?m�\�	�Ks8c6(s�����.����M~ �}D�pN|�:�O_���|m��qd��#��: Jm��T�b��>e��z~��F?E��?����ʰW<-t�<6'@��	�+9�)飘�=����ܱ���h�����:�W��|,���T/�Y�����g��u��|�{<� �aؘ*��7�B�����d�c����������ݤ�@<�B�N��8���ȕO��:�I�iQ���x5��3�V`K��ٝR׷�C��Kg�I:�WF�/n����{%Ց�-��`�� ��ȋl6>�9/�E\�{�A��>V��j��nj�/���~�~��z��Rr� 5��>Fb���l�#
q����X�.�̻{!�������������$b0��^��p;�o:4{(\$�[�Z��hE5둡z����b\�镀MB���Y*��=�=�m��[�vv��ׄ�h����J��7��젟A���mD~	4-�,76���wPy�hL���{��S�b�x�	�Fh���s&s�':�~��!Y���)��b�'��{_S��'ߢ���;�X��Lv�>a�s�y(MN�]QE��3ݺ�����X�y���FW,U˫�ga+3"�Ҵۈ5��[b;��Oݠ�����4^X{;H;ڠ��7C$N�2��~\Α�y�9*�ۼ[_�u��)�|`�4|�@#��؃��o��|�C[l�vztxtS·�@t��Y���?����]�`���<��V������2�x�m�W^
��Bq�~��s�����5�U�[�^]��ZO?3��ۋ!�f�Q#� �Tp����B6�]�FeԟQ/)����.Of8u�b����<�d�}��t�%�(3_�P����1�,������^�ZV��!���e��KN��������
t=w���B]΅���.<M�2��K4?y�f��ߔ�'Lx,����
E��}+ �e�8/ǋ�)T���6=�9_��1�����M�~:<ױVѶI�?���t1j�1KO�y�x����V�fJ�79�3��兂�٭�S�q����̀�;78�9�]���!��(��ٗ!tI��9o�4s��G�Cd�qQ����7�����ߛ���U��K�K�\�O@���?&GG��F8��T��_}P̨mc�jsJ#�9�e��?�~���F?٠��A�/��U@��A�(}C�~��R*��l���js�g��oA�^e
��"h�c�� 1T�X�z$�١&�SAG�k���;�x�<��ezt��y#k�,�U @4��ތ�.yGf��#@�=r=3�
�B��̗z5t@N={�''!=����T�/�wT�΋��3p^�f,��o�o���p}��R[��[t0fN�nWU�
۲x�F�d�.fV����b�H/K�ý(�i���ӎ��_�1F�U�Y�/�[iE�}S>=N�l���̠S��)�0��D$��	J+?iͶ&1�����p��Y}�M|����P��?�2�2V0v���ہ�4�I�j�0��� ��![�Qݣ�	=�#P�~H�E���x8t�;,~�:�הu$�Ķ˄�ZW��B�<©5��n���I�ϡ���̕/4�	�-�USZ�h$�tP`᬴Z�,�����)P��6������e<�&�}�ӝ@�F�0�$�Q�{���!�46O�����lZX�޺�F7��Rw�X�S3d�6s��Z�u�Q*�߿B6�<��1��\�sBD�w�V�J�<�TW�l��o ~
<�GkK�	e;�9����������W�r�v�~�3����a�9������U�\�L8?p9�d���A#�,�X�"nmf���q����;5h�:�-Ux��B�'ҿ����u�P~w�td�����Hy]C̼��Ԋ|DX�	����5��$�{�İ�YN���']��Ly�fX*�eY����z:޵�Hn������*�i���@ ([�ٛԪ���RA�0W�O�PJm+�zW�zF�%�n�U&�EV�Um��W"�J�+`�G�c�QL�(�_PR��w>���C����u����K�pf՗ZNQ2Q�Cs�����r�\�ha���Yӄ��u2Y�i��F�c4�+�E����f�������I�*�d��Ξ��*%�qEZ�j�U���Foc?߫8��]��[G]��Ot���s�F�����|��]ٱ�,� ��WSѤ��|��|����M�b�rl�0�i��7��]&_���RNkl'�b�J�H~\)<�<��Z�]�%�{�aBG(���V��BoW��^I@�����:���0�ⲽW6�c>Q���: �,�
�g1�dˊ'�<k�1d� �L�������|�
��R?Μ���GI/?
��F��CN��ei���ڴ�\L�P����3��7F�m�b㝄���h�������G�g��5��~�t��J��d/|��9�"f:c�/��/-�w"���[�0����|GedbAQV������'��w���|xP��$�~窫O��gw� �u��Q�3R�.D����uU���>�虡 �h>2)���]F��� o��FXĎ���a��􋣊De�����/޳q�f�T�z�rF�:~����a*�����U�W{OĚ{H]��zu,��S�,u͈�Z�[�.��Y�V�*H�TU��Uy��yo���93����4�L��_�iϩP����g=���$jLGg8����bX#d�-Si�O7g��՗Z/�����A�K�`�H���:��Lk��Fo�T%S�ȕS ��J�Y�G3�B�����mG~%Te�x�h��$a^�%�sP�4p%2�f5*%�zM{x��sw�Ֆ���k�۽]��J��/
 w����t�m˛�ݛ|���M�2C�4z13]��^6�I1�:; �tJQ��7�fR�>���/س:�`��ӡP����p��r�˻�Ƒ9��0�eV6x�h�������ܥ�x�Y���=˴���R>0j���B��A"�h&����&��>�'�@�7��8�L1��%��ƪ3�{�#[�Ѐ�	��3}���gd`���?(���ո�"'&M�G������݉hR�m��	)��|��֍�M�9?�z�%�4����1>�V���<m�.�������#c��N�:�A?U'U�	O;{��G����e1�����($VOg_�u�Ŭ�����ə��Iͺw�隻|x��O@����gG!��s�&�֎C	Ƣx�y��]���D��|��Q_pe����w	���bS�����A�R�΋�F0G�=i ��@Z>�꼿��Z��u_��Қ&�!��>�-J�Ǹ�u�bh���<hC��<Wd��F����p������R��-b�G��t@�R��z�4uLЦ���}�-�OD�j��`|q)kó񩦬R�����cy�V�/7P�**'^�돾��Y؊f����/ʅ��Γ�ELU��mֆF��AnI��9���x�v�k�������TZu�����Q������$�*}��?�6+疽b��"��-��WsR�A�8�nz�[<H|~S��M;�M`�[�.�	=,T���cA�{�դ�$n�Ͻ�yޕ��"Z.�Ô���3�G���ف�MyEm�����R �)Z��G�5�X���Ɗ3�)���ď������j�.~��ŗ{pC/,�C��a
z�+5R.���ztGG���s�ew��F`�C=·���6��5$�/�O��%c��5��������hGs���3��\�;]�z�T�00�.�������~����S�$���ϊ;�0fi�4��h��3����S�vG�K��ȟO�N@j�rL2�n>"xȑ~Î(�k)��i�8?q���R�mRZ�2��5��"�J����[zw|�OP��/��Ե�k1������qC-�gSر�Ȭn��DLER�$�%�b��mݏ�#@~)�Rqk�	�|E�}�8��R�5I��s�!zA]�Q;be�����kd�u$��M� ��!mߌ����8:������N!Mh{�D���mY��I��&��	|��*mW;ya�C�ɯ]���|��h�8b�, n�T2f+��u��]��x�r�6b� ]9-)Z><��2y����� _�d!@bZxѳ'[�C��cUq�m��q=i�}��g6$������қ	�����y77�&�-fR:_u����� ���>�'1�����2αw\�����xi#���Ù�i�k�gQ� �Z���o,�*���e�}��X�~jHα��V0�a�<���q�V��r�F�J�IꙀ ��>F ,PL�F��r�y��wZ6T�%��g�}�@[v��'�+���$D�Ɔ�m�ǻ����:���S׋}��֗�r�tD�%d�1ޠi��?%�a�8rW`�BaX�&�d�F5� �,�t�g;���e�a���)S�ײ���N�<��!�s�L�,	?�x�$�i�}�,���ߴ!��oT���gڀ��R�7¾����m#8Q�5es�l ���;zA�}��lv]�8Cn��h��!�$���H�����x�� �M�ȆK��?�R��0��`��0]���R���'��<ȃ� ��ˬ
u�e&��F
�t����KX�y��Ml��ܪ?K� ���N�/��e���UkX�Ֆ�c��$��kn�X����B��{|�ʜ��Q���}�7��#l8�lI�������$��e����
�S}�93x�y����ˣ��_Pl�!� K���U)��1����1?iݕ2:.Խ������_�;��(D\����p�4�|;�3��+�G �Ah��s����d4����ӳ�Kk�r�Z6��}���Xڇ���Xy�~l����R���+}֒r���2K�A�(��摷I��o�*o`}�M�)��B �
�7r�O=���UgJʸ���Z)�W$�6�֍�i�U�̓��Z��)C�8e�����Ό%D�jd�Ɛ���!>��\�U���ks��x�bh����}2��W��1�yWs1����Tp�/����3�]n���
�\l�p���!��o"l������t� |�O��>�ܫ��N}�$9�/^��u6l4I�m.�M·�$���?������@�!��23�@�x�R�@���AQsmRf��wux
ȬO4Φ,�ݜ��q�h^�����|ٞ����Ւ�u�%JD��F�p�aN��U��NJR'�:�c.���aiY������	�3�QW!�I�H%�f�
���u��l6���h��zn�]���[˛�s�-ʴ�����e��$���g�l/��E$�뼙����BO�AgGS_j���4���o��R:^����̧�(���&��p�ӟ��Ӛ�6���,U���)�r�2>���t�+���K��M$Ia>������Fi���|����+�!�(˾Ed��x�g�N��ח` �e�S�/��AiX����ڣGՁ<�SR<s�$�	f��t�	ڕ��S�� ܞz�ȇ)w-B�r���j�5\*�a�:�T�H}�V�!���r�Ξ$B���Ǜ�=�\���&�]\�|��P�
����̅취�}��?Y�1lT�J��� �gl��!r�dx�;�-����:육p�jы���q�;�1��H���aQ��Y�Q�(w��g��S�~O}ךk�JΥ��k��3T@RZ~2E���3S�Zҙ��Xa�[ey>���m]"�q�$�%6X�0��0�*����ռ�5��������;�u|���H�쭽�T;q�[�M ԭ"��?��,�%(�3dN��75�vX�����La�]���~���+ͮ���l�J���7����"��e��!�o��}5�R��)A��l��S�Gy�㼱���(U�KM��oإ�~i�y�&��J��g%��'� "㇮ԅ)�A���}� ��9�)X��(�����Ղ��$	i���1cf��]re�Ms
�*�gE�]?i=��(Q�x���8���J���������^��� ��*�N��B| 	�c�O�o4=�i�/?����y{>�����-��c�J�c�"���&t��I$�P���׫��J�[���BM���|�eG��JF,��#3�.�>��{���Wg�AF�;��s4l��~	k,@�#�;���&�r�����
M���i�Hzƅ �|�&��U7���poG�D�?6[dO�M�\~~N'�/�:b�qIb�5߱Q�~�%@�װ27��������>=��f�Ș/�[g˃i�+y{���Vh�Ȓ�?�;3���`��;�d��N�d鮳��ӵy��S����e���Ϟ�,�{y�5�o���n��]���̫a�zA��V%�*�Kn�v��A��s��7Ж����cg-��& },�KmԼJ~���k�,$�lhX0��Yߒs+��Q.\�^M	�%HL*�H�ax��t�챇5U��	���TI"_u<�6:�Mt�v���h=�G�i~�&)�B'L`�.����_�c����|�� �Y��f�}$%�
��_��\�?�r�"���R�H����%K� ��7��7e)������4+�̛�B�V0�7l�w�}��fG��� �;,�ܮ)��<���Arbr�@���)Do�.��nO�����F��Qڂ Q�SӽK͟Q�j�8��ݛ�-w�ߟN�E`
�P�e�Z�q3�xum_z�)G&K��{	 �J�(\����u�����Y�H<vǩ�{0������I��+_v��],�}`�$�Rq,�7�Qf�g���#=��^!�K�J��Ԃ��[��u<o��FUY��s��lf�v�+��<R�\���eߵ�,���w7ϫI��n�@�5���k��b�N�)5�a�F��P��<?5�d�CP�k�%`~�?=�=���&�Ey]�쉰�7҄V���&�Ofx7���9Sd8;�T:@|9?<S ,{�1��%�S�r�	�zQȷ<"�*Hr�?�j1��%r�Loϊ2��~:o��iE�U��Q� �\��/������k����2鿞V�o��J���f���1�ĭXI�CY!��E�s^mO)�o5S�>���|��oe��tn��������Ƞ���FN������s��� ��3�S�hт }�>B��3�R�ܪ.�C�J|�ѝj+��~��W\L<$���qn�8�~繝�t���W�(^c��ڮ;�Y���Ƹ�Q���Z�lx�(ݝ�?�*������3$W�줊�x-}`_v���rs�-�0���P��w	T�t+�gQR��@ndrd���|~%/"9�;�Q���ώ��H0����LC�;�����S�c]�@{����Vur].b*.�&�G��q�ҞBg���h�����A'�#�gv���4v�q{�q���XEO:B�v|�'��G/
;T���v�0���!�Uc���ݻ"�@`����>��ʤ�eZ�q�� Dt@R`��c�L������ � 75
Xŀ�1Y�V|\� )R�(��HbԽ��8��y:Ҟo�\�מ����7'30���D �F`�WRD�R��r��٬"����7x�5�{�ܞ(o����q3���nI��^���ǰPvν�&�V[�)��� �w�ƣ�Ͱ�XX�N�|���4d��A�ir#G_8���$�a�6S����Û� dkiq�PU�m�ղ�n�&S���:H8�Q�MD�  ��XˤhLr��)|���+=o-��ls�Y���Рz�\��j�GVO��3!}�FN@�n
�����<F�E�r1Sq\+d���K�G���G���ճ|����@r��b0rc!�!�C�a����r�ِ��n��;M���|-wI9F,��h��氋�}+�\�k��:��`��I��z���,��i��x�NP�#>
1��(]^!�Y�)'�_9�0��7K�eK}�����L�E��B�;���㘩g��|���d�̙<ʘV�C��bo�fɑ��-�kh�{�������P�F��:M��I��_g���6fg@�k�\���.�t��M!}�[��ձX%2�t��'A�H�A���6O1���5�p5􎱘`3Y1D�[k�@%x�Zs��OL����^����i��+Ǣ ���0iښ��X}�d�',v�G�0���Z�����*Q��C%�֐��Du��US�{��y�n�9-���2_��m�o4�/�J� ﹙dr,t��Z�\$kN-�M|��2X����jHH�@�Yg�Ϲ5T�g��c_]��0w�qhw�X/Y�=#��bX��;.`s������_
�u}1�>���S�����	���� .��}����2�>���uZp� �N?����kƎ�Q ��PW󠫢(���h����i�;j��t�\��P�7��	�O��2�I3���*��J��{�)n<��;3�*Y�o�v9�5���]���y�A�:&��o�=�c�?����>�I�]�!*큵��0����5%f�Qi�:K�*�\�I+$�ج����m��;/� f&�Cm�+����&G`i��8Y ����1OY�ի� ��9e�"�[�pLa��-���"�p�
�2�G����5��x��ɕb��N4Y*�^��	|>�ufUCxv�p7A�=Y�-���Ղ7�A�+��1�:_���gf��Ȭ��k�8I[���J�a���w��mB�5�֨R�WAW�Z�r~͜�&~� ;緵�}�VI��:fG¬���/��Q\ɜhT���jM�#����1uI�P������}��5F5p���{@��#� �טM%�\��񪬬�6<�+��������f��o��1j��67�@F�ǹS�/?a�8����GέϳgsQ@�l��Zs��EpӔ	�ϩF�!b�k����Sʆ�)@��wz���d�Ij.�#�s�@}y��5�����æ -%_���o.:�+��j
j�H�p��!k�;G?&�3��x�B��~�\+ظ� "N���E�҈�(3$ɐ{�������;	NK���c�(5-DL�I�Qm(��U��A�>�������v�VJ�#H���u+�x�9�i*���L�2�ʾ=i7Ե�qu8��2����%S(K��Xh5�M��J7`9���_G6
��j���]?ǟ���mF	�����M�R��m==.�:x��2��n��6���5A��oD��=�V�&4��`k��t&̰m&��^��R_k�껹�vut�Ώ���<��Q��s8�a��VvAU��s�(z����[Ͼi&��m�VR��Ԛ��q}/����(�W�8Y+��"�D�Khޔ�Hd���^�N���c�!Ay�(�|֟V}4)!�֣����-�B�Q
ܮ󋤻���5�aw��`���L�	��J��q�����K����atzbk���㹫�-�)��'�e��|'�7�Kd���K��T��|j@�'�����?������1p>\��4ȅ̡��]f*a���m��n��n�����:��G>�D�����K���K�T�W�!`K.@۲5���%��Z�x*I@�O���ਏs�<����	�<��,v��\���p�?��ۃ��߃���e"n.xs�[P潦Ro���V�{c��4_������H�]����G�� "{|�C6�����G%�R��u��"�<�a-X��9��$���X�l~��4�P�u��J�\���b%~� �-���q��#j�uF�ȖN[�W4�U�̜���W�>gp��pV�,G��k!0�!�:���'�8���PS�7��!ň-�jM�p�	�I���UGGZ���}K�qe���+q��%G�]&�p�tn�XI)��5�d,�p�hGGa��Q�8S�b�>���k�f{d2���eg4���Z�~��Nm�M�
����:�߸F���BX�L̎� ��cpF�u���z��]͇DՈ$]�H��q$"�2MZ�/k3`:N~��g��k~�����[K�.�Z�%����N��v�1t�nR�e'*��O�9p�{�^
8���n����/18ӯci��]���¯�d���u����j$����%!q$�w%��,;��q���ΐ�nA��f!/��PO��sm��aa����Zz�7�oAc��G��V���đ��B{��6�p"^��y�C�"w��[��g��9J���;�&<�_�>cfs��I0�\Ryao�gi;%�h��3g�#�e����q�l��> |��g8T%�n�b���y�n����^hu|��ꯨiZ��b��r��*4�nv'�����6��߰2���d1Àr��_E�����je	�_�w7c�`���M��[����}�N��v/*
|���@�ah����D:(����Ye�Gge��u���$�z��V38�$G[��9_��4�v�5�"]�=���F�� g�0d2�%7��e� t�����S����c�S�=	9�R�H�ْ��׹GU|l����E�Kl{����w?�p�z��6�^�Q+U�cAQrq��G�=Ju�.��Ԙ�%����d�l>^��4�l Q�5�!��X�|������w?�O�":UE��Y��}0|4> �Mt�� 1E=�Uu)�aڣ��d�� 70�`�J[<�����mP�'�M��Uje^�&G��e�'m��zc���岆��jɩŌua���,��ͩ�%6ڦ@8�������[��v ����g���B;�D�'c�]k�l��J�=�XUW����%1,3py��-���Ή���U ���0Ӑ�Ĭ�5��>6��G�r��PvNL�R��m�����K�B����d1=W4'e*�&!��豆��x�:}~חRC�W�����#�p+4Eo�q�@��&B��*��P�g�s��+(��T�E���E��x�\��|�,`�o���+t�$�@Z.�* E���\��-C؃Phn�
}��w�SZ>��Rz�X޲�I�H˦�>'	�Nb��f�t�*>j�� Ч
�L>)~V�*uuR1�%��n �]���v�)����)j$���������T�Sۖ�_:�]�M�՟��䑟 ,7��ˬ{���R�;��4����Ƴ�0kh�Ϲ��z�{���A��Y��.=��藦�ˊdu�P�PT�no@'pȍ�֕&0B2:g���- �lj���<�V���%5�AYY~�ӌ�>���,����%�9�7L�C�O��c%�CÅ;+���N�e(ȋ{a�&�^�������@��4 ��F��rHu.qI���׳e�+�,�F���ey�l_
����?���$�K�kL+2�FrǺ6�l��?��
4eO ��G�F�5�Q�/����޾�"KXfeD���.O��<�U,�0�o�ۙ8WHE������Nަ�jU��?������=��s
���c��애7�{E��`E�3fU���DTh,��K
��-�_Bw���o�{δE��wi����V����3h�,���{;䡅�7M�#����B�~݌���y�����"]�����w��-�������_YF�g�5�Y��mq�X�އӾء��V�>����,Ҙ8G����~���L�<d�BCD��F5�Z�`G�n3ނ�ᐲȋ`��3�,F�
?��UB�jF�1�c\��� �2�~hۼ��2��ј�#jw�!����O�$�/c	ŭ����e�}T?�	���f��u,6=xq����v�5A�0��C�cV씕���yŨ^P��P��~���w�!=��X;�E������$�y�J�=ܞ���k�)p�Bc
�P\`F��%����!�I�vF��˔�H�.G�����4�}=W��&a>s�I�0x/A��m�����#{T��Yv.�Z���N����Pn�<���R�����I�gz��9$,b����ØI�v�.aX��7_-ZN~D�$�g�e�>r�D	+�J�u�@�+�����[\�	ﰓ+�@S��j{E Z��γu�����g$� c�3�1�!�Qm�G6I2��]jH�H&��ӣcx���#0D|R
'��[�F
@DtI��&F�紧�\�lo1��T�Ԅ
�_��kg֯��x�S��]Udd1�y�r@�L����_��~���V�FU�̕>�Q˖߈�I~��I#"�e3�$W˯2>psBI❔�RZ<d� ؜~�{gMϠ�7�_��5vpr�$������m��m�0�S	�2�����`�WJ������{[�Hu}S�����$uxt,�pV�Wb!�7�zn/*�+�#���D[K�y�@�~JG#]y���� �B��?�ad�����:��!#n����%����_T��/�_Ј��ֿ��lӖ?%��/א��m�]1��F�Ȩ��)���P���D�S��nVi|+��0��64�*��Je�7W�����Z B�����w��o�;���-�� 9P�΄� �:�Gߕ&�;�eG(ag�m�:���1|E�ía��g��9,�����t�*\z&��fh�0��2�9��9�ub�Gk�An#z�����!jUv�o#z5��s{iy���Mo���2o�O�2�r���W+w#Q��U�U���:��#6��ꅷ��4,V���}NU���P��Nfr}4���MR������&�Z������` g���'�\#s�h}^�����PS]�xQ`B0�<�?�6B{�ݫ�CUQ�9���;��>��6���Li}����i��.A�W[��cӷT��TҟH�]}�Xy����uGa)(N��͠����㴴Uz�i�$ ��%Rt*�9��gt�3��S\ �T����9o��L�M�p�W<�׻�ګj6��	��qL�<uC�*�*�mӟ������z�szSn����M���)>��-Ė\�N�I��	�@<T{鞄���^�r;����Ii��w����ؒ6��s�g8{y��C) RD�S�hw:4��ۗe�w�������
n����cw�@���88��a����)(M?���c7%w����@	A������{�D-^X�n�4�,����>�{B�(���Z����u��\�Ѳ��e�1Ԏa^u�7*;yC���ʸ۽BHv��GpK��ֵ���L���7�$i/��{��Z�S8q�X���d�kKW�Y݃�s��}:A
���YQ25xY�=#��0�%����A�����ǻ{�rt�Y+A���yy=}�!�����$��|�]�Giq��؜���g"T)J;݅���d���%��(���Oa�e	QF�ZBe���I.LZB��A��r��meY�i��z�2�ӥ��.d0H���7��j	!��F��!%�t�Ѩ��o���7vM��S"��}��Q��t��_����$��"޾{�_J�R�**�o�,�9�^���I|N�P�@�P%����d��b ./�39Q�j��U�nv��o�C�Ύ��J*U�F�����:�79��J?����6)�4���~/�0Υ��ȈJ������z2���:����`n����^G�p���[V��"�א~ú��iJ3d019��@�<2��F<��x��Y9P���ej�)����X�r�1���[w��e��{+kz��<�h9�PM����<ó$L۶C3/�{�3D͠��I�>Ow�K�e '�5j�{08ш>���<d-N_4�����+�'��`�TR���lȡ`�j�´��|Hp�o���S��5�-27>.o2�#Ƨ3T��P����@�s�ɶٮ��d��]�P�<�zy[�.z�w�s!d�1;G����O�ۀ7���e�5��7hW�uA2�ѽ�����z�K�y�nǠ���*��F�\N������q�ٱ�k���x'��wcR`�����*�/P��
�-�w�9��PN�.!���CG���&=��\\ϘsH�2`�x+�E5i��L��A ��k��������i%cW��St������z`64��_��d�*�T�uDXX�}��j]^ 5�	d>��ȁ�C�,�a�8�V���9����?�$� g��$�F�fEσ)@fz~��1�L	�� 21�0�T��_}!a�
�;�� �����WdiX�$uPm���);f�3��rt�ɷ%BP�fXq�7�ίm���P����+M,�)s��sp��W&C۴��o�	��~ċ�&�o�']�k��'���ME�����Y����m��㘖+(W��-�����8^�+����N�&�	��F�#ʾ�t"Yz���:��S)�v����&o�]�8A����ҋ�ƴ��a���LlcU� �0��&�5ֲ��F���m4��8�����KO�������!/���3�Y�q�0��*���w8=�%X/���v��)��՜>L^A���-p���褪��m2�j�y\q��,�����QBCf0�����a�d�DŌ~񯧦]O��� L�:�|k!���&��m\�S2E�y.�{��<����z�շ2~��g�k��b��*Ӝj�
u�#e�6�{���g��i�+�V�7�1 0�C�{\I����3���湬< �Yu8���>P���9�o���H�4���k������g��v�}�ȿ���EJ�S������fN\"|�-�$e�Ǜl>&,��D��Yk��5��p���-�ay�4ɗ�B�X�h
�� Q������b>�B -LzZI�j��1�3�1WW|W�^��w�L�#�
��|����5��~@9�u�x�c\6w��7�0&z��;;���Às�� �a��Ȑ<X�o)�q�D��ʚa�cU�PY����Jo,$ً��G��u}E)j:ҥ�I<�+�X��:ͷR�WX�H�W��� ���,l<���h2M�	�H�0P��u%�G�=��t�Ө�l�a	�Af�;v���LD�uX+���P����Q�(�W�@S�hCB�p�3f}rN7t�}.��0�ٌ��&�Ѽ���W����K�_���J�R�IVZ�x׳U^e�*��&	��4�?v�B�ЬJu��8_�c21n��B�X^߸�aǈ��oa�q�b��y-�2ZY�tۻ�`i����|�P]����t\n�W�ɜ:�%A�a��tfZ�E4�s�.'�dE��Q�l:	���f��Pѱ,��o~d���I�e��>r7��12��Y��qhX�́�@W��~������?7��J�M"﹘!�nAٗ�߮h�<�����!����j���*]�R7J�_1>\Bvbt�ls�F��d�	��L���I�����/��cd1h����n$ZAÌy�r��7�[��&����Ñv?ь���]z����Y C���+B������6xz�M�f�_�V���!��|����t�Ά��ܣV�IR#�dK��#G��bA���At���Ƒ<,K��'��No�oA����$�b.U����~�Ѿe!SK�#$g�1���sΕk�>��h���Au�W�����-Y٥g�L��V�PT-�"�J�W�Ҕ�T�����׎���U�M2b`��<��bu�g�{ ����M���5�>��Lr�eo�Q���"R��V����j,�a�q��9��."˔�`*l����X�^X��?l���3�{����A�r�i���Ӕ:=��=e��,ѐM�vM����&��F#���	��4�O���uh�Ngz����C���ZY�F��{o�\�&��d�]mS@�4�:�B�\��V���L5k*9t���I
,d���-���k6�Eu�j̪2r�1M���,�'D}F��5!;�W߶Ⱥu���~Yz ;��D�N�,�t|���Ld�Gݕ��̕�R��óe<O�V4�[ʀa\j�`zh��J��x���,=隭(���4Z���A��~�0릌�1�D�����)^Ժ��{��)�]�S�v���V�9$��s�������^�8|�O#�6���>�~ɷq�?�M��Ŏ��?��]c��K�~+9s��o���-|;�+���ٍ�q�������Hɮ٦��$o�|�uY�%�M�n�,ň��,#�V�Q�<���Α�����.9*���r�0MSqVi��U-m]�B� tg��=_~0V�U��
Z�;�R�l�Ɛu���ǻ|�q�A���|0�R"X����=�� w	�V?-�x�+�/�@���[<΢� ː���d���S���dp,l%��(����7s%�����Q�X���ZNzਜ਼�Ùd�e��o�)0�$�j�e���2{Nζ�x�\�����l�K��,�B���SM�C~q(�dg���c�\�Ϡ4xq[d�;5ڲY�ѹ�~��e<Ѭ��ƨ�$|���-��F\m�3����H���TP�/.h���� ���?6!T�T/z:��r�4<���r���N�L���'�U�e�e�%����f�`��u�����!�\`<�]��?S�C�Z�R6O敨�J�1����76 _�Ϳ�~�ek!�Y7H�!�r�L0�F٤��3�h�n��R)r���5"�I�~�M�+����V��Z�;	Đ�3
"���q�À)FW�A���n[K�e̩�\�Y�\'�;d+ˍ��L�=
�/��kP�����9����\F�Ë�����T�(�J�ɇJR�E�C;z�ܩ��r�be0dFݩ���5o>;�1������ni��K��
Ϣ�r¦�F��̴Z�����GE~[�(,zE5rES��.�+>�t�T|�]��P)�r2��N��B�8l#w�_�h!�H�d'Y������O�<������F�%>���f&(d?��*���T�rכ��ɜA���av�����U	)=x%f�@_)ru�)�>�?ĳhk�V��2޵��,�4x�kۦ�#�dT�N��`��+��#�3���:�Hh�<%���9��2c�W�Tlw?̣��j	�U�,��|:w��7֨AO�ne�'����:�|�L?�mL3�؀�D���^$�k]�G�	f�&�L�߅���OAf�P!VV����G
��D�(֚�	��<����P;�{�h.-�dI�F����\ٺB_�ƤW�(�Y��X��4�9�ߚ�@�ٞfo�ڄ�1+�(�櫞�z�Z���5�)R�L�����rz��� ����#���8oB{Ӛ�A4�����%{��8���e��8��L��g�q��>Y�q��:R-��_D�WER�R��\�ׯ�Jv"R�P����M�n�ֹA=M����4{6��mf,�iuI�N#��V�+<"4��1�L͟ؤ���T����DGY�6�����m#?fY�}M��%`6�ri�\�LH�y�R��`5a��*��`x�T�es%?%�Dn���T��p�3� �b$�ش�$��tL�_�ͩ!H�����\�r�}��i@O�=G뻿�W����J�r޳�&,�з�F6��������4��+�dP�L�^o���I�3JeH�r�W		n�6ƾ�[<�o>��V�b������_�JɵC��Vl�����r�D�:d����{����Ow�"��œ�u����TT����*�@��*�r������:��E��'����o���6�w.򹬁"h$~��¥TG���������g3�/�{9�;�!/�0:��`�΢;(;��L��93X%�<j�6cQ���!H5Qu�������M�6�{6�-�u��J,��8�\�8���t�~�:���axG�Ј�N��I�̪ ����P%��i`�q�v] d�}̔�]�:�Bʲ� ~[�b���:��x�^Ʀ��I��/-�m1�����Y�4�b�s�����Сʻ��[4ZN� �p�8-�V"#V�A���l��.2�tpfk,�"$`�Y7�6C��Ǐu��V���y��"M��K�Y/�a����e�e*�1@H�hf���$�@?�%��*���N
n!=T��oV/��z���������y2e��/�~�97���B+m���U����"�k�hAd�l�����\ ���a&&0}R�W������ş�B-�^XJ��%k�ޘun�wy�R�y�,?����T�wz3ug�f�'�>����\��Mz�V�ptR ��x4�X9����m�I������^}�b������q�,/Ri*��ˁ�Q��w`S`�o2�q@c��KS޳���Q?��E���&���~�:ڗ�g,3V^8I��Z�`�JT/,���.��'��w�� �x�/�]|�ŗ<�7�NIG���D�٭��򘅬u��&nc��.4?!�L�#3o����~Z94#�����馷���@��-������#�>�Q�ƞ�iڇ�n-��Z|$���J7Gx��`�i%m,m��{o+㑲��G&�sf�oR<��?��=��q���8�j�Ͼ�)~�&��Ň?�=�LṂ�V��U�Cy�d���[�s�e�9�Ё ���o�?��g7�)�r�kO}�B�9�0���w�HT\Q+���^�$��n�W�3�Cz��������Bү���	�Q�$TRQ8Q�c��#A,��!`��������*a�&�|��
G�� c�1/]>����V��[�屳W��A���?�������Jz5��@�f��p��\�5vd*:�;G���T֪ka:�S�[K-�+�i�Ky����D�]�D��\S�����p�5	��Y�%��X�2K�l��M�nv�~��k�z$��8r������7c*A��5�ޚ�.�*U����甅��Y��s$�����F�q�z��d��T9#F�s�=���ٺi��w'`�9~�<����L�B0��u�3?*'pzp2q!�
mӀ9=u,d5��8e��r����th��:��&'ɝ?�c͗yv��E�O)���E2�CE���ϝSlo�<��ꬨWO�q��0<���2�X��<�	3� 	�(��;1"��I\ZR�:J�u��pؖ��uV}�}����0�1��epGote<</}OL�w��m���C]����Y�o���w�I�7,�b/^�S�K4��o1�,_�x�R�/��g]̐���A;�c-\o� Aq�^
x��Nַ���u/����]D���12-����Ѻ�����N*� 2�B�w�mضu��[�C'(8s��]F	�Uo�˃b��v_�����J��7�y�AnvӦ(�N�W�|Ӟ㎐z��[���M�����J�Z� c�?
W�Q�%�q�|��4��L��T{h�kI n�hn�c(���{*����'����]��Q����Lc��'�5�
y�s4�=wv6v��sB�?�~_+$���e0�H1뱯<�;z���@��j��[�D�s�$�O�vuvK�q�wi=x��X����~��l��&	(m�	9ndI�5��^b��M�[M�EC������{]�����}c� �3J�*C��s1s11c#e\���S~��igq�O���ƌ�{7W���͗��tu�Hc=��E�C�G��`$�Wܾ[&�Y�V��k�;�o��Y�b�=�|ژi_|�`! ���g�ip��>�2��u:��M��㸣���o<&�Ę�	�%��P^��R^?�Xj�M���Ic�:��o�7���i$��H��$��n뢸B!��P*����η���@y"ZJ�d�v��N}�Mf��M��R��w�z�Y9LY�p��G�.�$�AL`a��M�y#�k����M:?�R�;�����o���&y��z#2�	`V�a�h5@I-f��Cl��-�|4�(���JO8.�Tiǥ�����}��h��k���45��oƸڱ�&5dd��Ѫ�o���5�.�c'�5�A`>���3A�A�k(�u֪�����"�m�^�Ò�񮙛���;]6�J �p��ұ����ӽ��fW����y��[�Ġ�.�ŷA~�t�ܛ'D��y(��N�/r��L���I�E�S
���G�q���b*MP��6��^���Ȑ�h�k�$�w���\�*�d�Z�ާL��:�;߆T[ğ�Km�q�R��0�{��*6k*v�S����giԐ�w#.�ؽ��h��ߴY3�/�z$�V��k��B�����vr���4f�Ju=�'8i� ��~�����9�	���p�ܳz�������?+������>���ГnN��<������=�����M5�ZǩQ��� Qۉ��;���۔Y���i���3So�Q����A�f�b��M���]0)�
j�Rw��o ����+n��}Z���6٪h&/
����I�8���;�Q�{#v@�ͷQΖ��$'��]bu����D�J�S^�^��_�(���tB������R&]$4���
��'	fZ��.��{@L�btU�	��R$k�t�+��'��T��gn�� A,1����OP8'��`�F�"������� Q�%f]�`V-���s���r����н/Ŧ�98'�>��HWo@4W@���{��D�!ԯ6�}�������t�?2�r]I�|����*J$y�«!)��r�ɞ�c����A�CO�պ&Uȶ��#>�s�;c����z)M���36��,��ԭ�h�"ߋ�Ùb��Z�I?�k������6��UU|Q$�EF����4!��\�AbU��`��6�� �h�|*��w(���yJI\����r�@E���V]9�@$��A�U����A6��X��m�t�$v͆�{~,4�$(����۰�`� ��ZY��v#���ȯ/��Rٰa@h�Q���v1hh3?�r
�~�.))R2K3�⫉0�{<��嫈��6/�E�>���
�ɂ�T6�?k_)���r���Db���>���ۑ��3L	B�\"��δ����ؠ�-hN�G�� /d1���l�N���j�Q;h��h�ä�xf�a/T�X�ƋT�3��\G������g�$��ȶ7����!�0��?�^�� J�=��;�H&�}]�6�|��@��OC[�Ԇ��>n���9���)���k���~�"��{�_{��,�E A��!�O�ֆČ;%�ܟ�44���m�s�]���Y��&P7����ʹ|��4�Z�'�D9��P���(:+I�� �Ol����RÊꍦM(��؈� `�Zw��S��
�����F��)ڳ���	���,�Ӄ�����؎�a;e�>�{��@�]ap���t$��D�\����45�o軶H~�1��"�CZH��b?��w��R_f�_��+�"�'�$�C��ݾ�^Y��qr�o#AF��K�Hy��QZ-C|�c�^�������.��D�_�������gu	0B�;�;��Kג��" ��(Tj^	�>�}��7(]�l�B�zʛ릣ۦ[�b1L9��o|QGI����k�����ri�R,����Zll�^O-
�v�4��n�����^�At���u�Y8�j-0R���[~�nc�C����|,փ�V��gSk�)�����г^]��~�!�g�ڇs�(��/�1�L`u����iK��^ �Q=
�fm�Q6��k�۴�ӂ��"�qu�7?z��f�|�� ���/;��.$U��ݴ0#���?����"�C2.���U���_2)���%��� �]3�o��Nbq��0A���$�Г鰜#�B�m"���A�b�>^��ѱ�]ym��6�����Z���f�弞�.�>����Hi*Nt��]�O��O�F8_,O6�+W�'D�ǀu"4�b�<��L�a�cPd��~g1��Rŕ�Ƈ1��ƴ����)t�!xi	�M�LD���R�`j�����׎���.6=�;��U�5��Po��nl���a�lM]�έM?�� i:�S�N?U���r�La�.����q}��]�K �E��g/%�V��U�O��h�͠8}���h�	2w���1�Ā4 �j#�G)w�#��P�F����G>2,�tFɵ��kf�n��^����ɗ2j�]��؍�[�a���[�O<�_���5��F쾣T���}�1�������zmA��\*�7��
�i����J����s��'e1\(��=��[�-X)���*׊Q2	�%�3+F��R��j�`4���l���10sw&i��"�yȾe�8��G�%���Q���l�m?q�@H؈A���!�/��ޛ�ῃ�kGb��R��r���P+�ғ@,?!cF��m|pǨ�T17&����!����XG�Bn��)�JWn�!v�I#�, ���#{��6߇*m����3�vƗ��!:�p�P��y����͝v�����v+�
�C�o6����2���F�"fЈ�/T<�9�kY�~�u0D�����`�9 6"+no�vj��(MC�} f��4}T���ԤK�4�;�~����cn�id�s���iu#��1�0_��)xڰ+�ۈ��O(DJ�*:n�=�p����~�j �P^f^ ���*?&PY�����Z�ɦ��R�	W���Xރ�}4"P�`9�X݃q�Z�9�:d{��RXY	��Oj�n�%����P���A�R���>���whG��Ŗ*%�����w|yM_& �)�[D�c?e�C�Dn����O�}aPr��9Z��Ҁ�p�,���&�`�K�&�VeU��B_ä�2�C3<Y_���5�j���3-ː�z�ajj����`���0^�أ����?K�j���]S��	����!繋����A3��E�@�=p�O����8wT
��;�w�=kH�3�e)C�g(�s��c��G�������Bm�M��hN7ky�*T���5���/�*�p�V K��OG�(Q湟���9ZK�%d0?J��U�����#�h� �$�j��x��Kf!Co�1�6��ș��5�~�⥘��׭�uK��+���<<�\���!�ՐӶ���DǮ2�\o�U�+�p�`?�Oȸt
�c0[j���������{�_�kƝ��ʒp��I��r@W��Xuɍd&�h�i�����]��H8b�v�R�$g�u�����V��-�KNJ�:^��Ƚ�`��|�W~�3#��,��������G-:7��F}y�ЃYJ?]����T�����u�N8!X���(�Gٖ	K�ܕ��2Rw��k!���d���ӓ�Gf�%��G�}zR�-���k�"�;>�����x0����F5"�jH��G�åp��T�;�����%��2�Ч��E$��G�7a}���5o3�n�zrQpJo�=%]0O(�у1"6t�W��u����%R�ܙ��D���-+oz�j���Szx2\����|G%Kє�i�A�
� �*4p��N�]�q
=`���e�VMr�&�ԫr�|x���G$ߤA@;�<_h�I~E��mRrf5�!z@���E��Ĺ=���t!\��*0i�C�����@�"���/�?��KOځH_�ZvF�*���{��z�Et�/][%�������B�R�5"�m܍!�� �;�Ruս�4���f8�4<"v�κЃ����d�C`�(:2>@��:�	�F��fC�y��c�#��[�|s��2�[f�jq�{-����tqofN��Ae�K΀�,$�;d���W���N]e�f��B8�r]k���tA�u�7x�"�T��hQX��U�&�)m����!]�SnF���}���A4�r,>��#G�/tH̨Ohf��n�a��:H�8�U��rK�.@��8��}Z���x/�h$��x���)#�ebs�#�i���PK��`�
�@�b�;�}
"��ӣ�>2|mP�U8��Ry�HkBPx�'	K歏�MG"���&j;n�q/�yr<��:��{өy9y�X6�c���(B�g���T1�ώ���FS]
]��8�x�{7�dM�{�q".����a^��
�2����ByL'����$_�����GŞ(�K�M�et�yt�E�8$�2L��%X�Q��,���ƅ~8Q���r"�K��jQ�T�&�2ܓ���I�ϩ���n���#3x���ӎF��+��M����y�pl$��V���J]�������p�IgȖE�C-_�% ��}g-*��k m;�Ǭ��6qa>$S	��`���4���~6��s1E pЩ��� �p�%P��׬�I
!\u �\�4�H5��d�b� �B�5�>?ctwMT�F_ԧ8�o,q�48t�
��#&b8}�p�3]�M��L�G��<�P��At����D \��L�|�F�to�PI�q���?�I� H��X�.M��q|�usXY�=	���ԥ�@'<���@��V-z3�=S_�}NB%
�'N7w~�SF�[99�$�S�����b�絯 ^�k,փ�s�}Y͕Z־)8��+̺�2ʇqqlC�r�Z��j��ް��"M��=HxB"�\�H+64L��W%�}ߊl�����8RDS�V �jg��{2�ѭ�b(Z������_�5Z���sճ�~AR	���L<��t[�x��I5�r�#%6�w28m�^�&�x��!M|.�P�!��㖠�)�YE��69��em������&�8w�R	� �IpC�0ҍ��?"s����WH\���Fh��4����Rsq�#q�B��+O��v��BI�S츫�YG�)�m[��	�Rvq�~(���lH��\�#5`�/s�/5�ҽ��n���.{�~Ң1F�yjz��K�M���V�ԇ�Zf��G�Ő��* M�&��p�R���S(��x� ��|^�\���W-���&�V��]���_@`�w!����6�T<�Q�Om겖 ��*K&�� ���`ԀO���p
�s�zod��u��ޢ���3���B�q0��x�'�22A�Bq��zH�L�k��=D�R��D��ڑ�1�+I���R�?��݆Q���-B�;��y�x�V�����ޏ`{���bԸ�C3� ?�_��<��D�<oΥ�0/*:� UPE�k;j�)��9� ��x�S;��F���a�Zi~�aԈ1�b���QC2�(Rb����Mx�#^R����C�|:��g�F�#�q_-P����v|"nT�wVOX��|�t{	��������H]0m��E2��%>A�R���->�=l90ZL��r�j>�T�Hb�mZQ�u �'�Yd�5�Q��uB��$����oik+������f�6��E�c��o։dTZ@�~�m8Nq=�v�9���	��Qd��o֞F��b;x$��ޢP��}�&���e���K�`cl~۝��m�c��c��MZD�A��bF{/vg	R���V	��ۧ�ɧJ��[tIk�\��+���t�5�x��Q���QT�+,�+�-�UȰ5A؇�Aa}�Ĕbv��Ŗ�P+T�r�;>�
�O�Y�U�^�)�?�N,�\xm8|^�ln�HQ������}�/�gYȠ��U)��P�L0�9��$`�,�CFb5x��J��DCoRNMy�޶��ǘ��U��ܚ���3%)V"<PM2�5�㉎�����*n6
G�y�k,�!�\�_x3ʪ����BO�&X#�#�L4���dT�����e�ް4�|�{du�}~dB�.D٨��-�O�f�Uu�k�S�K���*�� v�~�gm�~q���7~���"�Y�_�M�#`f�ҽ'�Vs�
?"�@�X���۰jXS��'�$ @��'�G����v�g��⤹K�&�`-bط�Ip�`3ě��S��j�A�>���"�E������(=>���D����"��%W��ȡ�2	�&��h�(y�|(��aG��m��p�1��_�Y�O�����@B�C�\��{�q��i�H�ng��D������U�������3�+�NkC��,�f����<��'"�B��*�rl2�j<���(ƩS�-AՁ �[�<a8K�����i�4UC+�[��_S~��i���=I��<P���^�>��ے}C1v���Qe"i�񰤹��2��|p��:�ۻ`�A�:�d��y%���
���̶6�?c-8'�(~-�L;F'���P�u���H�]i���#;�s#֨�5A����yב�H)��V�����st^/%����l�0{�l'~,�q��ݍ����ww y~s�~�\�3�M��Ed��6)��'��"�d�Su�3�s���>�aܹ�m���w���*��~Ԍ�B��Yr������9]W[E�'bA�ޡ�u:��z��Ag_��ķE|@?S��{S.?��c8uC��	��������#�0yՎS_��TV�),&�)�'���j{i��¡j�6����=׿N&��t��و�= <�X����F���M��U�F?{[
�X�%!%�O�_�}>�^5Y�8��{�L�PFք���D��~��y�X'�a&�C 8�7q�]q��A�8A	������%s��q��W���3$ �*�S(���h�@(�P�TB7
��?1�<��*��@���xtʹ��+���t�I��5�0�y�Q�`�*"���X�gdV��=fE�v?5�[���7N�*�=���)j�mb�y�<�m��0l< ��c��R�Ռ�p�4��t]ҪG�l��h
�B���׻shp�~tni\'�����>��U��'%Q��;���F:Ϋl-.��į�-'.�=}���t�Q&��RCth1� ���;&t-�-������3^����U�����1����7�'�95,4�����Q�n9��w�pW9��`��qI�w�6 �R?�k��ė9�ⲅ���H�|S88P��b��|1��3.��1YD�0!�<q��|�DA�u�c��"\���E�P�K|�E����3�
ҍ^F��C�����$�F&B�i	����wnhDM!HC={s�ͰD�UA�(�?Ғ� r���U�)Xhݔ(��U��*�ļ��u��L�#(p��j�9��j�q�o��� �T�8[S�X�C�R1��8Ɲɑ�8��Lhw���$4�j��mO�jY#�����K+y6%|x�렯S9�4W,W�%����2Z>���Q۾哀}0zH*�b����w�_�!�՗�?���g��AhJ�n�1P�o)y�9G�S �+��=43�`���D��g��b��sws�@YR��`x��ld/k�y�I
[P�vW`�DD�r��ؙ'j7)>�	�޼��ܔ��f�ǁ����1�g��iA�(��[��@��p����H=0�1�%mGYf�wR���&1}k{A[����U�!R3��<,�R|���^C9��t��N=Fxf5JؗY��Z�R3h�&�SuM��Z�V�&�F�0���~�ۀ�6��5��W��,?� I{N._yF܇r��ޙ4�]Q� o�)���D�=��{�RCn)���{��gY��㥹9�mn�S!�Rb��K�d��#!���K�$�%'�M���]c{|���sy)�Lʦ�c�u$�l�h"w�E��j,�~!	%�@	]-�2�������M�՝q;��pRg����Y���a�Y��D>��H�V=e+���B8	k��i�z@���I��;�)�U�����Rŷ�maXM��wF�֏Шz���}A��]�a=�hhw9�����Reζ������Ӻ{����d�2 �ؗ���7�ʸ#Խ�k.��o
*r>`A�9�u�߄\?f��7/�t�4�X�j&�ڂY ƜĲ�[@@��KK�}1��s�,���]��β[�Sv�h㡰���Z���0�ȃ}��?,*�w�u.�P����
I�G�=t��[���@`�j��:]g��DZ�a,w�A��yq�j�o͜g����5,u�8yfM&��vx��"/�\gK� $��ś>D�����n���Kd #�k�zL_������h��"�h.���d��`�lw3�3ޚ@�"|���p�/�,��j�6�����Q�n?��iL�<�L�h�����(O�{ե���.���N`1K����@<��VWD�5Ũ��$���Br�"�+�p�E�(:��%N� 8�79�$�,F��B	�����l��?�l,�h�n��R����o|gļ@U���ȁ#�ȥ��������
ddJo'(�EB��ST���N�[�sD�H`�>1��q��V��!@����Y��Ǫ����@�p{��>'@r��A�X2�n�g"�GD��޽"N�o�g*e����׶Ho��+�9� ^h�����O��ޝ��<�r������%Y�xxM�&K��>����5$��G�Q!�aF�A����<��u��x��]�O�/��$�jE�H����m,,t��������0T�a��exH���$a���]y�	���SF+�q*�%����􅎸�9����Xmg�/`:j���My=tZ����PH��<%�<��%�xe!&��g�ߺ�:�}t�L��>H��oi��0�K�"|#	�;Ψ^%e�-�;��	ׅ>����� J�eu�z?Q��	�'E���j�\<ggY��g"'֢�A%�w������)mZ���UwO�A6QH}�J�()��3N��:\6A��G�>��*�v�b*����Vd�.����7��h��fk!8�>]/O<b4����:ǷfhY�9r7hoĂC�>`"Y%�/���S���S�n����0���3B�B��7U�zc_�C�����x�&[y	ݘh�U���?F���0=7�]�hk2����T��c�͌8��8Q'6 Dv�Q�sS�>p����) ���,>��e{G�̐$�pK(�%=ʘ=�7�S�@S��>��̠{�JL��q
0��.U����Y���O?i���e6�f��CX�D���\	���Rg�Io����ʜ�2?�6���������,�h�5�;�C��,�|�ۑ�a�6��q�K�J�u���Qأ<���'3�����6\�&J&�h�v>�ީ\q`A�4���������`�tރIq��YG�QEA#僥00z<��>?�@�Ev���8y/Z�Dਚ1��3�b� �b��&��*�ݝ4�]L���IY�Y����W�Wk�$����C��3��Rx�Y]_���}��3��1z�Q 1仔�J���zs�(�htDT�[�&Vh����u�u,I4e������?�&x�� >m��b�L�5�[޺�E��K��	ÿ����ޡ/�3<��3�Ȼh�C�W�Π�
��l��ná�q"�YMt���z�H,|�"uː�;a3/p~���QSM�F�d���D�x��v�[���b��C3��c���vU`�2�\�s�g#;�Z^!���7��{8�x�{ �H6����V�Ҩ㤟�ܞE��ɡb]�vjƎ��.�/��ε��^8@���w���M��ݷ��`*@�cb�&�V������$�����%}����fh�MPis�X�n�&� ن�lX9��By�d41JzI�1v0��k��wų�'�
�Qb8�t���8\�#�e�z6:��aLh:0eY5�&�@x�b��5>������#���lx�r_}]řN7f��tT*C4ǈ7�ZGΫ�˻6�/��y����&;hcP{L�vx�V���4l12qR��`9y39ϡ�jK<⹯Sdsv����^
�C��_���_I���h�F������0�1=þ�6�F_C+V�	��N�k|����C19�B�lی7�Zm��kqz��'��ǭ+�;x����T��7bæ�. �EGi�]N�Ȁ��IĔ��"��co\�z���țe��KP!�D�:����%v������cS�h�|�k�_�����w���LN����g��6��[��?ڻǚ�v@{J�@zU�6d%�!y�F�
�Ef���A��K13�Uq`��g�<u���Ů��^s�֠	��G�_��m���X��3=0],=�,-3R��xg�g�l�hu��IT0���Tg��~Y��k+�)�	oR��\1�b>4��Ϯ�� ~`S)sns`WP�R��y,H3g}���Ǎ���i��[\���rT�a�!����O�-�l#���Yhq��E����mC�z������e����1-�$�IHr>����A�:�`J�|�G!-��c.��ʟSU˲6��Í�QW؊-$�v'�}�1Xw0.�7}�#Kk�2
�/��q�C�h E3/XR�ۣn�y���=���Aױ�J;�eO�_�\8�%d
L��O���r�������z}S;6n��}�񊍆��C�a$2���N����$�AIa��X��k��̨/���n�/��N�Tx5��)��*#*�V����ῡ(��ۓ�/Dn�M��]�`�� ���\�^��3��j���_�E|#୾��=�ص�b�'W�� 9I����[�"m^N<e�һc�`��yjo_@��L�?��~Y�$�XKJRtn����u�hMU��/S�˟)M^
}M�N"~�����Y͐ �h�ˊ����1n׃F�m��N:���F��QlԺ2��Aө��'�y>��Ԍ�usMH�q�����7Y�� )�?���ߌ
�sR�zf�e5�v�`vd"�-�8|C�R{�'��ٟH���ƓIJ����m&σ�X@R��Sdt����c�snہ�z]�zDb����k��U����!��&���l�<�c
�&j�B�W�|Z�}��ҙpi�*�y��C/;r��⯋�s��hT���_�������5�{�ﰂ�眶��@�z�L���XZ�sb��@�&��Xd���x|:�QK�#��4���G��O�k�9�����5�h�x;��c�Ln�m�e�j��wĥ��uu,�T.���m
�*�M��*m��l(C�v�	�]1G�@�
Dɾ��3r+5�=�����a�G9��X�v����;*��_���CO��~�G��H����S��D+��Ø[jV��/.��9>�:zdw�w�+���s4�n���Yy(�܅�g�:ﭛ�;��Y&�-Y������ŷIHM�bơ�lE`m,�/R@9_���jK��e���o��(8P�.e����(ǆ%�n4={�{L���y��'֍x2J-*�QO����sU��'�0��1^��3@[�h��g�; j�2:S�PX��v�"bp�z��?��C��!���#���m�d��ˋ��cyY'�^��.�X�w�ר�<.҉[�ы`�n|�f�AEL�o�$<��ڈ��0��O�#݁�.An��U��IU\��ަO��;R�z;^m���#�]1�(td��~���k��,l"����A˖�S`S()7��g=�Bw�����`����~�����#�\���M����&����@�R����T��#Su�	�����FYV?*5��U-辰���\B	�+ X��Ӷ����j~�n�da���U���1��U#�6�}HS��·��'�Nt��ب��Ȼ��@g]��t*��X��	R�f!Z�i�:��>��S�[ᄮ,DL�j3�I��ۯ��l�Q��z\M�y���Nj��N�;L��D4W"ni��X>��V��;�ˑ�
^�VT���'����j�+k߻hq�s�(Q{��P����	>������N$SW	�^����n��U��cRgb��wt2vk��z�s5�#����`���҆���4�Q��1-.b��3��V��]�=)׸�Ϳ�<̅*T�����p�� �M-��l���r��|��<�7i�2͔�F�'��Ea��Ui��Ό*,/�䞶���v�g�ȘפO]9�荢���O��υC@W�65�J�Fs�-�#�ŷ=��p�hf_f�ș�v�xp�!j�����J�V}S�:���H�lʹ��ϕ�2�]��8��c�p��-߲���/3���C���ج٘��.4�Z!��CgFc����)�Q?(�qS� �z�P{]�[9����\I�����=|u��_�~��������yxMq�����SԘZZ�Z��F���zHW�N�z�0&�H��I̛v�]8����u+.���(�N�B�6������l��&��S�d�� }�r�Yg8�]PW.�R
X���T^�r/�yF�m���N���[@c��gL2ͿT]��M���d�ڮ5����R�ʆS��壑�
G�9�[ㅺiw�$���G>+n2z���csr{�s�Bs{�W1��u�}�t��{��&��{JU[.X�޺'���SL�4�E<�uS��&fz܍pik�֦��>j뗗���vf�x|e#����}�/�z�O��]��V�=�_����}⿌`�]jv��݁$h�I#%*�0u���w�������#1����vk�gu��r��.�a�2i��c��:���h�ʤ#�pGJo�p�`=�((эh�������;��&g�c��.��[$ҳ�8�z9g�1��?���������� O:������s�����H4����f��p͎�E�5y4/�WW��~�y��첷����� ���� �v3��ú�����#��՚�4bY�Ң`5R��g#`8m���e��)Fk������:e*FRi��%g�/��"��RG��u�
����ۚyL�*�Z�j�j��+�Wop.7�{γDl�|W_�@��2�h|y��<m�՚�ZDf�⾒���r�h�W�Ei�+��)���q�D�M��D'�H�s4d F�b�W���*��q2V���6)`�CdJ�Z~��%��v� �� ��/$M��~vT�w̷X���eW�Bw�k�-��̟���44��S. 2�~�]�0b���,�~�ɗ��bcm:&]V��P��a��1#�O���A�E�U��ƿ�<�彊�>7O۬��3jEX���>��Y�^7xA��*�ĥ�;���[��:����HO���������7���o`�ꀓ�����?��rH��Uj���N��?L�
��oK�L��ĉ�A��n�"�(Z�i��h�fG��� �X�8�k�Y x�r;E���p%W�Ք�%Ȁ+�>�s��'b�y��h���!ݠ��U7�V�6$���gٞF��X@PV�md�0B �I�r	��L�����V䝶M�;��xI���/۪WI@���S+��;��(թ���3eKz�.�'����[.�f	�r�s;��~�#�H �5��}���Q"���ADMr� ���:C���i0�]���G�]I �4Y��=Q���ʏb����rvt��y��""�7ܑs(�����g�0��� K��J';�m���螎5��vz)AsCj��	a2}�d��z_�wH�#s��,�J����ع���a�����Q�~�>�8��AC���v�>�Y;� OvX��U���o�řS����1c��o���ɢ��۪��s�A��Gc(�
TE���o
Ro�\�*���.]��N4#��3��_�%�
���xL���(W\�1~�>Y���
��߄��3r��S��qr������K��45�ѭ)�����L�`c�Ք�C��9z*z�={�'9����sB�Y�Ʈ�Pr8	���u��y��SwDZG�{A�ʢy����/P)DIP_,LN�K��p���$���&�����t׊T�ăv�x�ș���<h{��~\���2�3&�w�Q�� �#{$mE�a��R>�%R�k�<��k�8H@<��Cgv]��?��`��l־}�C�|�R��$QI6 蓏D׃A������l�T��d��?����0lK˗N���`��bB �-Z�p��I���L[�q�Y�7�$:������}5ءO�ӓ�A���<�U3ʨ���~������T�HE�`q܉�#�ZVb��M���]�4M��8N!��rݞ�j�O�[��^�=kG[�@ڡ�e���X�Tz.�ap% ����e����x�ܘ�Ur�����x��a�5ӊ��-���H�T�*�y�i�D�����`3��2m��ڎ�>���7���r���'ŕ-�P�`
��8,�`�V9w���D�""�E>.��
���⻖YݑR!�V���/�I����S�|����6�M(@3��{�І�y�S��*:X�O�Ԩ�^��B�<;my�a\^[�]hİ�"�mq���\�l���h�d�k���,u�_��F����qrxG=�~��	�ᄪ���H�����acX�Î��U���ϷC��ʙ���E���K�!rU#�$j��L-2L� \�˛�Y��0=1�Ǧ��D.aI�be��.�y��yE/���[ ��{�r�g�ʚ��6��{�i����J��a=�oJ]�}��"���)@�ez�Q��P)�}�t������ԁN�Ⰾ�J�*�j�.°�d��L�3C��PI2�����I�u�ƻ$$�*���ݱ\�
�����T�y0V-yP��N�J�G_�Ak#LO�$$X�l��P�2�`%0���R1@Cg\̺Xd�+P�8꯰�T�B9Y)����y�T�Y-n#��x��8�� �B�u��М�����m����9t��4���9��c���l��j�k�ԇ�.	�ẹ*�Z	~s��)}����f1�4()���;+�{bu���ѱ�s���F0^���0% ���I7�G�\����M�M��C7�n�4�o��-�!lDI&��Ct`�>�yB���,��=Fx�]@�@iaM�L��uR������op���[�\�0YO�d�G�enK�5k㵛�2���|�@�ܰ�2n�zܺ5J��� ^�%I��7<>.�����w�7�x8���ӳg�SJ%}rK�5�br��"j��#�r�)�)�e?&1ʵ?�H�v\8�n��T�J�����	J�����6Ri9�+��յ�#{.���p)��o]�>_�G1� �тh��#&����z � X�oz�X�������"̬�C*gcƥ���~�W��	�C(oi^���M��9�Q,mG�܅�x�s�5=��.�%��X�J�(OL�"��#H�`��>�5e���9U��
�y�������d+{Pw.MC�2�9/�<��H�� MM�=Q��I�B"�X#�[��XpyD�����i�~�����P/�5x q{�TvlW���N)9�G���Mk�����`.����~e|�j�Kt�/WP({��7�ؑY��	س'� �{жR^X��bj/
}�v���,W}�%۽�:	?���4���J������P=��68T���L%_s4!���n>�S��l�A��Y%x��e����ȹ�g�M�xsBv���\L�7\�9+�E9���n�V�0��P�������?3� �>;��s&�E�;�V�]2
[l�Y�_J��vGS���_+���E^���o�NE�<2����Aˆ)��<iY��,��a��������UD�k��n�f%�>8���-k�CaD=�����I	-H
�����,Hi��Ls�Ih�����O��W�Y���҄HUu�W������e��`#alMg���.R'&��5A��nx�6��M�1��P�ʣ�^�S��.F����Ǝ�p2�K�-�����)�����GB)�~�l�N(��V�[@r��&-�������vq6�n?V���_���_�b�'�o�R�����&���J�n����#�u��~8�aam֢]�*����+�[�Qgx=�� Iu�j֨	%���nX�~e���r?�;Y��D�r��n�L�5����ҙ�^�$U��S#��Q��j��� �S�)���:�;W�p66,&����B���Hr}T��׮���[({�vQ'6j ɳ�Q��<}f�7���x'ph	n�(�XJ���"V�f'o}]϶
�{=-��S��7���;`v9e�~|J�3g���������%�4�����G<��8��q�$����2��̑�-t��W��L��0��%cD)uԲ"'���]Ї�F�O�*
h+�%i���3��[�m��-��M�^n�B��h�dq�4��繓u�ũ�?�|LqK
��/��4�"-t�ťi��7�O���("�{p���i3nbvP�	,�)t^�!"=T����V+�(/LfXL{��^��Ht�j�)�/US�q�l4���d[�y̑ڷ}�Du��u\�2<��i9F�TO�(vM�Ay!�i��p�����[�W��t;��ǕX��+���K�l�	:�mT��
�-Tۚ��r]fon��:!R955�eK�����c�cw���q�D����Z*�Nԑ�Hq�'Q_���y��i�4�qN��I���/�(�]�4V���;�|�yQ>_g���T��b�溡���t�.�K"g�5�7S�y3�Z���>��s 6�ò�a7�﷡�L��icq�K��,d-zv��5�	���"��g��)(I�I�@K�n�B�U^�(��k�
��l�b���:M��xcA��\Y��eS��~yT��ww;Aa�7�j��ٹ(u�z��訂��3���qZy��:�x܀H����5;B��_���p�M�#.�Z���F�s�h���d���s�P?��t3��k�d�u��B���K�=���t�
a�-K�+�EFה��&tz�������G�"�߅����~p�����<�ݬ�J�Hu���?�s|E��)c
^��Xe1]�B�\1qD��QI��-[p�P��~J���l������%���7���ػvk�B���I�=�3�W!f��[���@�־�=y������[�z��슞�o���k�Kn8�?�#�p�K��	��;�K�e��A�`�8���	TͰ�R����&9fI6򉃨�m��>�H���5��B�ؿ��ٜ�g��~�s=��--����k-0B�y�P�/Rg�~�kUw��_K���g�v�J'�[R�袽gu;�q6���j|���~}�o��m듵�p��2�|�g��u&/:��gbo�����ex��P7����"1�.��#�}Tn%���T."�jW�'4������0�ě��{I��5y���!��_�1'��"a�_��Q��"�&ݑ��vi�Y����S��;$�wJ&��Y���˕x�aZ+}qpSҢvIm�m0B[�fm�Jf��/��P�]u��K��w�2�`��
�3�G�P�l���%P��>��j�k#��z�J��Ђ/���C�Pk����g׻5@�_۞ŧx	�{�Fg��ɠEsF~N�2C�X��"�7	��o��9N�ZH	�M���W�8e��^"aF�Y�,+z�,�4��cAtj��p���{�el����'e*RH�1�exPzc�aGq)\�)"���z8�" �4��Qk7���?ǚ$j���|�"�p]úy�$N���(�jWd�_�q�P�~V� �?p�R�cm�CP֖����J�������E�5�Y���_g]�v�E(�tgp0a)�����w�i���*m�TY|�@�����%��lx�xEz��+��w��d�*�\�NԼJxܞ$�I�@�}-���M���	�C���J%�Ud&���:��A�W���E�|�b)F�b�wj���вz�X�5C�G�([O� �f��ԒۛB�SOl��N�CH	��f��ϊf�E*g�NV�rh\�
h=NǞB}�!p��&��(_YY�gydN� ���VHѻn!s BP����(���ɛ�����;��W��V���I��n����k6�z��{��Ɂ��H�]Q�"�tj_�oT��%�	?��q��q�!��Tfx�z#� V eDN�����"m�9S����Rf�3���`Q�Y1�QC��Ph�{}�̭�k�h�9�+��,\6�7Op�f���y�|sVԒ�5?Z��]\Q�)/�q�{Y_��/e1��>��5hǒ�D������0Ỿ��
���Cj°�����S��!K�Fq���V�w���-h����P�e�<IB���d������`��A��	#�_�9��Э	
ɖ�^DG���aǶ �Fjq��K�v��I������`(I���ۊ��Ō�<9Y��A�
�Z��}a�'R��➚��c��x@x��ݨp�Ȇ	�I�m  ��b�}{>}g(���*�7]��rZ�Օ�壬D�7��M�C�q�TJ�q2d��w`�y�s(�uσ�.L���Ee��v$3^]�H/����H�1%����^.��܆�խ?hS��Q}�ũ\׮\�*�4�*u^�Re�B����ϑN�1Z��yW����\Wbo�,+d�?/�[L��&��܌�%���n"[d���8B?t_tq�S��-`m]�q�K0)槞��_�g���z�`H��h*D���71�U�H��^O���~��Co�xID�W<�K����W�����7�)�^����zP[���adh|�x�e�	���0�3���އ��'-���2�i5H	����z�X�; <�lө�i6�t�Mh���N�	`bVn��K�G:�Z\l�� ̕i�&��������v�T�Y_}}�v5��$�˕$�;7h��Ө?�_O�Z̓�����u��VM��e<>��m������Q���n!�w퍓���4��ߚ�ef�vx�,�(m0���F;��<Lv�����s��	W�ZN@��Mo;�܋���~a2����| �J� z�X�+����)�2��\�����q�ܭ볨���a�f���L��>����4�b�V ~���YtԔ�u5��+�ziR�A��"*!}��̅M�9	R!�7�M�P��љ������䑤�[g�:ם� �n�A<�?f#���O��5�q^󜒸u�,��B75��q���& ���4)�]O7`��h6߰�C��J-
��@G6`l�w[��;�g}ͭyB%C�.�,�&�ݷ�o=B�J�˧3� �������f�UJ�[Hɴ�V���"���)7��鸴�Wb�1lD�������KZo���p�j��B�d�����D����>��ޢ��8.�Ok�sK��+{��'?��6�=����L��)��4H�	��%YI�D����,�i{k������YKR�S����2�}�����z�VKR���L!�ӖH���l��l�B�QD� �-3�󢥕�9���0h��Y��:��2<�*k�mM���)F��6\�<�����c�p�8mrG|5��I�qL�lϸ���g���:�
��;��T{+)�� e+|%䁜S.+���p��0y@q�k��T�7�ϟ�Q�5�..��*���j~W6������[�&i|E�}�o(�:5��ɭLe�2���[�A-�t�H�<57�L_%�9S��8K\_zJ> D\Mָ�}�j�'㛶s��b%���M�g��G�n�K���z���S�|�=�o�r�W[��:��Gwy�&�D�M�dܴ?������3��� ����;6,�����se�2����]}*��':1OO3/?m�^�vm�;�4"�H���-S��O��@]��%�A�0h�&��o��켺�g����ե&�U��C�䢍\'���2�Q�>IY.8��g�5����t������e*Z�n�i]@s<Ҟ�v�.nV�79EU�w�x0�^(�n�)]�vKʖt�u��(����&jN� ��L2���o��(�3�M�Jۤ��v����(?�ț1[�����O�!�N�-��Kg�;���\g�o�`�I�H�������� �`Kp,�BP���__}�*���\V��t�P	�J?G��]G��2z�W�a�k��1e{>�UKݗ��N.`�x9�R����ob���4ʮ�������a98/�i&���#�m���ϰ�����@����b�R�B0ڵt�`���N3���g��X���K�~�7	v�xz�������[�%Y[~Z��2`;|�ጘ�O����;6&%�'�u�ީp]�p�Y
K��Ɍ���z��E�|>��5�=ܮ����s�<��'��Z�m�J���yb�:��v��Y��SqS���;�)��[�
lm�ΩlO��20t��}��:�a�c��_��,^�tg�`�*4��76c<}(��`g���ɹ�\����_��	t�t��N)1�>�
����M_������kW��������!�}��_�����s�,/A"�Y!k�H�-s<�g��;
z�w��C�z�+Q�O�Z=�]͋k,�`x�5��n;��*�[��{M��`��-���?]WW!��Y����p!ԨAz;��ۏvB�H ���1��?��WAK�C]�{*�xxẀ��P��:��:<�'^���ᐬ ���ü�#��^~�K_�[����QP���pk��O�[��������b�e�>0���?ˎ����0�F�d��'Kzf��c�����*iD[5+6���\۱T��)%B�}?����L].)�~XY�G�I��o,^#�}b�G2�~�qh�`J>%�z��LۦJ]�k��K�Y������	�H횫W^XƱ��f.���ES6��Yhe��~���^�_��HO�?�������P���6';�k�ؖ7�_��!�ޝR��v��#������U�(�Kb�U�7��5�	�N����PR�����[��g��7|�S8��dJ�/�C����<�3���KQ�2%�j#"��$py�۷�Hڪ���Y�n۳h�9��I�xqA�V@��f�t#2�%�����jЮ=��y��+��>��@��b��f˭u^,�cK��A�8�9�%Σ�+�:�dţ����44wW�m���)}DZ��:�8u��}q��D��M0���0�m=ZI3^6%i���O���fⅤM�,�m�De���V�`�.$�̚ɛ��$p�����*r�,{��W��Zy����N�z-cj����&oO=�I�6b+�$�V�#Z�e�G�s���7
Z�q�H��N�5e�
f��X���+�ܔ���x��mW��F�$r����m�n���/��
$��VPV5���Y\��5�>JF���/zv�e�Ϙh3S'L�G��f欄8ͫ���;\�ve�0����W�p�X��j����x!�h`�dI���i�lB��K���n��#?�o S\
��{4T�������Kk=���j�����+w�d�������2|=�,I΋�pV�i�|'Ҫ��9/�-J �"tA�/%W"�j�])�nSʈ5�gr���>a3j�����[�3OLc���zA2$��SO��1�VmvsJWm	�'x�Y@��>�`�vj�-���0�_őS�Q@J޻���-[.�|]��>�	�%�!^�N���}P��f?��-f1ǆ��VQ�9e��H���*��L�"���SW%��,?���˓)d�e{�m����uB^޶�lQ�-�p�O0�Jx�yQ�j/�Y�R> >/m���hW�J<��|���0e�ZXW� �F%���7'�c"�2�E�^O����K�����Ŭr0ԾkT��i��q�nT*�bB�����>�k���iށ��H�ĝ�!xW6����:r��l��� ����KG����=5rܰnx�B��%��C��w�Iof��0��.���M._T��#Gv��#�-X����3�p<oY�(Ncn�Z������)R!��A�WZ_��2i���,��hX��͍�l�mL*ݨpH���i���Fj�e!mI��B�IK�z�<9 |7�ueǦ[�ӛ��j�c������1:X	G���k�>�����5�mg�1��Z��hW���|g4�f"i�.���쏳�ޏ��h	kUl��������/�_A��i�m!=�%��I<S�A%Ĝ��/[,SH�cD��WOd���D��B�Y�>"�$-�fx^O����6���*)?��?���NYZ��zdT�j�k�=:N����&8��z��47l���������������?�!�����POR#��~!�p��|�Y�sx�����5!<�]�%!m�\��nO�G�[�<����ư��c���b:þ�.�?�/s�<T.D�>�9�G�4���t�\x�����*FB5ǉ��_�_����f�x��{I���ۼ%>S1�p��.��g����1=��ux@�L~�l��1��-����j��X�l.)�\���;1,u#��J�G����>�
�1ل��b]4�"�71��
b�"h�8F�<��{_j�O��Z�\[��ע�������`�c2���h��M��`B���/�D��*�QyZ4a�R|��)rɼ55|
k@��� ������K֫u����{�HTxW�w+yb�<m��aӧ§��Qg�3��,�J'w�+z���Fq���.�!{)�$f��eׅ~��ӝ�3���@
-۷�n��
�D$4��"�t|8���`Ϋ��X�!zf���B&#���:,����ە�����f��vWP*��v��( ��������^�a�c�q��b�KÆ�#!�ߎ����l�d�֣<	��N�݉�[�����f�|�G�5��$���f��;��.U��b�;���"3i���Iq�Þ�j��~�&�9Ƭ=�������aW��Aҗ�̆H0�!NP�;+����^��	�zʃ�q�ο`����@�>]|�b����,JЌƅÉ�w%Br-g��j�h����ٌ^�g���+h�ܝT���;c�L���`�ж�Jf�I,ȇ�\�vօ���H��hd�DI�2�B��ƫS�y����T��"�4�GT2*��w���P��:KRa��N�}u��2�Ɋ�I�����U������V�iý�#{S���Ka)*F�^Ӆ�ai��p��5����V2Plv^�H,P,��s�ĹD�J<��ݬB�l��5�/�x������$s7I�.q��Ռ��Z��'q|!n{�b	V��YZL�ڱ�Fc
�+��<��
�F��r��a��Qܨr���#������"e{#�ٶ�D��_��'��*&M�ĒkF�ָ��BTK��}���?L�S�5�>��+9F>��X���%ڹ3�I�X�޷(�C��u[.��X<�l=|�O4(�F�Y��q�W�������R���l�lӭ}�/�� ��(��%���x<	t�X���n�al�6��r=d�:�Ȯ�i�B��QM�ќ�{�)�A�#r�p����K+k��NX�dfq��
7��VJ�.at��Y0������@�X7;^�1��t,�`�'k��LNc�Q1�����n�E,�9�R.���(v%3�V�����V+xEl���W��K�*z�q����ő�v�V�,aA �|�(��Jb�=?ӭ���r�HG�E80��O��G�#�R�]�B��;j[8�ѯ<ݥ��uO1�+%v�t�YFUp`�1#
<?�S�<5� ׋��lr�7�s+=�"��qg� U�&���¯�i.��S�TVC� Sֆ%/�XD㫬4@OJ��`Jtb^cF��uml��Ƽ�*��x"�)���ɚ�ƣ{�@o;��'�cDkP�ؔ�e�
%���Ć7��p}Rq��ep�|��$���f��V��,����ɛi�v��-���0'c���A��e��سt';	�;��t��U�8`uG<�4.��s;b�Ɩ4P; ����dR���Ŀ+����5+[z����9��w��"��ۑ�/3Jk���I�Ĝ�D� ��]�@�BX���p�p��vfjr%�"��6Nd���v�)p�E��'��l�����![� C��s��ԯ���Ci"�(�J�P��a@��K��?��1âKbb�0&�{����GoT���e7/�K��h*㿽�Dnq�#��T�g$�)m�2��_���~��qLp8˪���m�lRCR����-Bu���,CU�N�w������2�$c�KV��:����,0���.�Q�亩7:;͠�fz�E���m��:��:i?�6�!ZUA_s0xx�`
w������ �O��g��Q7N�Q��nn��Hqx�o5�b��Pه9�\����NlQ��Н�E�kd_��,��%���aJ�1o+�tow�X0ڨ�h���/K0�0�V�3�`0e�h�`���ɠ��X��P�FD}%A�:1�u�6m�¼ʣk�>��l��p������S
��Vy�L�
�%�c��c��ق�e��=�P��(;���%`&E�UO�f���:�4d7T�_6)�]��׀u�����$jR�d���[���`,T�~�GA����#s�j�>�wU_��?��i.!�]�@���Ŗt��g<�V:�y�}℅r6�$V;��^��' �Ӵ���G�-	qx�=(��a��߰f������}_{�bBU��;2��I���ל7��$�c�(�C,\��N�hD~m��OIw�Xt�
�10C��
d�v�ۦ��[ط&���0�e�D^�Zʘ��p�`pMRP�AZ�y8�����Ź¡C�=9�
��GQ�B��T Kvu�:���K�j����w������ap���pyܰ$���b��3�/�?���b�h���hK���ł�Ϟ{��w���^-R�c󹤐����r#.ͬ�F1Y����Ȃ�09MI��®X�?�
P{���*u����LXoJ"K�Lˮ���5Y��u�����H�
Yq��� ,:�k�tm�����䃎�Z�.�JlX�h6bm��o�򒥳Me�;M^��՘r�oG�͢�0�+�<��yI½/�_���mX)'�.�����N��
��E)�%PHSe�9\��^�A���/Gl������ٮ�>X+�X�rD $�.��#��r�̊*��zC����m��B�oNHKCG��m���ݽW��g��_�q
L�o�-�m���˳,��RK�+��,!�4vt�J�l�_,В�B�Xp�.6��	�SJ�)3)�.Jd��[�d�Ie|W�w/���:q��{���:"�q�̡*��c2>� 3���5P]���;x�L�KdV��E���~�SL�abI376Z֝�V�ar��������W� 3�ǣ�!�
ӦJ)_��B���I_�!�~���l��< b�"L�4X�'r.u����L�"ֆ�q��.P��t*3#ٜ8|�M0�8�槉���X�{�+�OK�r��/���P�y��]v!jD�
7�Nڨ��JNG)�,.��>�A�gjD�#@W��6�(�{��Fr���I
��/ɢ��b:5\��O�}��"w���3E�a�������|J{�6�2S/E�5���_�9�Yz'� ű�ׯ0&�eR�:)��(�?��3���t��j�[b�OyP&kW��}kn��d��*(�bP���Ŀ���5-V޺��S�~���7~�� �(_YL�������,��x'�z��qmD]�I�*�S܋6�����
ճ���+���^���u�s�w	q�	Ck���=��z��#"1$�}�i�Ԭ�}Eh��h3����ʅ��ʍ!�(&��G�X8��y�m��-��+��ɋ���&�6	≩�����B$��K��{�S�6�����$lh/�G��Q�jo����%L���X��+W[H��2m<�]3��֐�EC�g�v����ȦٺH;�ן<��X{�xz��`�q�k�cN�f��^]�0�g���V2.�EC�����MQI�p�2�q�/�p��z:y��u�͠�t�~c�2�̈́�:6s��:������5�Xѻ|�����U���
��s��G������%�NE�F��;@ls
���2|�QrR���_�k�$��y�"k��(^�a�>h�X�>�J��[5��ׄD�sY�P�g���P�('N'\X5*��D��ˬr�m����A������a�fO��~�=/%o��>�*��1�K�3%�o�#>�Юx�X� �vmL?3tE����uѿ�"���wh���#�,�����x�͢�=��ɖV+^a�9��KܽM����:lM������c��%ۈϥ{;�~�ٿ8�Gڤߪ�Drj2���qD6Q��f�*[ �(���ډ?jz.\2���沧	���c^6�Sӫ5�.�}>Y�-�$`Gf��誅F⽓�Q^��t������G���	�u�5������%���m�������֚w��H�;�Z�TϳٝT�x����!���3 �)Q�����HB����^N�5w��O~��	}��P��ep��0�-T�ҧ�:cx�r��v���O��ë��������;�����˛
�^v�����]�\���{�+��OI��]��g�|�B�G���u�Q2��Ws�W��~�|V�� yXa�Q�j�<s0n��X�$�:�����s��{�I\i)��P;Yi��"�1+�g �*=Ul::�,9��o�P� ���T�z�!�3�>OޚZ�����^��,ş]��@�^���̑�����f�~aשN[��������� ���4�:e���⧬e�w��r.�I7�$���U!hf03x �r:(�UvKX�.T�>����T��s
�Fvhk������e��**��;�n�����z#W�Ơ�m�G�C��m�ﰠF��Mn�M�����׎Ƞ闖T�2�7�d23�P�- �M�H>9v��E(�o�s�Қ��П(&��P�v�����i��ڬC��Hc�<F��^d,,/7��*-7'&����l�D��j�P�Aͺk[ ��4�hzӽ�ְ%˲������H8է<=V���N-����S^�-5���c���A�Z��&hHi9G�T��2���kg��#��^yp����x��l�1���lS�#E�c��©Q,P9T3\�C!�=ݗGd�I�)��Ȥ
�nb�B4*v�%w��]X�+�E�i&��^����Nu�w�Y�5�����'1�雫�Rί��v�ܟ'7|��0�Ц_����w2�����OmpO���HT��T}��΅Z�TN���o= ϲ��Y��ȗP6_6݅;����E������!����P9�˻s�jf��4]��C�̊���.{�srJ����Z�A9�����>bb8�E��S�T^
dY�sՠ��1!O��?y�O=aC��O<H��A�����J(��5abQb��S2�q�zt���W�OQ��G�(����k3�ݙ� u~�r��~}q�ה��?��w���7@곴�7��O����!�ڌ��(��I�r>�t%���Fu-l���s��Z�Xj�i�vpt�Yv����iN�I�$6fPw�G�uC�1V�ԁ��A>��s��P>��ے8g���_��I��*q��]�^�DþB�JQܴ"V����/PFGZ^w:Nk���$���ߍ���-d��üK
kEV�E�;X�� g�\̈@$7-Zr�|R>�H�C!�tLt���d
5�7��m�=񾛜��vA��g�J�[&{n��6�h��
�h��H͏1�����Hv7��"��3Q:Z9�����N��F{2,�N��n)T��?��H&��p�v��ы+�kF��nK#WZ���V%ɤ�k� ��̘���n�/�!�뫡�t���W7�1�N�ZB�12����1�AM�M�s5w�A��t�1�dd�y,WEl�*��8lُdH��"z�h{�0��ąYK,TY�j�
:��ӫh ��̹���L�@�]4#�V�9��U��s\&cEw\���
�`�v9�'!i�@MjbF��'$o���Ɯ}/L������oGZ�v��#�_a������!O�5�L�x���ʖ���;��b�:Bёi,�(���v�c�w.�Q`ڤ��v���&��_��s���u�h�ٙ��D���4��ޮ���βp�c�Qǧ�^����$��<Cn�E���DJ7���\�A;�/>�d�݃tKݼ��?w�o+�"c�S�h@�����o����y/îuv��k��f�o��� }�W���'�L|�ܷ�u��n�Ɓ@�p΀�	ծ�:��rk(W`/a�r �/G�h����9@�S��nl��iɢ��)��ooM_KL����}�-~�t6'Tʱ��2��W���Ʋ���j6!�d�����8��͇H��E�T~:�#$2����������Ȱ��gQx����o`���9l��H+0�7��n�蟃P����++��k��'_P_Ί��ct(hM�㣶2o��QF"e��#����R���?e�i��6w]�t��ʢ���@�*�VXq�Z����Mt��� `{�gV$�
]/���F���㌖��&��Y�A�2��$��fˍ���5܇��upS��"�q)>�.Q!;�Q�(��Q<벍`+`"�֋����Θ.&��>�A���c���ف;�QB���Q�@�I��qJ�����;�,���q-B���G?��V@�Q�MZY�=����~��2���u�,����'����d![� 3��j���92�8�/d���6�k�"S&�`}��PG�]=�zL �N��t�>���F�Y�Z��(Dp�^fώF,�s��J�D���ȓ��$�B��W� �6+�E�� ��T�&�pD�Pz����]z��A8��Q��8� ����T���g��L�L=��~C�Y�&�8ҕZ���;7��1Y�;��O��������*�:�jx�%#��DNNel�ʲ��ҋB��M��.��� �NVF�˻v�W�?���N��r�����*w���W'9�F�����;#9�q>^�9�����0�Ws�6T��#JX[~��T%�?86������C|����g�V���~��f��KBx� 	󭚩��+fCݫg��[ݶNU�����V��3���W���w��v�=#W0l�Ô�c$yqnyOeF�WY3@��T�Z���e^\��C'��S�#��=zV���{$���PU�ø�2)+�4�/������g�b���������p�����+�2�*�&�{D��iHܱ�������7���V��%'�FJ�&�~�b�����h���������c�s��1�o
ܭ{U��K�n�Z��\WL��ae���K�[�'P�mr��\����oP�ʳrV��R�j��b��`2�9
��^	.��`�d߈�~'s�y���פ��x$2�c���@:�
�8��1�p+x*>z>L����о�5��3=�jQx���SqNp����.��!G/�z��{P���!��
���x&��D
玩W��[�6�q��ԟ��':���I5w[�x_��.�)Px?�O�G,4o�F2��inD��ɦ��O/�[����LC�k����NkY���UY K�B����R�v[@��:2n�}��S��n@+ϱ#�����U�Y���n�;׼��0Ly- W �Z�~�yV�R�~\���`�f�����t�R���$/�M���ώ������E�=b�\\���vQ~Ͱ*�on�(�l�z�(� X�r�$.`1Z�g_���>rQG��h�g6z� ����0�:�!i����̙ij"�ɍjM28�؀���:�9�@�fW�LT�d�W�	�]�ƫ����r�`���E�]h,w���y���%������Y��.CsjGޞ�Db���XV�Ay����x��qf���'�O8��p.>����W���&`,�}Ml�,v�=�V��\K�X�R�cW��H�ց��EV"7056J�.?��]�OO�r��_�tg��{�1l�����|�i��ƌ�V4X�.)-T_��F:1�T��"�x�	B�ʥ�v�h{��:��L��ܱ�b�� ��_�@	��l�'e��
�d|�E�f���� >�xB�D������|Y'�i��#0��L�ɟ�w�g.Ѭ*��'nR0P�B�-�ᕬ�c%�NK����a�]��Ƚ1�P��d��o���
�R�2u����Ȏ ���!�m�L�jjB.q�d�,�
U�t�v�-u��<(.���F�8v�qnNrrJ(m�#ST��J͸L�A-��3��ha��E(���|��\b��;5�3XDUç�\��KMG��	جc.�E;���XOXn*���}֡*��N��r��>t�V��Z�wE��xa�T���p�l�*����]6�@k��:'Ќ��fb=�\�EmU}'��qj�FO/��Żd3k�D����I�Ee;q�|�"�I�*(WD�U�p]�m5gQ��B�Hs�X��w ss���e����*k�l�c��{ ��g�MёH��s�T|������A�����G��bȎZ>E}�kr�r��R/�,�$����"<���@�������^�4ZD��o����R������F��[�u����fѡ���:��*�פ��{� �oS����g{H*��B����*S��P����GWK�Nbi�뚖�+�����GV�G���&�i�>�<�kj17C<�,yF�#�9�����Ϥ6=/ ��H�FF��M��P�t�.s��>�<�&{�o���/R�q�!���3ܦ�N���.�ܟ ��g��.�~��Vb�i7����=8sKU�v���է��A��	%	~+�|�J׀���D��?.�e�,�i�ՔXxO=�_��?�|&Q��Y�g��:+�(�
�I�^��P���Iv��� ��Se�4�a�m���J;�)&�N�2���\6�6���v緲� �q���@$���*/�I1�	�d�1:X�.
:�]�u�����)&I���GC�bĶ:]U�sz�nҮ[5�����I��@cb��b�.{��M�ZI�� �Ǻ�x�-Bby�S�K��f1�+���6�7�I�G�F�}�@�/u��kY�F4w���/)�WC|_Ş�h�kXy���"UT�ѣq����� ��k�]c{�3�>�ƴ��;���]�6��3�8��ץΙ.�T�@_�Z��GI�l�ses������=-�����f��0~3��gР���p���nQ�m�����3ۋ��W䔚��@]�Ζ�*_��l�֤XU٣~����,�{f�i�Uz�R��4�h�Nܞ�K���}߱�F`�7�X_<	_d�t��֘��ts�P�#��Ve[����K���_������q\��� ��%^�>��:0N�Ԩ;������K�]C� �, �ne���<��Ձg��e(��۴}�e҇7,*T�!�u'��H!���W�% =�09{O�/���h���xxM�,�M	;�8౱�w�=�rb\�mD����&9�5~�fiL�o~�p�TQ��U�F��yM6d aA9N����."nΒ�J�h�Ai���C�4���苴���0	~� a2�뫏]֟t�#�Ͳ� b�B�Sߗ�it�zj6�C������Ks|�3�@ZI����HG�x�)#^n�4r�+�`)�,(h��*�Ty����5��Vy�%}]���7�8֢(9�SKKl����}�դ�cs�_� D��1%��"��b$�O��K���>m�)�V���3|�'��%iL���N>�6�@��@��[b���]r���B/�	&�f�NfQ��/*�֚��zU��,]sMa�靂���ϙ �@��y�
8m��H��v���������6� E�Y�E(R�yd�39��p����R
�������>X�߱�_/Da�I��"&eTH�`-_rbPR�Iq�NW:4�Epx�ȱ�t*��_╀Յh���=� -�C��V���6��V�A�mXdq��/I�vO�pr.�G��3�(�)��F�|�'��=��d��vЌ2�X@ʌÒK4qoW��비��M��o|�Y�rz��c����imI3����weo\�%�Ҁ�JA���b�[Q�3
�˶u4�|4�~�EN,y�*�L���w袨��@�޽���Ş��q�i󯆘'��/����ԯ�C�.'x냦+�U&İ��e���h��U��"ck�SMo�0 6s���o�`�V�@��'���)�%��>HL��Z�M�V�߀�T��a��zv"7�^�]�b��;Ϋ�o�������n����r�09x�;<�BU��ةjRD}���>��_Mqo�Vu0���\��y�l��G�e��������4�/D��˧I�)����5�4�巤���҈�E�W�&��Q����� ��Is|��E���=8�8?�ȝ��^(�`�n)Z�7�z�<�т|�>zk!��P���Q�혹ϸ�SJE��.Q��]�چ���������7:��`_�����14=q]��wKՖ==�,2y	A���ت�2��j{�IKV*��L�~V^�I��� 8�Ui���Z�����e��Sj��`�|6hK���_4��:S��2��� %e뺽M��S0��Y0�����]�9�$�A�i}��QP���Y"l�liP�eUcX
�(��5h"Q
��1��� qf;�l�+�-$�y};(������Q����ݻ㹿m`��� ����M9�����x��,]�f�c���G%;�Ĳ��Z��<��G4P[u���pҡ�pG��_v j�v��'qզƺ�@���L��_�.�U���]�)�ן2�F�{��o�P���2���e|d��*Q7�E	�I26]��+�[H�ʚtW�_��Ҥ�~�.x�C�ۯ�ڡPu�fT���J`�l0�;��7 ^I�1� ?���-���O�mk%y��Lx֧=vM�nkw�-֥$V��^�>��q��9 ���N�V�
Elx²�k�h`���*u./?u7k!
D&�"1����������W �Ԑ�8����¹Nog9O������$�!_��O���fj�ŭj`r]/P����AF�&�V�|������`��-����)���kxߠXi�ʖ���d�73������k0p�c�A��=���t�zY+�"�(����Ff7����%��k��Vy�d�?uw�p6�e�#����fq��\����\� slـ¨�ӣ�sr��e׬g�Z�3� r���%?��z�?�з�� 4��ׄ��+^�U��0g��K�6��_�S�3E�#�{�<r�S��C���^��H��lE��1$�$��D"^ԴWd0�S�=.�2��vQ!�R��jٹ������$w���,�2ڵ7��b9d:\s��!��_��1�����C���{ki۳W-IҌ�*a��?�H
~U�l���|�W<	<�Ʊʞ�����s4i�9�$L�Na=�]�+?��#�.��"�s��GG���J�4RE%ƄF��c;\�6�*T�A�9Q��C3U��[QJ�_Z!���n=�ޝk$)������B��� W[�t����%��
t�*��0$�ZS�-�qm��}�H�˲�Iq���0�z����gRw�a�*�9{e}�^ɋ&�h�����;$W4-eB��S��:#��*���Qj'%�zL��vl�:h4:cQ7��˂*	H !p�����r���*ML��d���j!��/jK_Me���ԾWZYt��J!ܣr���s�P��<�JF׿���#�I�;jNaB_��$��2+~*s%i��>��L�Q�A�s�6���߯�  B8�xT��e���V�5�*qv�_k/�}	3��F[Ĝ�k�Qo��(i�c�P�$G�x��0�gT]^�_�HSQM�u��g� � N�lѻ;8��2�D�礿��rF�������+ȕ/���QsyKqc�]�_�gR��+�S���Hd�h�yyHRW#���H��o^�XP��u#h�����Ok�����փ�?�6NZi�i+�����b��Or<|9��\�:"�����˚�A�x��(�����W�_�	 h���j�/�#��Yv��YR?3
z���Ԋ�-
�
Q��^FO���)��0����G}&��|ea9u�#|����I~�<j���!��j��ȳM4�w�wLV»����.69/�i	(<#�2A����8Hmt�u�=�� ��ӑ�&G�|`l���E�c�&�Y%f�����:��(0a���Q�>sdI�u�j�/�� Z�'�9����?Я�h�|+%�?@c����U��j��~�4�+����i�����j�2�!�g�ݫab�"}���#}	���|���g�?��DӽĽQ��=<�1�� �vڨ"�Ƹ
}���f�����
"_)Hxr�����Z�1�7Qw�3�V�<%��83���^�u�ӭJ������^�?n�b�ul�o��	�K�zR�^5���dը���6Ն0�����6��x���v���&IJ�3�|�G�tjyj $�`my0��.�_�zmX��g��9�;Q�U!��B�$��h2w%qZ`��l�cT�:a��nhDl�)a%As��`�1:�$�df5��'pv��KZ���~���4y�i��xob��Q��Nui'�,6�4U%�� �<�fۂe��[�RT9��3�j����u�Gυ��&����+.My�G�k��o�%A�%s&<��Y��p-xӌ�m�C��z7�ƽ�\��Ѻ�pM�w��tEC$����he*�U!YK��gR^{Y�.��zr�]��������s*�P٩�	���-o��7�t�;ZXmQ�RnNo% ^9B��f�>r�\�Y/�#K����)I�����C2s��-�!9�2��i9u��+Ȝ_�؏�E����m|�����f8�/zC2�ؐ�j�5�/�[Y�b8�I�z\�R'AO��4�}�|�¼X�*�镭=���������- ���`Ո��~�Qیeo��or����wt��� �߽݉#ɡ[t�ew"�Kԧ{�ͻ�)CM��N6_�~ՠ�F��d���RU��vŜG���\��:l�_y��k��1��<VEpDxaqpf�~{�=��Ty��@<r���T���?�������P�p���'��w��^N�����|B�L9��&��	EX������yVj����x�?M�b��q�������"4h��4�zS:�;L��a��5�`����f.	�te
rc��O�����.z�E��\T4���푃�4���ȶ���7^�,��)PU�1����Gڑ1�>TB�_�_�������ݲ�ެ��~�ux�O��6�̣G�Y�"�rl�"r��Ip� ��Bз���(#c�L�������x��Ӣ���ڱ^���.f/
ßZg-q|�v�.@+�D>�Ƃ�Io9_�<����0q�Yf�S6����s֦��l�'�F���i3�ru�_��8:P�v��G��{�7�nfI�/.�t޹o�I��P��jL�J���d���|�{V����HlAĆ��^�j��].N��܆l0�Ti�㞣�$�]�:	��X�9q��>�`k�_��S�_u���`��e��{���/i�: �o{*&�r腖�^=�&_mi�1窎�25g������Ԇtt/>zR�Y�KnEu-��!2�aJNޥõ�:�[!�+R���K���؃�\�ϲ�B/i�GUĎgїRڞ��ݻS���p�X��K�| �b���<5��ˋfG|F5�?1����A�a�.nz�u��Z.���C�F����e�ꉦ,��dQָw���^��n�sr����u�,;�m��?�W���T�,�CT�X�Wz��f{c�K/���4.�J�L�N�YΜ��_ܹ���Yq\{=j��<a�/��M"H�jvӁ*������2i;j���bܶ�Av����	q����2?�2�ө)�ss�t�ڲj˨����Xp܌�7ƼO� ��۬��4�{�o73�� ��"�u�ݎϮ�a#��a����)�f�fl���%Y�65n��������΅��᪅�b�y�����)�wA1A�]���j��Z���TC8��RW+#����s�&��Ƭ"ł�z���X�F�6��Ү�bH�l�6�A]�,�(��=өr��8�?m�yY2a���^���:�7�e��m�dO��@e���88Gd��s��!xJKL�5f ���Ƙ>>��K���������a�v�7���n#E� S�]�Ҁ���[nkmb9�3�G"��<4��$�.��cDj�ZE�R�$���c\yiSjz���x���m�i
d;*���AS��?9��';�ؼ�w�y��.(<��>��
fǘ�I?f���֦�X�Mo&�&M�hBpf(�E�]��hG�2$S3�t�u�����V��/S:�&*����̕G�Dp� �ʓ9�� ? ��)�0��{(���D@��++���|&��8^�u.�h@�\>��S�L}�̳�2P�c`��^�g�K&�
�Vc�QK�]U
��Ṿ�ƅz�=.��/u�Mzpf;��t��˩jLk}S�i�=�ݳ��p6��q%d�����2!g<:kDNc��\���W�G�a�2�}�L��^����M8�s�yCu-�
Rk�n9�H����Y �{C'�~����e|Wd	��K}�	)릲T�fP�^����Y�q�=e�� ��ş��b�S���i�&9� z��,����!� �<��;��y���ݬ��|���+R�$�������qӆ}���9�%�ϒ��w5N���U@������c`�A,}�|�ӣ�4A�V��î|�Y�GjǙD��j\�L�%��G~oM�QU��sF6���5J2W�E�N�t��N�����m9�?]٭��L�� �E<����P�\nJ�O��32�F���]=���\7��KJJŜ@Z�Ч��L�q��b�E.u�UH}Q_��J1o����!+;㽺�ia�T����'�����H������n�?�o�_,�`�9������%E���0�U��Nuxý��8�x������);�?CۖI%��iVM:�H��^e�d�ґU?�ܡ�B,S{X�4��{��r��)�\6�!�>������1�?{��݀��+�2���Ƶ��FLSxCڋ����\��ԟ�7o�斕��� O�\|��V��K17��ei�[�:p譲�eI��D��p0��L�5q2�G,���oB��sn�6�| ۖ7�^���w�!��R�T+�;�{� ���0VY/��[���"!�꣌��O�i� z
4�e��]�	u�(ų��Z�'6���Mb����R"�RM��\��3�`��o��`u"慯5��O����'��\��~U�(��O�U����#9���~�w׻���-�U쪴�gy�{�|ߣ@�J!�i�ǜ�DN�Ɵ>�4�������b~��I�oO���?M����03)�M'qF��~�`꣜�d��M�8�8C[o�a�*Q�*�{v�`9�����pr�N�q�d�f3#��ͣ�-�{*�8%�!;��	����)�t�u���Բw�1K[>����c�f������`���H�[���s.�[0���5��� F��7��CҠ�ӵͳ=�����[��骔j��~�Q�h�U�#_��,_#4[�0/	����Y ��{�U%aY����&vI#��lz�ɵ�/�r�)��:u/�� YгɋA
�B�SD�$y:��`�p���`b���'��)�L����zs&����OW	��1sPp�;^�'�v�n�꾲D��g`sr�ʁ3;I1hX�W���=\�}�}��u6�]|�)���\F�hE����.����7�/E�G%���k.�,�Xȉ����i:4>I����8*����Y���%u؋�<z�LE�7��G)%}y�b���[��2�zn3s}e��k��Q:���W�Q����� $ΧƱ�NZ��ǌ`A�-���T���>��3�r�B.�����7�%��Ͽ�2j��*�EEsҢ�$?���A�"�o*��K�Δ��Y�L�]��6����|�6$��yS'��	���i��_{r
�\��K�����!q��>9��7SE��p�(�'�X۲����+���#�V��i�C6��t�d�Q��)��XfM�Vs� ���6~���U���
,W��aRz8�ev8�����fV��&(���N��9��H}P�upFR��"+cw���Ll0uay\搦m�F�P�����t� 28�c �m�x�~t�[�
�d+���QI�rK��V���`���G��E�c�b�n�s5E�yQ4(I����#�p�9��<C'���a���P>u��AN�����5�4����l��.� ��U�5{aO�`��P�b�G�4#��?`aab?j�ik|�%ɠ�)�m/~x�D�	T
�S?qy�y) \t� [wo	�$���0}�A�S����rr�ܟ�{�S;�{�93��{�)	H�p���/�Z[s�V$[#���A���0����y'��=~����A���smG	�	r�_��NG{�E`gbT��}i����;�&X&B/@�P5c"�疢�|u�N�^�U����눓K��!�����s�vr���ѫ��=L�N0W �_��k�}j�0��J%�7��ҪQ6��0��}�9�́0F���]R�Z�r6��IBo���x���~���J�=�a5蓇B����ԗ�p�/���z�mR<�(��14��?��΅v��t�F�	"5�.���`Œ����^�B�b���^j�"<W��RJ](M�wn�4_�R'��,έg�� ��:�����^l��X�%��P�����.R�YR�c��4�F�F����`�P�e'|���K�P����&腅�in�9��,̊�:�d���%A�-F>4T��7?E�\�Km�nV�@�߂'�(�]�NvNR�k�忠g���y��j���t+s�jz�EAW��h�}y���䣁���$ˬ�{���{k�+��6���Ac}L��4�5�Ȼ�H�G����q:�m���#aB��ʝ���E#��ۚ�5\�l�	@D��(���y���u+�d�NK���4�!����go��	���ň�g����p�'7�x,�"1Cn������S�2`GOå���i��(���!d	6�R�T>m��G���#C_p��"2�'g	���O�lr2�J����:A�/��'�q��de9R�{p��œr�Q�S�8Gv��=~߄�n p*�I���c3��ŕ�?[��̡_M@B��<G��� V��v�����%K����&��`����BȈI*T�}d���.
�7/x7��,Kc�����6@�����xA�P!����Q���^�����k?���P���E'�ˬ逺%j.�l:�Q����J#�p��_�6R���������\0��<-�����p�֡�=�h�q��j���@�3���PX��x}�a����ъ	�|&���d��qZ2'��*�CDjYްɏ/�,h���lL��>yA�7_����c�"��͓;ܧo��?<���JU�*ͮ�ci�JR���-2�,�(�۰ZU�MC��T��qwzy#��8�������"�(����A��1$`��m#]G�<��[4�7��z,Z�mF�I4k�����nt��3�#�Y��]���ˊ4!2�,��%� 0���!��$a�	�x^PZ�ɍ�p�H�*E��ad�hrQ��z�60�PE5FJL�̎���R5w!��S��y];58FU�H������WB�o�N��s-~��#zrR�P.Uq�$��� �@�<C��L*�pO������� #�'=��0س�����U=>��{R�v#�f�n��(��'��H��y�9$��[��d�H�X�%�Z0��R?��nf7�&��$�xk����V�Ê+Lx,�߂'�$&G�-3D�Ou�x���_����YcIߗ�d�H~�}Ӭ�j�]�k��{��md�`G���8x�zk�>��:}��$\V��H�k��h���S�n@���/�7�ITt�ɑÙP���E�_j:�{v�q�W���t]hள���CEoۣ��}c��T﷍@ &��%���,��gX���h�MJ��cT�/-,����`q�S�CԥA3�Ah�!j�T2�����	�!�X�[�6`��Zf��814���~8ȧ�I��h|>�{�&R���޳�N�\4�� p�i���s��1Ŷ�^
AY3.I)B-h�X7��C>l�c��u)���y�!y�8�c��g_����BG���|W�qF�w�<��c�~�V��Ye������I#Mq�zT=ǜ��94��	p �KO�믔B.u[��7Z-XyX~a8>ђ��eC@��UՍFޗ��)�<3����@���R o��Aw/���0jT��b�O���� C��$�i\:G^%�Z�;�ڽ�j��Y��_��5��5�L/yek���ۤ�GG��bO9(E쪎�� P��-zP�󳰛�fT@��T�d��umC���5{N]m�yb��~g0|���ǈ�.�o�y��I�`���^�2!2c��:<��	��.�:�!����P/5�-+ƽv����r���>Q�/��t2�`��*�r6X)Na��X�J���t�*�77i8
n�����(1O-&4IQ;]��M�/&��Z<S���Gv{��qQq�䕑���>�Tk���jf�2+����3��4���ꔗ���*"����U��0Y���B����s>H�- f.@�E�����F�}�A�%Gd؅75��H�|�#L�c&ua���MZ��և��_�Oz��g��F\ra�ou��F>��va[��iH\^+��/��W"���I㌄s���U�y��'��FUJ��0;�Vֳ{ϰt h9�-vY���Z�9)�7� �y����
��59��HLz"%T�3@��5���Fa��+i �mΌz3�vrwsΚ)[�V�Q�pExᝑq�aj�nR�B?So�CT�?,>����x��R�����r�pU������Q�,�5���a����];>Y�/���=:Wq���s��+�<P��3W�ҡT�lD�Y�E�����Zq��šB]Áq�ؘW�Ws/7"}�I���PPx���\�L_D��e-�"M����uJ�E�4��<�+z���T�����𷏕�x|"U�����6}�#��5���{d�p�ϭ�s`5�uD��A��|b�PuH���mn�c�0>���"[Q+[������oI~�,IIBH�଼��k����^�?��~�h�	x���uǖ����l�Zk�X���k�1�H�� ��R�w�qB(�>MwDR}|l�%�	��W"����!�6�G{�6(�/<8Ǐ�����MDD8.�g��u�6���Ol���۽Ωd�T.B�S�������f�*b�����])S�⧜���	��H7}'����܇���=U����� �Uك�ߡi�%}���6g��Z��BA5"��v9��Z,��`+o���Ŀ���M�⸟�J��f������M��!�,��߂7���<rmo /���c�X2�PM��v9_�������n1�����Ez�x+�J'�M!P&��\;��l�0 y���P�� �i��$=z����u�����ϳ���	iK	m��w.�t����Y�D����!��&��C�8�Pv+�c}��9tom9bR�ބ�u�җy�$�[�~�vT�RԄݼD����վf �����H`J嵠����:z���;.�i�l�O�WE�睚�:_=����|�C|!�
��(�a�$����JČ�r��p��YH�HaZ"d�3{��M�7���8|�׻�����f	9��>���|��YG�6YTf(�<�]Rdw"e��".�B�%��Ơ+7NjTO���$�%�#��@������r�L
Bcg'�_��
����L&�e�[a��DD����l/���p�M:�]�uX%�{D�nX�!��t�^R|x���M��^��hc�%"֍�T&�T�^�0S��ղ�!�np�F���Rn���H�-����u׃!A�:躚�	�n,^&�iɴ����
��qyߙ�[���T]]brnb),W�F`�e���d(�G���51��b��nj�^�7z)o��ߣ��^W�b�T�\��u#ޠeҺ[w��k?�V*�eUR�v���f��R�����De�܃a��z�6��i�]G�%�_�w�7�ڌ �}1@�n��lW�O��	0v�ń�@�WO��& O.�j���"'U����cu߅�O�T�h���
�J�؊�@$����V���8���1��Fy�L��|<�T���A�B��l���֭�y�������B�d2�	�!1r@}�tI�i�����4��J<$�>�@��6�?�k݉o�ž\�[�F��Q�5��"7�7��Ҕ�n.���h�1�p�A�k�D؅�'�x��狱y�v6�kѳ�GK����02[DF�z�{���m:�O���خ�L�0�)|�K*[��+������3����B�R�gR�^e���K��7ٌ\v	�,�W2�򚊈���d�����/n�iV ����H�J�@�O;�箾r/�O��DG���g�� ���K� ����$���ʜ�7�s�=��pG瘔~�^�r��W�¨��gJea[���%}�`_΂�$�����ֵG��ك㹏V��Ր�݂0i����S��}�(4���Q��R]�|��*�Ƽ����F�D�X���>�j��љ���Z���h���IVL��E�B���
C�7�|u��#��77|���*��3R��h8�Zs��L�����8ݳ���m8R���4�z[�� �IV��@�F�K�o�(`	p��d@�qkK������\�݋)�d~�H¸*�4��`+�AD�����(H�I!G��苔��o�}צ��zC�Qb�v98�Ķ��8�e�yܞ�#%+z2I�8]6eaP�*
�1�ǅF�W��(d�}���;j��4:���&�&�-[* �
�J�M]���rb'�&"?GC茷bG�J�O@l3V5�jF�[�ؾ�gY|�֏�$�|gN��I�m?�޷g�p���x��'�i=%����b�"�s1�"ڣY��*o��a�i��-W?�)�/7�䲣B�S� ��b+�	�Ң�SzX-SP_!w���"�\��ڤ'�3c�4��mY�ϖ����:��׿�XR1��.X��v��޷P��+�W��5���VMf�Y�֡�Gw���c��ɻ�90�7@f��,^���s"w�b��?T;�������g�l���T�o�J2~�K^���N:�'tL�l򅽿��;���9e�"����6������W�?�M�5h�籉>�3ޣ����B��̀J0��֩�0xN���E_FC�i�U\��G]�⟍y��M]mLY/S?��N�B`�\�8$I�`u�;�^S7�r7c� ?Q����W{��(8���I3$�����}��;�8����q��C�0�����b�z�|��7�]��K?N�����ƈRz!g�������E+RpؾF�oݓ���'����IG�33�C��&i�b)�Z��M�P
Xl��ɣ8hQ#�	�wOq�K�f�sK��}�!y����a�f����J��z�c"Eb��H�g��+����Ou�8�V�B��(OoG0$�7�Xa(�,狕�
��C�����N׃w����ns	�_z>4��X���v�I�M+��k%&s�G:�F����43�0Dh�d�3�v��}d��Zy� :[�AN�1��Ѫ�h�HH�(����.���>�˾����]��e�b���$�;PO@�$S���Ģw�|1�g+|	?I^&^r�u��1��� [�.��� �����~՟�h�65pTAj���-1�i�`8���=y�;�K���XRŰ��["l�47��3>�
��O���?rdY��)�1�Y��ҝ�WU���pTU>N�#�����c���v�z��w�\l����;������vܮ�
K�s����BIJ��Ԭ.LEZ�3<8�Xm˸�]fo���A}���֦�!��c�ᘜU��O"=��*�-�/�#_Le!��٥���+�%�-eIs���	e�z�B�����z�u��OKEe��)�,*9A|=
��Q|�Hk���͠��h(7�/���XC�uD�4�m��܎yO����BGg�\��R_,��P�޾���gA}3_��9�]���%� �"����7a�YҢ��d(��R/|QL�ѯ{��ٶ�`����F��j2��S,-�T1]�$$��s���J��%\+<����w��]׸��@4�G�����)}U���� m"n�T�	ofS��by��:���Oj���圷��=�S�YcA%1�듶�2R��KY�z*_�Q��/
�_\��0�`&����hhU�̆&2��m����Y�	���{����U�ߣW*k�q*�K�'ۉ)�}�CtP����~9��x	�Wpμ�pH�7s)�%��E�S���#������W����+������^�y������cy�����ι��g���Ѣ��<�ȧ��ђ�z�\����:a�x0N���Kr�%�����[�i����]��9�k5P���jo������k�`�����G�'������Lz�:*���83���p?[C�9.Ո��5��އt$�?u�ь���"�E'+����|�1Zr���������1g��D�V7�K^��&��'���-",���-�oh�����?b"[���&�"Q���Zg�5��^ξ}�����O�U��GD���9E�,GU��y[���L��V?p��'�8�d`�o�F�mJM�2d	��� �d ������D`9�x`�ȍ�e/�b�`\� J�OL���ڱ��x����y 
�
5�c�G2���s��p�����/1���?|z���E�'��m~���q������va�t�$<OȈ�=�oF�v�z�Y��K�F`)�r���hb�-����z��a�f8Q=�v�' d�`�XㆭP�bi�w�7�D5��F�������I���>N�-f����?�a�������Su�8CM?����R�$?�)��n=������_�%��! c1������C[gep��/pkkz 8���9`j�z��(�h&K�ĝӨ����������N�醶'9�S�V�/���wM�)7��qK�U��y�i��e��W����,:?ƅ9�1b�L��{�Be��
g�m�L02;P��{'M �.X(���M��,�ܞ���geʩ��8�D����û�D�ܮf�g��N׾�)��Oo{iE4ʓ���O��u�a��E�w���{�U�#B*`�'��d�',7J��4���r��nl�_KZ�F�F��-��X���1�B�y�:�I*�@�4��k�XBC�.[h�H�]����U��do���N�eaE%<��QA9b�C�ܜ	���.bK��'����$ �����a�ӡ�X�oY��!��-C��YTL��c�$F7"e��6�x�lC?�I<L�a|����k5�2vg�6HU�@���/ܰͨ����gw읳��S��2�'����<( �ҙx�"�?�`@�k���1A"������ ���(K�e�8��$w�u�0��9�F�"��fԁ*R_P�b��M� f?%+�f�qW@R{�jlKa�&5V25�n'P(A.�6}��?A�%ɵ�V�qf@E���鹵����_�gOcCT��]9y+����*������am]ǃ���8*�7�%�F�iӷ'�'84�c��@�*��l#��y�	Q�f�N����b��_�آ6~f�\0&�E�z�w����I�\��qi�8� ӊ��?����D�kԯ�?h0U�*�R�l��7_��{
�x%�cD�##&�y�i��C�� �n��el1���qh˜�,Hc3�_̟�i)~�wZ� ���p*^��>�]!�D�/��^(@�=��#BT��[�"�c��붏��Ӽ&���\��u�* XSѧS�!L?)�z�u.��ca
�䉂	UG���e�b�P`�ULX�ߢ\��gЦnջȁ����<F��
��:��ޅ�cU�F0Yg����%�IU-��CC0�N4����C�/��G��'EnF?n`�q�^-��w�z@�YS6
��aG�PC�rPX\� ��qa5�AN|-�\C%�(�&mr}�:o�(�!L�U�h3gH��*闿�5B��_� �|�F�5��R�#��x�n�8�l��
j��U(��
���$V���
�*\01eu�0:(�U�9lc]��l,W��j�Y�ȋ�'~>�����!�N �r�����ܦ�;w�b��ȧ9�k[ׄ�|�ĕ��3�w#3�So��N�R������I�Th[����{�To�i}k�i�����4b��P����G월��8E���o�26(�j.���П� ���ݏ��CjO'�V��"Y�M-2�Չ:�0�~ ��N� ;\�~GhK��(�i�ն��IAl�'/���IvbmbH��r��譧*	#wf=�I����B �fX�*8B�hb�l��?'��&ğ΄&u�����\�x�w����߹d���vMT��C���2\)f���g�n�u�����A�xw�����MbN,L�[�k�����oΐ�=�4�Z�iYQ���:�P^jyJ����o*Ƙ�H�-����w#�Zj���QY���j�l&ڞ����K~�������;�+��R�p����_e��L\J�ՀP8�Ys�o����a&�����'�]B=,SH*��A�#e>ш��D@�߭~�ɲ(���kl1;�m1�c������v��&3�wV�_R뮪2���oI�ѭ��c�|%��)Z�`���Q�ՎC:������]�����Do2��=EHԗ��
��i�/��쫛��i������b�;��4ESb��	�z�
@��%��2I�S�+]sJ��G�_ ��)b�K�9@n�[����E�*�Ƹ�W�rs�z'���������3��M��p ��p+���:y�O�;�7whɫ��Ӗm�ؐ�"�+���������b"���B��p�<ˁL�.n��$������W�Q��nk$~�%!���z��̲O�)��8lx@�,�(���zgp��[��J�1�J@�SYe85Գ��U=���'����׍���C�X��5I11�p8X�����ԖE�������Ea��-�A�-���I��jg׺��/8z��z��6����w�
H.^z᜜U����T��$���\z`��O�řj���5�����\(N�	z)��79s����|�$�L�V�y<7�f�KKDe	r�������q��s8��\-���;vnHT%J�6�̀�|�0!#PˋX]L%�?�b��x�1���@��cI��{f�b̠k<K�}Y	�/�mkMM']l]�'Z^�Er��Z�� Z�O�X�x�X���b~��8C�!�<u1���ڛ~����ٿ�Z|����D�Zq�h(c=�F������U%��|��j�0Ky�xC��.6U��VE`i5����%���HT6�V§[��}H]$M�9nf'����-�5Ԫ��y�t?p����y��z�������ٽY�k��T�>�U���Si3!��sG���n�Y� �2Ǜ��Y�4�A�������LF�^fEĠNTڐZ�PoP��W2��_�YojGh�5a9� ��)�j��<�Rs���@j�0��C��R_tە������x>0Q#1���r��JR&��!Ә	��~�Z8|���IW%ؘ�ǵׯ�4y�>�7�B'�~	ʨt��\�4���b��n��<����⟜�0pIR��7&�dY����)3��?l�I�����P�=���/��\��4_HOZ^��ZQ���Gg�U�
H���
R�K Wֳ4��yW��o��� �sSA����!�4y=d*�!jSQ�>��C|�eqB�������H�5�rc���+�
�M�WVܿ&t����(�sI5���CF�Y��DT$�;G���3�1�O<���I�A%�H�td�0����M_�P�f�-1�[��,�;,�"���;%�Y�e���|�������3`cEն�%l1En�����E�z5���\��I'�ؓ\��#��ʤH�[@�1{!�J����cM^c��`]$k䒃]�fU�j��y�Uf��������݇_�2X�����xc��!T@��|F���&#$|���J���9n�IjrB�b��}I����[IoY�iVF��6.��n�g��1��^.�$���!�!F��+�� {�'2ըIx%7��� M�Rǫ���H�5��!�)���̗h��1�$tB�g�@v��A��TD��9
G���2�K�8��a�:�'6�C���n�Mk��f?�$�Y{�l!�p�2�6d���3�c��x���3�<ӎ�.�N$���c]LM�Z9� �F)G�IaY�2#+��}{��C�Z�,��H��#����Tv���%GŢ�xmb�}s4�F0��0��$���kNKz��ڥ� @՚���Jg��(x�*Z�����~\6]��Ķ�*O�j5��J������^N�W,�zZй,_�������k�ND�ؚ9N�@#��8u��,�=H�u��L��O
��n"!��:� ���:V1���[��/�!.E䌼���>�gY��T�q{��dGS��8b�cX��B��F���Dr�2TS	�e��Q�Ց���_���"�
<���Eݝ��=9�C���Q���I��T���x���&Vm.Q� ��<����o;Ķ_jY�lĐ?�f�d#�"e��2��-̌������I��%ʉW��� ����,3E��d�1��؞�"0�W=@�����l��5��F"3�2�a7�(\�,;©��
�u�pC��s�o�2'A�:Ʊk湒H����h�� R��\O��e������r�n碌��d�6u�F�H��8aKl z���"iY֢[DFuqC�4�apNcB��	�<{΀a�Y�T��6��0`�Bf�k�qn��%���7���T(�ć-��&���P�T�C�ܝ�N:2��i��R����e��$7�`���"+X�No;x�&bG�ŋ2�cgd��}Ћ�$�Fv[l`��MN?�ZU�2e������8��&���V�d�,.�-�vlu������RCGew�fe�Z.�(����S��t�}7���{��o�;��d���+)}��h�Rũo�%�5���ޮ�w,l:�>BB��w�,�e�T�߅�ƺ4",�x��L���P7X�W��9���h����Ą�7c'����'��ZrЩ�����4�Q���b��,����3��W7�0�C�Y�{n2��ͬ��v^\������T�GDO H,���HHQ���A�4mه����3�M�chz�X[��:�~�F�O#�N���u�Ff��2�2���Q�js$YA3��fH��xP$�(a��V�LޚA�R³(�MN}o:X�qYr��C�o�����p�B��&i:�Y�T�
����a>R�+�$>���`�͘]6O�����X���Ӝ:�_-A�撥f�y���p���ǋ��L���a��U `}�`%H�<E���'2�>��UΝ����Z�c<���Z��v�l2�CH$j]6(�Я �ZN*���S���aDjӈ�i%A��B��������w���ń
z�W�=�We
46s�K�RS��%�¥G\'zz�ڷ+��G�:%���L�_��N�yQ�1$�d#��>w-�<�0PM��vmf*��̭�=�$�$������no����I�Aͼ��_�ٜڤ(j��!���v���ai�q�v�G�tk+ǧ<ɲ?�+[��~MU�͋F;��!����Y�a@���� 5����n�^@���i����b'0�FZA&y{x=w��Uò~I7��B��>��A?�|����P��H�đ�fqB���TR�I3֗��92��9v7X��+�|K�K��oG��%�S��:Z�}�M )x���T�G��=�L��M]�|D��<�֒,Y���2�X9�"�08���lM"�c||�M����%t2��g],���Fi��u� �2Ύ�
0���=�c���� �|��/FY�XH&�B���"pL�,2`�;���Z$V�n8��wՁ�I�7/w9h���tƜG��Z�|���3c\��U�I�T����F��3M��"�2��P4Y�d-���ۗ�wG��|,�2�OG5Y�,_Tͧ�W\)�pv�(�P��Z��9�]�߭�\{�a��E�c�@����cꕯ�Z�*��* ����J�<��3�F�v���=�n<�R<e&S�'je��19��E�k�}ȓ���W�8�
�f��\�v'���U 4>��phVM"�z1h��PL[�ws.�\u�Ξ�ߒh�Y����֟�#O+��߳�n>{Jl�o���]��NX��u��{�<(K��;u?�.�
�Ƨ3��3����w{z_����k�l�G��q��\	��F3��oΠi��8�I�W��J8�@����Yo@"�w��4>�_F.'��3WF�^����#�Ds��W�6�Sa����]�(T�ń�0�|h&YO��ޥ��mxn��'�P[H�=(���wQXIt��.���<9U����{�+��2��5/l��W�Tdw!�B]�̇8��p�`3�GG*��w-V����!��Z�=ی~�,�t�A�2��PM�Ju�4B*�Yy]�p8��w�������ع͟���2?R$�*��U�qa������+� �F�t�V�{��W)֤��Z����͇H�{t�B�c�|B�e2r�?�4�R���?Aa��Z��t��z$P��ʱ2(Q�}H��U�P�`�n/ ��wG���֬,Qm��7����$��юLx���O�g�h��m�� Р��+����2��{B�x���
y�Sb'��)�/|;�R���C��s��v�~?������m�v =�a�
�ғ���q��b�7��]�(�-����I�]��N��8[��$F���T���z,��x���� ��*�ӊ�❝��o2�$��pF��]�;W��VQ�<&حN�Xs�J�B��S$��y=*ؠ}H�HR��>-^�h2Cf��|~A�>_N�(���4պ'��ޕK7��)������YI4�3�x� `L+�����T-g�`�Y�O�qb<���s=h����f�l�,*N�1٣N�H��<Ḁ��8��-�*�ҫH��s���&����͢��cv�����x7b�y�Z�
�VG�l�8k���[Ze�Ӫ�ӹ�Î%�r�~.��)����Dѝ6�d`XvUXj�@*ͣ�
5��U'�iu,��[ž����B�����s_U^ O�����~��9�\�����{5k�-v>>u��h �(�Ᏹ��5�L�фύݐ�@3=^{���J������|R���
F5���ۑZ�a�|X𙔵!b��5#m�#�nQ����j˲w�nj�&l6�|c��, ��P��C^�D@�"�b6���r(�hQ��;����ca�c�����Q[��lyΏ����]��;|�S�kq�zKm6i�f}�L��#�	Bo�A�G|Ő�-�ŎduW�\�}�X}CW|Zf��є}����b�!��D��}�qdv����T"[3��EB�p�d 2� ��	���dt��y=Ÿj��_�`��j9_�C��2=���2�\�q-a^��J�&��|<�P��d��X���q	^��P�J�4���K�&�wubc�we~�W��ǡ�ihT1��Z�L��6%k�P`�%�l�� �aI�Y�E������R��[�)���ו ث��d�&U�1PA�Yk��e����%�2&���B["��l�Dqd3���t�N6�O�F�-f�a���p�t��5��L;yD�i�����@.�4n�칀	d��l��K�\�5R��sC�H�ƣ���-Ʋla�
˰A W���yI���bo5&��'��N��+����J���!�x������İ�-ܧ.�Պ`]���ޒ�aL�`���
��;�-�@(n��w��㢢������~� mc���t<2�r)|��!�~}���rQ���Psb	Z��9/����6�%R�}��ZQE�_���JX��l�T�s�ͼ��%�0u��t������4�]�K�i
}ℑ��u��������3x����F�wv�|f8չ�X�m��dā!���0�)ۤl=-|F�L��J q���K��>;���������%�ttx:�d4f��J�\9�Ձw�-n�ЛD��yvzN^����~��zs��Z~�(#��O#�_&x�uN��"�v��a|-��Pܙ7��٢^WfG�m�Y�# ������,�-ŝh��	�:�cU)0�̎�����,�
�7�6���J�ֺ�%Q�_���˒(� ��-y*�-2r3_g[�`����s�k���!-�H�k�h$��9�������:���(`�ȷM��V���DFJP�[+�d��H�c ��kE��coP��Il��F5�����-!���l)Phk�&�F�/k+g3@��Φ�Sl|���&�0���<�g(����F��{�W�~Iۊ>1֭���N���^((�}���/�'OZ��,�{��-�o^Pj�xZQ(�j/�u��Z2%���I��7,Wr<-k}�Q�-"Gύ�~ޒ��OR~��g[��W8�3���V����@7G��ՠ�q�ة�M�e=��n�?�3I���`�F�������FO��4p^��o'�������.�<#QJu|�TW
b���(�=Zq�2�@Z&��@	�����KkCHBY��Lk�l-ɿ@0C�!��O�ݩ�&Q!��	�N0��mҏJc�id��Vzȼ+��[2a"�9x�����|)�P��
�����E���qB�?�33�"���x�	�>+�"�~`�AX7�"�w�Iu�Q�j}MZē���%I��/�P]X��\�C&jT�s�1��J�._ƫ�������3X��" VƯ�.�3��M�
���ѫ����G��$&g�T��v)��a�t7�Ɩh{�{���O��g����m1!U-������(��گ�kZ���)�Q/���}Cx0	�Mr� o�p��uZ�I1,���ؖ��[��L�Q�"�aNcqhs }&s>=r1��>�{�S¡��U� �b�h��mD�;ӕᘎ��e�����&�KJ�[��1;�_�qR����+��(�qf_��L��2�3����ӽ`�?�)��s3��)��N�>�k@��_�zӵ+_�`w*�.i�K�Q�����%�.ć��_N=�e4�9�IXji�f�s1q�%�w'�"0��g�!^�0�U�>�`C�f�������2���[W��.� �⯬�e�gJ����Z�����Y�)���J��>זS�ы�þ1�ԉ�����N6�$������W~@�+|Mnm���)SH�a���2�o� ��5W��dc-�'\ʢ�Jޘ6�Pm�j��]	e�F b;�c�O�B�>������>��ýjP�ն�@ހ���r�W�3���9�Z|���X;P��W�6[J�O�W-YJ� ��}�D�^9��% 0���~*ݗ��J�?Fd|�x;������|o����a3U����%l�g�0���ݠMB��t@&5fzn�@S@�l��y}sh~83*K�m�P�N/�*� ��[�����^�o���A�q1�e�B�ϥ����ꉖ��"P�
;�[/;
Iԙ�F��4#�ӫmo�^g����x���@C�J�AZ��JR�Tk�~�{��3P�fD쯭ŏȪ�1�~�+�s����]��N����5��J�Gu���@��+�/'����a�;��^;9���F	߆3�#<�30���ӿIh�:����	��Q�� ��B�1���P��x�q�4��V@\�6 �{�iJ���k�Z��d������	�
4���V>H. �*��[��f9%�6��^Q���-�M��Mq��N�g��i��i��I�4���`�U�>�وê��fV�@�ݒ�W�Do�����@��Hђ��@Q�+lD�Cѫ_���2)K	gY����~���x�z�D�F��o����������BV�n�f���a�Qź<p��*[z�����ʕ-^�[=\=�hl����9c�P�l���KS��
�1^	�x>��vϦ!_eJ@=��j�b�� D�EC�O�qz���\)��<�=a�j�]�M����-0����&	�T��E�z��m�"cF�$�,/���������^��^�
/:�!>����x�ˏ�ϗ��ZE��(\L$�V
%)��hy�T��
v�9��m��o�RD�g�9'�Ɇp)��@��'v�TyG�[儆�����k�LqI�^z�x�gU�TJ����&���(n��M��L�i��K��	�Ji��p% &k������i���z��z���Rv���W���Z����1��s�/OV�$D����|ɱ����W��j/�Ep��1?���@&����-���Sh�wraAճs�$��6�+�ĉX�(8\I������x�Q�R碦�8�D��,A�|��9a��]��9�4/�����`	�l�e�����b�����J�xR�>��]��3[q^�䘠-���/#�j*�b�����-wW����H�,�&O��W�i�mZM�ncy��}Q���}{#�V�C���n%"���bR��mj����R��B9�
}>�ŞI�}�ް�'�I$��F���(3�o�;���B�g�n��9��T23?�6񚪐�˱})����L��{3��s��$�K�4	�&�h���s$��T�n�i��Q:BaY��
\co�71LD3[^X��LO���R�P��Yr:���G��웋�D�8�svKr��^�Qy ��CWْ�5j�\P��$Q`,����_�R�n�U���餡�ÿR��,��u#��B˅���%�?���̐C�
T���4��]g��F�9j\z��-�E��`i�Ĺ�z]�w���_Y�r1�!�Rc�.�Y/��~��b6��Sk��.Id0§�������X�{w��P��� ͟�a�f��`ُ@A�vhx����q9x���Y�P���,Q�Ǚ�@�<��DM
��m����U�z��d�y��x���M �Ü�>���79`p��N���%��FH똷_��u79�|T,�Λ4�$����6�a��W�::�T�-�����$Z�ȷFj��[�Y����'ӗ�>R~ Y�d���?�9��{.�p���LM�	�،TW:U(�<)�����1r^k�d`�H՛�����]\���.;�*�ZxxF���,-�7�&f��Y���-��s��9�zQjZ������|��t�$>�VJPV�� kC���ד�3G	��,��Sh�`���f��w�Em�-0ǣ�*��C1�a�*4�H�����8\b��y$1r<��3�N@�D{�ʜ��;�7���X��p��0&�&�H烮_��8��?��������O�
G�t#}?��)qP}�,;�_p��Ÿ����[[�dF�*p�����3�~��%g�	��)��%W= ��v�'z���H�Bgw�\�`�p�BB1�g C�EU�{|���l/�efע�g�.��憡��#E�r��
��PK����H[2c�y� �tV�!"��7���޼��$5����uB�B�"~�m�rm\C6M���]���[isCt�����5u�;��=#�m772�BZ;��S,(5{���( ���g�q.-h'�
�I�bhK�+ev=���_�����'��=�J r��LjՁ�U��ްy%{�u?��8B��ą�N� �֩�O,g.��p!�Ǚ��m�:��^u2�RT3�Z����)�kٵ��M�(��zaEG�Z̔�<��"t<�"����3�/h�|���\
�OV�@7�ʥH�*R�2i��'��� 9����N�LKy`��Ņ����n��Q�ݟ��M(��ܘo�����H��$�*��y*��|�S���F��;��H�޺3R������Q��S��mb�놔&��6�����R��ZYe�������Ȟɲ�H��-����w�'�7M�����l �ȷ���W��M��y��(v�l����:%�`�����ތ״[3�u�u{��83ft��dU��C+�Wm�k�-,_#F/\�w���y�c��T\e0v>:1-6��1���r_ zSr��������P�}?�zh�9+KX+ٛ=�qh���pꊧ�-1�N��:����&d����絑fV�"�i=!��P���8�KǸ�w'	�(l�e��ٸ߱)H��9�'���9���:����giX���|p>	}�2������H�q���9�..;-_���ߞaJ#�St^�OX���Q��\��\a"H���zԱ�K��^\�������l�&H9�?H�ϼ{V0e�"�?8�;�9�|	�Ȕ0tB�WaA�+
:h���#ܨ6#M����:�G�pb�&D��Q��)�lY3���f�z:Fs�}<a��Ϸ�|t&�"`�N��h�3��x7v��ڝH���4?��\�@ M:�81�:^9�Ђ��>�U���Z�Kjt�׼a�l�(�>K���2��+��ʘ�خ���Ǡ�?%r$�ynND��g�&��  >�S	G]��1�N�[=����5�h�	���6S����\ގ��h٭Gfe/}����V���(�Q��)��"���Yz�&p��zd��F� �7o��$%�s��q���l���|�R�4^'�C]�����#��jt��7��B.n��-<V9ü�f�S:mz?�p6�خ�i!�^er>�'�v8�����x��_��>�^R�D-�y Yo��xD�a��!�js"�5DSE�vO�=�3�X�@�g����j�`T�(�i��	"���	�l�oq�bx r������|�dW�W
�,�{��\\x�\1}�]��QК+���h���ڋ������덱�yF-5YſdD���A�O�e���mq�]�0�Z%H��m�n(���~�j����+���:�8t�G���t�`�"G��H�U�V&���/�}�\3�l�!���?�߭599a�\b��X2F����k@���si��-��)�D+�x���IH��_ܹ
U��/������9��9����[��=	��+6Ep�p�d�Zq�����W.����������C�����c��Sx]�Щ��*t�!��C)�2avL�O��;~,c��ݫ#a�R0��E�H3f�X#1?�"N��
�v�2ܝ
�!
�J�s�j�B��]���I6��`1�z��Ǝ��2���&5�3H�,~�����,2��u8t:)��������a���s�,�q3"��-���̀�4��2��e�z�zw(�a�1�=���Oj��6[.E"'�]FD7߾_�Zr��dDt5���Ws�|T�@ʡ�����
 ���Lats�_LO�A��i��';��7��g\���:��N�rP.z��D��S0�J�<��d��~�fH�Ʒa����T�2�������������Qpulg�^V��8����T��z�) ʼY�?��.�݁�Z��O�/97W��Y�����f��[ի9���Y������H��C�ү�,�@���x}�5:�؞e���q��i0��Q����v�X���Iyw��P�)*,��n��0A��4�Ȝ�yE�u�)��c�J9�0��$�%]��[b��<�pI��t��tNn�ZiS~���q�L��|�R��~ϟR�����ty�0I�c�to�����h�۬v[�����o��,�4�{��u�/v�(�8�	���M-�����f��U��j�O�WB��Xd>*E2C�m�̔��.�W�$d�u���
�I\bʭ�&Ay�T��� z1\�2wL�t��YbEzkO��E~�+2?�������M	�N�K�]��󪬴��(�<��h#q���PV�s���=t/U�`|7Lyb����'���}�䊰��0��_�k:3p`�����g3&z�ג�X,g�8 ��a5n�]�`L��#�n�D޹�};�>�ǍEp ��坉{��3�I-4����D6$#&�W�0��2\qj�bf�\���e�`)��\�Llj�u),�A�u7ٴY��yŽ�����(	� %�z��	��\mj��ս��ڀ{1L&����y��gOPD��6c�^�S~	����*stׁ�-	�F_Z�{:w2xB��â��19#����Ȭ)�0k#�i�#����y��H+��b�:���K�X:�!�H�����)��4Z�tv^\=;k]8�����riN����	&�|��x���
�!�5]����,X0?XeK��>F�D�&��	iT���!�
B�+��t	{�IOJ,��Z�C�=�o�cc�����q{�ʣ�)#��Q���[�Ni ��5�XA����e+���[�qாLX�巿tM�MKz��j�cH�(4��F���ϐ[fY�L*�Ul�;p����WRC�;҃@3�q�Vj�r�yܳ@�ϙ5����](�����Ԯtj?`9�$�j��'<�8AC�be��ǖF�]���
Å��\�z�'��c 1�{;�$��^�Vc��\�꫌�X��-#ݫ[��/(�Y���EDPd�4R��$���2�P��#�c]�5[�{�U�o+��L��Et�tǃG]�����r֧��ʐ���I���636D����z'�,�Qi��ױ�9�W�D����QA���fy�O��'��nf�����<�Т��7�:������� g��+%P��"(3ȅ�&��ǩs~]�_uI��j��Qc eeac��5��͵�t וG�	�W�Y�$P�d�p��m)�C�,��w�ar3bB�2�-M�Oﾋ��k��!�`�� y#�|��JJ��E�>���S�-pE��G�B��*G� *�-�qGܣ�>E@L>2�R�9:[9���ռM�i+�9E���샄l��E�F�����5���瞼����y�벝�K�R΅�6;�^,�YK�[��(RT����ǂa߸�	��x�	��!_�ݮ���P���F}�/P/�jF�E�9��p횚$�!�(B���ρe?�U7ae�$�A1�F�hPd�#��B�C��������S8�q>aV���zGr�<_�:�8�AKq��s�RoB~?O���>X�l��2,�<Ab���A��n�埬\e�@{�?��U��m��l����6[��EA��b�A�_�S�Ģ��i��0���~��L�]
fn��ߝ�~��;1�`���Щ���lA��[ܐ	��7w�҇^��,5��!��POw�=�lU���"�?k��c���y���{��6!dfW���ƺh�c��2JK�^���m�m��^�{�f�W�]�ED����kr�+ʂ�[�܄�)��,An:�u�.�����m�K�r����m}~�%�=��^oV�E�z
de�=Ї�K�.V�88��Lh�v�+�9���?�%ں�e���%�{U�n/���<�1N3�ԅ=O�<�_��>1���ǲ�l��#c�ު��b��E�cO������MS�B�Z�ȮAb��:^�`�g����ծ�R����������%)o"��и�z���t� ��I�k:[��d��B�K��<���b����dd�7[=��*M�ҟG�[ L�z�nb#:�&|=�i�]~k�[�%�?��	~�LDG���ǚ��ŤE��Ԝ�܋^Y
A�_�kɳ����G�A�ɤN��[�= ;�Ҁ�����X7,0dl��rx�
)<�0eh�����FZ�Qٜ��6`:�IC���E�m�{6����%a� i���;�1��l��-Dd�zj�o�ҭ�cTzǕ*h<p �B��p�7"����ck�r��]o���'JV��t]�O�8+������q@ٳ� �e��H����;�M�iNX7�+�5�(�R�T�4`�MJRҸF�[�w� A-���3�F�-�!W�8�j�A̻���%x��[����FN�n ���� m�hr���ݓ�,�SՒ֊.���T
)T�#�P<��7%3�5��{���HǳV���M����v�X�R��+W���gAa��8X���l��K̛d����-K�3�y�i򊀁 ��Z)���I��ό���Oz�`|��˵�*H�B5]R�fM����~�Xݠ�w��ݠZ��X�w&��_��ɛ��%��j�8Z�\��G������l����#�B@�\9���Z౼�X�ړ1�Wd�=��xm�X�*�Wj�b��?�`��Nqs
ZJ��4���2+�ɍ-��Y9~2�w�`/�#=1��iQ��B��)�ܜ�0/�8i5nZ��T��-qhc;���ЎW�-~n�t�����������E���v��0'�pd��t�\�{Wtq�<�r��P��;Q�6E.�IR�Ҕ�&-�����ߺM�*LF��gF"��Z ��o&��W:����D6��|=�N_��kITwE>;q�P����1�r�RE�p�+ƫA>�b�딭��}�:m�F��)��Җ7ӗaW�ֽ`m��;��V�c����_�	p�{+HUa�	+��z��0y�s��8�0Y��n����׵�s׎���oA�N��1B�˓^���H�_��]/|������F_��m�ҳ#��Q��s�S��x)�	�&�P��1��)�[�R�^�l͔�Ӻ<�3���Q��x�H^:��)G�o�̟^�)��۵[mX��:��u,�b�5ZAd����}'2�W\��Ce^٦���;��[�I�����`Ԋ����g�ު ���K�O�_q0_g�,�D����`���`T4st�~��3���-.e�8"���"�ѥ�C��W���۳�039�)<x��!s|� U%�ttr��ƀx��}+L�IA���+�8)�A�"������؉4�>$3 O��&=?#�;ϧW+d����e�>���zm&f8׷ѥ ��x�^�͗�ѢI7U\���q��&+Mz	N,�U�%.T^��o����'T��-3{�_ݪ�b��@7�P7BtKċݾ@v�c�?�P�b�U,n�B`(�3�\��B\��5\?B���W0+�O�T�e!�������l7FfKk��#e�g%�T�a�?�nD�j�w��9{�܊��d��*��!~vA�������ɰ�ii������F2��m1�{���E�X�<��G|O�q��;j��t����#KW�����{��� chn}0-��ͤ��a��U�pS��F
*� ����#���7:'�Ր�r3��뵑��;B(�<z1�����L6�hYw_�`J^	��h�e���s����A\/L��d(���nBz��i�(�`)uz�ݻ\\&�{ "˩��$#ceK5��h��Y2%�̠�[[��=�6�� ~*X�@W���p�����r�Ռ����
6�瞤�v�����6W�ZH��_��k�Y��-)�]	�G�**s� ׳ܷ�J���Zݒ��si�ӅS(���^R�i'~�`��Ay�u�
��oF'QF*%z\m�Y�����S9UpC_����C���
8k,���,��e�0��?hTR�9˾&P�q5CZ��{������*�Z��F���3{hLEz�q�Z�Spf��.$g�=�[���b0ՇT-�܎����e2АQ��P~]�d�+eV(Z�GV�ŕ�Ƅ�Yg~ ���%h���&n�oV�f���U�/����OtjR��h���A�H���3W�5%j����������u�1�ȱ���`r�0[�"���0�
���'���eJs;�n�W��>�)`.l�A���[�`gd�4E�)R���禋����"^=����^խ
����?6���~����E�+^�7Cc�	�[0��C����H2�;�Jŕs�'[Vk���(�.	,���c�@���O�������	���x�
xT�4^��5�r�q׃�d����b@�/��Z!�^}P��y,��^���00f��jt�	~�{���=�HB s썾� 1N�sm�^(�������(9]FS���.� z�t��ƚG��Ex=�U�[o�!ۇ�Ȥ�&�?�gf�E�i����� ���K��''���qk'J�e'��{�G�?_��� ����r�v�)��}g�5'���Od��%.��tA6Y��R���0��yHX;�?��c�Yp��Y���^�v�.��h��;J��X*�ox�c�
H�S�0=/�+��Zb�y���u%��];�lM��X_c/�DoJu&U�7����2^�(�<G�U}rpev��T+�B�EK����߾�o�AE�=�u�}1ζ�㖧[�Hn�xM,7��Kp�:���33*�q�4����ե���nϛO�׸���O��v=�ޜ>,��8t�Nf.�ٕl�Q�VtX
���?:�Fu�<O�J�����j4�K���<�aS��ʀ�zz�B|��Q�!8Dk��ZV�������;�uiB{hYU������ ��s�����d(J�0@������0
���5s��,_�<�	1�b�=Ā<ٶ�J�+)^�Lu��\�H�������K*�f7n�e�H���j��/�%ſ�˃`��B�D_�c�K ���S�(�偱#iY+����kCH�^�	k+��<*E��\�m�"�b@�JCX�)	"������|e�ϗ�.'���x�E�QFV&D��	�ZW�����J� s���H(U�����S�Z�Ӛ�]�����c��.Md&���o�(�A�!��p�;P�������ǚ�`��*���;�Rh�;+��Fh��ueO�7�E��En��uץu�:E��z���i��R6����Sё���S�KbёF�NE��ܳ|�2L2�W&#T���PX�{]����
l��e�2|���p����p���`̣�Z-�S��c�5/Y&�O��>� TZs�t�c�7}#����"�Wk^�,�����5�����f���viFC걗�
��E�����TM��$73�eT�l�bp�����k�9*�*nw�z��y�I�:Ƅ#'�erܫ�(r�Q�N��#� ;���oK&�
�l���$��r��p�ut��$tn��+��Q��`Q`�����}G$�"[Y��5�����6�lt�����.�%g<U���O)'�����0y�h���6��XlR(��p���ٮn �XLX�3XL������AL[f���
[%d���Ad_�LF߲� ��F�Z+[y7f��p���Xe@��{�ƺ�Ap\�)1(dP
)�̳h.:��(jk�����X����l�yp���A�n�^"V���bP�(�����C�� �J�:���c�C�R"�.��<OY�<��e�4��<�1�P��${����!��p�#��W�|a=D�u3��m�A�WA��X�67���L�?��Lݔ۫1�G���g��NG��Z����9��Q�rޥ����X��������M��[����;������r�U�k�h�V+以��w��娽&�����r�3���y2�q0��3e�k&3�u_O��"y�,��(k�v�s0~o�"�H�~^D0ԇh�&��M�y
���6p�sŴ	��0�� ;��[>V�M�=�U������RZ��V�,ִ�fK���-�J��n� G�Y���]
O��d�3H��dm�C(�ii����C�X��͇�_�;�#��y�WQ��|5�*M=S��e&��M�q��+��'�|?�����8�!57fe��G)>���b��lj�����!��$)��������_��[�Z`�_aڕy�	�uQat)�ҳ�4�g�a�b�3H0�em�Q��.�М�^��u��d�����p��胃��أ�����!>��F&��1)�|��"�@t�Ò��-i� Ⳳ�R�+�:V��f��X��{ṍ>�b]%^�EM{o��B����[�ԌS� �y[�*Ed�F����}z9�fR�j�y��9����Ɂ�WߣY���V>�?���h����̰��_W#��7U���RU���9-5C,=I�p��[-���
t�bjQ�/�f��[�Ӛ̨u���\�7;���WW���5��l�#��#0i�q8�=����]�q��䤅:7 �%%1O��z&&X�����8b���A\�ú�	x�F��h���G$�Y���_�`�	�M��`��H"ތ�<�6��#.O�O�"�t`�wR�s$��Q�R	��擪�FY�Gx�e��!0"������j7�	t��K�ht>9��cr2��ae��E��@W�y�y��S~��0��iN�ߒ����=a}�f0ͯ����u�(�}+��@�O���I�M�J\�)EHW � E��y��v�i�M��$��jW�0H�0A�,"����IA����aQ���ݠ �z�n*�� ���Z���H�{W��i�:kW��kN��Hm�kz�>�c�;���l{l+�+�oHڽx��C��<@�Q���U4�{*�.��@�as�>���%�nP�h��l�[L��"�\�ð��4sC0�؄\O�)����m���!<���e��I8,�c�H�n?a��>�!"L�*����?#tp��J���kwњ:x�-�Y�W� ����{���a���4Ib��c/��Y��cH���X�z7����5o�,"�n�;�$�J��G����FjmkΡs�����Ε�yVx�E���45B�R>o��k��)m��bj�:�PZ��b�c�>�0���8��7_jwKA$&R�Sc��J�&b���C���c����0��d}�P8��r�@?.�����`>D��J���9,L�����M�GZ?�U�����O]Q���y���lo�}��*�=���4�#>$Q]��]-�3r���w���췵d{�TQiV��a���z�?\�]��E�}�^�}#]"�O�=,�O,#B�؎X̓���Z�
����W��gr�-Б~'M�͏a��<�q��0�l��|i.��(R '|�)ݎ��J��ʘ�&���]��~A�l�X.W�[%��3Ё[ok�  �㵅S\��Q�w��Ŗ|/���!����XJ
�{�@Q���QQ�f�%��U�=�PR�o]榀��
̷����Zhӆ���C	�Dv�Q�u��k�Ɂf�D̉g��W�a�2��ѥj��t����w���Ag�ə
g��-y�o"�� i��lp~4�~#���)OMne���`G����o�f������ٟ���N�[�8��IyQÑ� hr\������b�m�{;��̉��7��ظt���g��=C���o��G������%�C�:Z�{?���� i�׺�Yi�!)2
3꺦��d"O'���|�q����W�%&ɋ����
�R~R�5��h�����]��]u>���IP��P��r�n�gI�K���T~)n	��A�SE����=b�{?8��P^n��H�]a�u��&��W8&�jK��4��e��� G�J��_��K{�j!S�SG�2'��D�G�����+��	���X��)
�$\nO�u�65{�3�BMb��@|�z��B�H>��f@E΍G���\)�7(���Uܩ�n��6�$~F��������D�T��!�%|בH:���+<B�������$����[�z����8`�D��`w�4j�40U?�<ۚ�o�V$���gm���q*ɰ:N�҄�1��.��]���I��@c[�q��LSt�
dW��a=$YمGX�Ӿ!?+�)��;04Q`���1wo��`�$�* �8@4�BL<|������R���D�枃훯������r[�a� ��>_�34a��[�t��Y�+��U�	E�2���hE��&4Ă	�n9�QĴ����u���s�x�����LP ��p��ߡ���M��b�-��G����ü�����������%��4mӊg+ݬj������[U��?���t��S�t9��4�sE+�څ���"���h�䴟��$&�nl:��}j�v��;��u�m�)�HV�z�x���SD(N�5��������������QJ2K��!��?.s�k|O�.����9i�S�<� "n"aJ�'�&i�s��]d��H�9Ds�)�:qd�#�	�5�N�(����\C���o{�:]f���g��]9u'0���E����&��I�QC�h�z�mֽ��*��v�R�"~���ѷC�p�z� m�!�?���<z��� <��@�?�P���$p-����u�D���z�/��z�!cJw%�H�"�����m�D�z�~A�Q��u�Y|�ukQ1�8ϕ�8�XcO�a�u'ogi��jN�䌮ڗTq���/X����1Luws4E��xfΟ$�Kp/\>���?Ϻ\�	���'t��$;pB�R�R�8���1��E���*�H@ǔ[/\I`8���ϫ@����]�	�Bm�Q60J�1������EQ���#�K���>,2j!�Ý���9w2Oa�qO�zZe����)P�7�<��h)3�ea���`ӯVV�92J�-�|e�u��i:A��6Au��G�I�P`��ϝ���Ҧ��wkM,���P����碚! �2+ķ�N��j�l4f��, ���~7%�uY
�]J_k�g�.��Ҋ�e$Iq��s�T��*����s�.��7��W9)vU�3�H�(�ޙe�a�P����X&���߇�m� ����N�0*�Gb��O�.��;�����s�30�0�W�P(5-Gf����A�R���kɶ��P �J|(���Ma���Uͻ#i0Ã5LG�62�	d���/��]	q9	�����67�O�nXG�A5ى� �����fT�yu�^Z�����QXP�����:$^NK8�:leĩ��)[��ę�ƀ"�R!�w�V9���D�ble���\�'�T�EG'gIbf�7������zqgY��都��)���ބt�_H��c�%uf�Z��7�7�'���gV������1�܁?�C�k�u�g��s��� ><:C�)��Cx�lz��>��f�Q"wN�c���Gob\3��3�S�m�K�=����� kɿl����a���	. Q$`��W�#J���f\���,ց�F������o�~��_uc�F���!d�f��_X-^O���z(`Ul����,�2x�
�kY�qk�J|G��.�msS�M��/\^W�t��p3<��B�� \LU���WM���VMu	�L��w�9��r�lm�*R��?�\�p�Μ���9���H��������їW;ճ��u�q)��;J��@��f������E0��ˮ�ɡy���c3s`C�s�\�1?���t[)�0�S�L6��V�J��d�a���*��(������	�uv�=�_ )�7�7�6У]�	��8�b\E򂽐����5s)+�U�k��j!�ZwB&^���^M�;��A�)����.ݡ��<;���+L��Ƶ���t[�h��2Kx�� ��3�uU�Q��T'�;�Qr+�+�1���
��`�iȏ,�2��Tmɚ�c"����/B�,=���1"���ې����ŷa�����.�T3��400ȕ�k���^&�v��B�!��v ��ܿZ�%:�y����1�s>�M��ڻq;b�G?��A{�-��2��Տ���q*u'����҈�u_+�q�
R�,=nZ�\r4�8��sF��˳s|y��e{��\�,�p��X�XÅO����$��&��� ##���H�����˄"�[���%#�z`VL��#�p, !VKGJ�1��߈%H�g���4���D���n���Aɱ��x*R%2���!��Y]/誸�l^jP�wl��" �+�F�t��s_^+a4;��w�_#x�%��5�L����P���+&��7�V�(v�aMޗ��_Lc��#Bi)U�'·�71���/��X|������lRC}}�J��5ǇT7.��L��GAl�����Ƭ�9�QӞ�f
�zhJ��$���L;H��jG�q�>���|���RG ?�oH5���.(>0r�_�>���op�PW>̱?."̋=�{�����=1�����D�2���&���7T	I�	�;����
j4\�3c|�j_��e��*˝I��~8�n'a4b*��.-�3o�)`~Q�����B�|����7�xg�ګj8=�7�*gM���%̷c����=�5J(��0v�6�Dwe��j�8qzʦR{�k�H��ۊ%e�p��^Hz3�!k�%`�3��[r�Jv���^L�(5R�u��?�?�cmlX���)ݻtyu���1�F�4:�<�T�H����X�N����Bc6�[���>�q������!>��.�E���ξ�3��ٽ������s���3�w��������[��H�GE��!��0�4X�1��KJ�Q�+���AY`�`jQ���t�W9����5g0�C4Nb��}�I�cK>�j� �Tֳjb������l��$����p�]U�^�6G7ţ��g�آ�)��nfJ:��ޢ!'��w���]K�F|`��� �`9�9�<����H�[� >����oKC��Y��
ׯ�Ŷ�O9��q&��������u}�D6]����7��:�n�v%z�ga��J ����~_HƐ��9�����N��(??3�a�*�:O&�1Uzѷ�>LRd�W��Y�B~=��W�B�^�ЪE����]3�y>A��JQ�i���Ș�ļ�R��x��Y�Θ�����zЀ�qr��I�ƱLi*�S��(���r�wGR�N-�X�H���z�o��hT�:3�k��#�'3K��B �G�o0%lԒI[��a�.�>�^�g? ��4Y�tv/�z�V!/ m�`�A��Ң���(��Cy+���E�}2�oZ�L�v���6FJ6�M"�vx+a0U�D$;���=�)&�i0>f�lH�VU��;��juf�4û���gg�hE��7�N�}Q��rʏ�N%= dQyg�b�S鹐��{d10V?�W�`�w��)ո�F��*-�a�HA?�|'R�JZ5�1�d�g_fsޥ¹[�������e�0����c�6��*Ñ��\��8��7ڟ��<�p,	]�Z�NHwjR�k��'}������,�m���\Ӕ�h����a��VZo�~>r��F��O�>�nq��ab��dm�8A�6�lR��O��b�B�ɴC��Y}��t�*[��� �A2H���N�>��k����xo���������H�4_���]��B������'�9T�esXG�L2]�5v����7V��|�_��gi�=dέٱ@쌡z�2ΙvRYi ����-�|'�z{Xal�n	p�'T?�py�ł>���Y����g-u i6�W�e���D���f��SVY^��f�5�E��Hc��p2�S�f�ڿU��F)RBHS���*Or�;{�e�D���n���� ��M*�EZ⤂�56N��u�+8�ή9�x`�:4+�OyL{f-�W�&x +���Z��rE��M��a�E��@-���:��7d1�Vͦ>�`4<�$��3�`�V�˸g��?\j��gSgI���������"-���OMoٌ(��Q�n�����?#���|vC��ܕ\��2i��[��y�z��<9�qP3�����c��8���یO���e�&��/�.F�wl�DNm�B�x5����]������sF`�C�<��*��$��X���?y �~g%��w�:�@]��eN+��.z�ɒ~~,�<b����4�����Y��N��(]��Ƹ�Ֆ� ���1(�J%N�Ğ�q�Ǐ��ُHiW8���*[�?ċ�����	k�?,4��t�8HTֺjZ-w܀7V���@V�L��:w�p�+� ����j�N��3���WO��󹗁��ނD�������d�]Ã3�lK�*d��+��u��FPG�^����3���ؠ�(��݌=z�T{��	\�Y~z��o\��,)U������sG淿	��vO�y-oO#cR��D)�cBlQ�E{������t�WMk}M~t�W��-L?�L��D�PpRۘ7��?����#��#2S]�\��DR��M����8����ښp���;�����-���K�D�կZ�Dizg��1d��$��{Lp�$���Zs�Y���|��a�q�Ǚ�r��bl��;M�_�1�5�5�����Ɗ�x\�J�8���D���y1��̼��й���3|-oL�n�"��3h@��L����y4uˑ��6���@�>["zU� 
JH�<R�(/2C�&Ί���m��B���L,4�i��ٌ�H�
| �13��a����NMP�@�4CP�F��Rv��|9��Hw�clQ��׊k��>�<ovb������;f��&:V�ꅂty!&��Ya5�'fH�5����c1U��G!�G�W���
��#O�E�G����_�Um��َ��,:=i i�&շ��TsƃnC�7�0�[�.\:�������
�b��ty�l,k:����$;�p�Q���}��(}1�δꁇ>f!����-Uw������( �=$�4!�\����E��(������K<^�]�=�n��[xY�z�|B�4ԭ-D�!����
�����w*���Δ�������B2��-]���$&^d�`�v�-�k>�3c��f�<D�Y�aX���o��Q�Ȱ�%�N�C�\xL�f��V�6��E��FւU��a�lw}J�_\{�b��c~nVʝ3Ap��kK.>�Eߣ�7��DC��=_ӣ��7�1w����yVi��$J��f�&+����r�y�� J�R�n��Dša�7��w�.��R�M��+yg%R����fSlgu�x�},���]�T��ᰢ�������(/p׺�8-��+ [i��k�y/�N����Z�n��.L7&Ι2�&�T2��=������ߌ@����q?!��&��)�>�g�W��0�,��X'�_�֜	�	ٺ���@�;���CG��	���G9&���@M��P�����I�8}L��Lm�"��=W��RB��5/&A3�M��1V�}?u�{���Ra����b���!g"�4C�oþշ~S��`�g�w�D�����pNO\�{y6B���{�J��^M[K�A˵!ű�%�_��i�Q�H-16>$�>�k��p�M�c܀��Y)����BV�K.|@�V`����#y����O�˄F�y�Du�4y~�'j��'{�6|n�%Y� bWt>��V�bk���w\_�6������tl`��빈��y|��ً�;�6�Joˏ�v��bE->�קŻ��u1ָo.���yA��%%��.Kk�J��Lw*�hN����ݩ�h=7>-F���CA��w����T�"��l���&)y橧��zm�`�;��S3����-���v)n:X��ݣ���k���^�j��_�So6�8�n�"?S<t�X�ZR�� � ʤ\:!8�7��ަ����%�R)��ҴN��fy�Ts��H�gu.��N�Q*�:��$�NQl�4SUB�\�~�܋��������7s�B���7�+y)�y3�)�o�s�/��\��1{q^һ^�6�����h)�RRw���83�$5��K�V���t�4��rrT+���������5����lJ�	�g�&��~�7���t�X� ��c]�3w���))Lo2�#��r�0�?A���#7v��P胂g������j)��h1���R/,��Ю��������P�t!�����å4�3ڵ��rgz��>��	�ǐBJȶM����}zԗ!+������Ƹ	��G	�
�L�
�%G�Ӗ����b�Rz���Z�E0�g6r�B�g��V�j-�/3P6�.d��P	� ��g�?�O� OG�
�-C�x�3ri�]'~����DRT ��1q����v��0��f���p�t�.����p�z 9/��<��[�zӁ���B8~T�}�;�^Ce]X�+�͂�8d�7�}���O��C�*���S��ƚ.j4�ûQ���k9��k{�絚�5����v��;�j���*aJ�^�K�4�E@�2m�B�(�fM��"��v+�WE6@���QPWk�!C.Z��"OЫ4X}��A,D�&���rI���]H+��nbԡ��r�L=�β2V�3��.QX��E=
��U~�6��G�&.�w�9�x�yV��V|��o~�:��e@ʖ}��	�"<i���HvOa)��m�B�ί@�-L��m��in��+Ca�jή�ޟ�`��TN�J�9�Xˋ���`{���.c�w�N3�j���wA�<�����U�
�y��#�v��Pm����ax'��}��T��3�~tĠ_�T�3�N\��(߅~	hȱsz��_<	�mƋ�u��N�����9��Q����_9/���\i~�_\�D�������Zqf�7�i7���_����i�q[�%�.d�@;|&�ӵ��g�pB��8��qG���k���x����3���s�Hys��/k�M�INw#�È&h�Vls�f�� ���6Yk�+�H6@ѻ��Eq����Β���vV�_��P �#�U�VZ�b�Nv ��J"�d++���1}��A?��xzRU�Z��3����W��PS}Zy	Ne#Xm�h����Eo��Q�g�z��������5 [�5�`��<�����]�:.��-l��^ـ����G� ,Q;9y���e���UM� ܕ��ðRvл��z>HRi�ƨ;O��)}���84�q,��cnzS�f�EP�e��q�g�;� �c[�T���b]N�f���kOA����n���kAɸ2	O��E�~���g��.�f���	�Zؒ|6���{�d��:����wJ:/�B�_Q���/�
���{4�)�@:H���� ]< ċ���Sĉ,?���`���W2�:1(:�#(�"4Z�U��!�*����I�$%��pw��V%;�04@Q�(�E����u=~�g��#�����(\�4�#�����Ьvvj���д��5������RN`��x����@���j5�+M�z�n���S�d�Mc�X���wtO��R������a���>����!��r�c�S���Q�瑼:�����9�ǔ�ٕ(��kϥ��u��Sڡ�Zgc�:G��UeY+εh_
��V�M$��R���L:�	�8�;^�^dk3��1�K�[4���({.c�'�q�u��*��_���y�����C��,*��@�j}�d��yɥ$d��]w�3W��Z�6u�>:�gBVc��M�ػ{�c��|*1����~ĮD^b�'m���������yS�h��{�����i��ًyA׮W:5�!� ��C�zUZrm
�PAݝ��HoN��eZ�������k���B�� ��8׽m_�k��FX��,}�]cz�%O�n�!���|�rqy���[���jö����+3b[�؞�q͙ÀC�pv?�:��ۯ���C��d���xD^F��*)&��;�n�(�E�T	����S� ��P��h�ݜ/�3߅j��|N�1a|���5�њ�x>�k�U�w�KoK��qU�;��4�땲XuwU H������z����y�G~�j�T��V2�҆C�I"�d��Cpca2��km�{��K�����i��ԫu��E��䋢��Q�=��k���\�l1Ҟ��+Gq������1�<����*�C~�z��d�2s��"Z0�X&Dr��H%�4���:%Lu����dN�#�׿���0��$��_�W~ط&S��, �^J�]�9���:"ժ�"�cfG��Ѽ�>sZ�r�W���j���Vp~[L���~h}���in�jےNb�R�(�!C�N�ѳ����<��(��~�������5=�$z�D���yGOے{RS�Q[n�vU@�U�.<;E2:YQ���:[�w��Iu3wr��G��BhrvzܹQJ��^'j��h`x�Y�;��d��r�	xelu?����r���({�F����h��O��'�!��O^�=�j�2ء�6�_��(��W�,���lH�/�EZ���HK�f�)�!�㐙!�.���#"0-6a���+X[�!$S��e�T5 Q��"���[$�NJ�¡��WE��,�2IV5�A��ox�=䂧 ����kM���s�a	�Ve4��:>�<���1m0l�� ����z[�(�Ε 6������,^�"��0fw*Vtv��Jl~���NߧY�&��(�?2�`������u����靥p��\yYxHD F�6g�1H^�{恋~s�.��$�#��a�d���f�8��di}u"2�������\:M�
]��&��ңva���o���S�~��������S}��&9���`1�*o��غ�nA��z�+mt���D呞W�0ٻ�73^=TD��=E��bu�I�6�(�i��j�Ϲ��t\4jC���1l��APX��5����x�D�W��|�,����<q6E|�R����\��D{�K;�ͭi9A�m�[�z#uۖ�*��zqdZE����e Te,pZ4���̉��ȹ��&���	
�(<��g��C2I�����T�����"��	/BC*� �^��'Ȳ�����"9��A2�y�<�����Xl���jH�"d�魜��)��Z����������l=*��_�
u�J��09��:h)�<v�om\�4��u WM]T+��!!^���;f=ٜ�X�6g��$E=�n����\��ʟ%H�\�[�'�}h�^�f��0ہ|N�vo�y�S��eH�IZ.%���Jv����P�Pi�N�����B��w�BGx����w�mA��]��y��:�\�L*��9+R��V�������3�U/�>�%���a�q�27w�q.mp��/��VU,鷁Sܭ7#E2����B�s)g!�l]/�~�-O�b����cٌ1G\�M�ҫރZ����6���T�	N*N�ӗ������`{:܅�^g�9j.��t�!c�>C���|�߯�q_e�3��Vb�;t�E�~��?�43����z�T����6�6�s�н	�K�13��"��p�x�^�h���з��"E�Z+z�+Y!��n/�֜:�9�,��J��, 
x���@�� �t��Mʲ�b¬�`���q�Pv�%���N=�_+ -������N�5�9�H��I�w��ݺ��ER��:�����<o^^qK�wGo����t�Ր�mhrX�'��M�+���/Ųjyi��Q)j?ƽ��G�5,��&o@-�+9���D�$���ģ�G^����9�MPT���}ɽӕ?Sϸ�8�M$H_^|�&���E�r9��Z\5ٱ�̈́`��#f����2�r0��t�u�\'���;_,�:�����ct(4C�A|��[���'�*E��Ԛ�}�a� �OK_��j��SI��`)�mh���y�`�(e��F���ǋeE�I�#�=i
.��~D�&�)���`~��aǮ�EA]���`�~�,��F���B��r̛m����ӣz���,Z��1��E�b����/�vh���$	sV��P�۸�k_Ʃ��<��I���}W��: 8��G������3�g�/)ʩ���T�?n!N�F��r�R�@&1��<�`�.�c���C�1����+2UΚ��B�S��h�� �.�.ZaB�;T��>L�%��Ib����Va)�0 �A�a�4�@Q<E��;ܨ��6$����/�0oRs���)f�ZZ��b�ݣ�f6�P��L�?cbߔw�WQ�t�8.�+��-Ϸ�����N��`�Ɏk�����[��d�<�OY�3%�}f�]��&�{GARDz)�V�l�:G��4.�l���0
uƏ�;~Y���8,�~I*��G��H�h�4�|9ax�"�?���^Z<иX��a)E��dʽt��<a�D�(�d:���j�0i$��\R���lT�����0�?�i��]�o����^s�/L9�$N+$�Ͷj������S��HOw;�{ �auK}�"��F����|��k�p���i�FF��F�v7��m�/U���?��I��ܥ���`�j<��@I�w�6x�
��-���I��e������{�ñ$B�f9+�,��7��N�mO�������D�sl���6�h��x"��V#̡2Hi�^✢#�|`E(��w> ӝ6�œE_�)q��V.(�QCb��f�i�i�Ձ!���5v4Tq�҄�ŝmD3hh@n�_ݚA�\>�>i^ �����ɦ���ޔ���i��s��t�vu7	=ϕ�H�>O�6qO�
}���?���os�I@�P0xD�㦳��?'Q�L���lv�g���P&��+A�!UɆ��	cR|�H��n�=��a���3�>G��½P��~y�0T��;����"B�]Fe�2~LW����i*8	�1)j�7�­�B(�L�C�����X�
$T�*Z�_�4�&�$�Y'��	$H���cc��.eB�e�'F �:�z�/����E�n�
�,6��iI�R�FUާ�����0�)�i�6�<�P�7@����N���e[~��L���en��j^OA�u�k��ɳ�{�rV�8���p��Cu�"ɹn��|Gz�f��^o����Xp�v���pE6P�B�$.�CL���9a_���s{W��oIS��S(�B��x]�5����.*KV:ȁ&�΄�l���<ō��]�,* 6���#�Mۦ�o�l0_�
���|���ZܝDrB�}4EH��٬�#8���HH��t�5*�/�����N��Z���+.+�2��k��tz�'�m@��!a(���V�d��}��eދRSbR� �6��Eǽ���_�[B�k�[��d��-���D:�!-���w�G��o�#O�+L�ȳ<��K���H����	���Ś4�X��K����3�U���2���' Uk�K%��񞨋�ov#��B��>�0���k.�]����|c�L0E�/� ��I���(���=�yn>,!TL�?O�G;�.����:��4 2�{�>T�9�t��BK�:�ރ��X�����j����4z�(��kV8X�c�@�;_�¸�?<������	4H��%W��z�ו8C�u�7/J�t�N����H�J�Ԡ���T�u�1y��͗�+��ٓo��:�ӵş=���TPB�w{x.�Ƃ^��i�#�M�RalE�w�;��'+!�Hu�G���m~o��ڍ�|��:ƤlkF��!�b�f���y�3�70i�W���g�&H.��lO�{��PصP�y=?�M�^��>�d�m�{6�c:0�Y�%r�|���	��d@�l������jo=Y�YG[�B�~f��x�Y!��F>#����y�wjqi}�+ ���\��������W�����U*�G@ͫ��v�U���0^���9:�[(o���`��=1�����d%M�u_ti6n��~�и��ލ)�yX?��e���xx��[6�:Qsİ����q2�^'�������I�s�Fz�ly��<���6`�ˤ�#�E%��cA�v����OT%e-+5�u�w&��à�7�1 ß7�~���M=��+�ا�7�� ��H����L��∩���g0D��
�`�x'�# �B��Κ�hZn�
�`"%M0�݄������o����U	N�q�__҅O���w����=t�פ�:#�!2c����TU�&��$`<�Y�L�6+]��]���;�Q�TM*����K�dA�r��Xnۯ�a�T|M����0�:C��ٙ��wm�BV,���\P��2���A* �yg�&��|X�Y�^(i��8�BA~c�i2��(@JE���>B.�SJ�i=���S��;�7�.��}�P���g�������ّh�e�G�Y=Ь*��Y�����*Wq���"�7���#�8�Z�rG�n�ey���so��7kk�`#mp�h �+�}@lB�7�8\��h��śjF����G�gf�]eq��7���3rP������}%ts��y�����\�(�άXD!�5}�vI_}9�$���N� W�c���8`�,{�U#�h���,h��sɠ=��v%a�L�����9� &��P�hh�3����1+!�sD���7���������܂�����pZQ�|��TN�F�#V�e��6>�! �%�a�a�~��gN�{}�o�i��.F��g�La�b�B���{ўX�0j��)�ᗁ�������~��۲�
�;���}9��G(�_��d��ܘI���e����]�	�ѐe7	檴��)i������2������J�h
`�e,��FU���L�]���l��Zo�H=|"�R���D�#�t��Ѡ��������o����
3����+�(f߭���`�jt��C�Ap�կ��_�5�kX�J���e1L	���fk`�2��IH7<��X���<2��7��LY���<
f�q��Qت�A�zB` �W���=ʁ�=�q\��T�,���#�ʪ�T�Y8Fh��:�� ���0Ay�\Q�O����5C��_� �����(T��Hυ(R1Y��Kg���q/��c��ǳQ�;~�y=�d�	J��Th̊���G�*9����9B�����%�f�jX6�ಖ~�p�:�o3S00,��	��ZS�kc� 0V#�< �@�su���w�J��'�#���_"�/������Ͼ�~P]O�[�>geL/��G���bs���$+b�k��u-�ō"�c�n�UH+�q����zF~�F�7� ䷠b��bIc(P���&�+�ck�B/X+)�u!�!�Xk2`�SW��EM91z3 �:�\���k����h�v.-R'���� k�@�r�������g�n���
n�p����R2����B��	&��j�_Nxȿ��o�诰�4�

�]8��a��0YW�4���1�w��_�Zr��7d�cp�S��x�AC#����޵�V�{ot�r��$>�m*����x]4%�&��TM%��45|Y~�o��R�����;�,��kr��c�&*<��G�Ōo�i��+���`�{ G�WϳÁ,`k~G<a;�.��s�����W�e��{d5��-+�7ǃÔ�h����V�C��+�CF��+#��L2�3\6�s�J��CsG�.$�*8���3�y�D�^��.�[�E�����6�z@�z��-}�Ğ��ܶ!=q��r��ɞVՓ[<�M���3t�M�%������1�}���p������X�U	m�*�V�d=�z��|<���܊HG�G
~����v��p�3�kM���O�襥~�� b�ao@*�/	�Ie�6�JS^���[��|��f1Z����:��7"|xT�z\�w~��+�/y)V���:���]#]��'�Z�F�U��4�Y����� <��Q�k���yǉ��Ļ�� F�!�d�[�e�)��<�n�!{0�?Z���������ۙ�ϝ��17n����NF�<��M'�/a���ٻ�bt��?�7��]�ŐZ�XSᓍ�4�A~|����dT�
���)`�)�]�c���Ȁl�mĮ�k�Q���RH}�)�r_�sA��SS033�6������WV�:5$���e��m
�tU�t/�"M?�n�I����s��@Z�ǣ}�=4��)�cN�^�'zi�ڨ��:A.�۠�O�����1��K'�ƟjI�؋��@.ըI7�}���-%+(y����7eL� ���,�0�����8�(�A�:x�+b1�,�o��U���I�t��k�a���Jl�0�	Sҏ<b�E��l����ɿ�E�)`��){�?%��q�+n�������"�MA���2��� 7��W����x�o-�+�o�*3�����aK���Y���,�g���6�`�I�+O���,=A_)�]����4��-����4�I�]��d\�������&:|�*	u>�j�@7׎��N�^���t�B��)���{���w(#�m1	�KҊۃl�
�T�^�������
͢�C#}Ҙ?P�I��9��ѓs�~�w-�`�b���d��>᱄����r���LDd^)��3�Ԡ�u}:\[n�@c~K�Kt���JK� !5��pOE;���u1�S��P����Q��^�!���
��v�-6���( �/M�B�dS�/�wW�e�����ȍ�e(Ȍ�CUD�m��kQ�vUs�����5��[��r~9�W=5%*�-��w����4��6�x6�����1ː�}���/\}�	�0T�2`i���9��NA ���Ԃ�v;���;��4��g)�Y�tP+kv��V_������3K�[�ȍm��ԫ�����\|Id���r��[tp>u���;\�r�ȽQw3q�zM9"` ��~`���n|l���4\Q·�!�(o��*�_%�K�+gw�����;*�ñWl4�bW`  n}�:#R��@d�N%�ߧj���%m�M�x�M}G�e0���'��Y�Z�"��;�2���~�I�����
��wkf/{Oo`p�'��M�	�Do(���ש֚���L|ެ{6K9h�Σ�)$���׷_��#���W��M�l�ˏ���̦�͍�ȗ�jo�]o}�Lۄ|N]�w���A�@Z��c����M8iЅY\��������Vl<y
�E�Ko�dD=���(v �D��h�Ȧ�pؘ����}����s��KpFZJ��ݯ�/-��-�[<�,�j�H���u�����XM�/�ip�8��_
�f��Axr?�ƙ���nL��(��uR&5^�m�zoc"7��'ԏ�]��;8@*<G���Y�U4 ah��f�d�f`dٙi}��}s�n~������	2��
҅˹q���V�
�K�lg��)��������A4�����p19#�]JjɊ�h]&�������~��}���9 ��VdBX��<�R[�V}sa��U&�7��0F~Q�3A�!Z�m"�c,���m��g`�d2�H�InDH3���մ��MLb4����N)(��T�Ϻ�@��y>�̪�_�.F�F�FxD�S0�	������ۤX����~�a�n�rt�J�)�����9�Ow�'�<�=9,�2c,��w�-��Ĉ;5�PD3!7U�;��R��)����+�^S"��i;��;�T#[�;/I��MS�������Y��f��l�۴�,!�h�lh�ɯ��h�m3d�2��>��X[ fH�X���wtD�T�w�+�A}�T)՝k*z̐	�:������
�����J/���@>�e�V;���� �矂S�l"|�b�!u�^a-�$���,�y�3'rQ�շ��lY��c�=�q�d, D�|ӆ��s<��B�
_���ڈ�����7�&�֝j뢮6�3�i���*�~Iz���Kb�s��R��xN���՟������>5�'�w#�vQ�J��Q�+)0�P���ܧ��9��z�vW���[��9��q�����@����C4I'U!��)�k�*�@�\�5@{ݤq.\\&�1��&	U>�p��*��Ȑ�y!��'��7�7����z���`���˃8��쉝�e���̵��_ǧP*]YD����@���#��}�p���sE*�&��8@����`Z�v�Y���$ftCp���2�tޠ+�܎Ñz`2Ę�]ڄI�[̙VD��Z��Uo�Hzph�)1�x��?y��� ��v�G;*xq�"Wc[@WI��O���y#Ӡ5���O����U���XK�*Cs���Ʀ�%h���VӍ�ß!b�[�G!%ͭ��0�ATF"�		U+ւ3VN�I�k�_���嘗��s�ls$F���z4���խ�R�ű(dk�h�b��O-�{tv�!��Ү�s~�l��u�� AJWf��Q�Ė=����{�1��<�s�3�oWlA��kAJ�޵㠶Qq�U� �Z��Mx����=W>�߿޽C�g�`���7�{���h9"����i��Х��/?��t%�\F�[�NH���d�7Pwz�������^;�P� �g�c-O1�1�q[Ѽ@7�LX=2���;�- ��4j<�+�ЊK�wdo`5n��1���0�^�5!�D:���uC��������YOe�!�'i*�1�w*��܊A���tI)o�q��z�?��/�D�O-4��nX�X�E(�*�x���'!x��S*��P��wݜ���q�}��粳���+����5��Q�־V��f7�P�2�U���ɒR�3o��ֽ�14�x�o�ɀ��#��	�'��Ǣ����Av7�\,���x�أ�.�y�D=I9˂3�!�i��6Ԣ9��W��B��~ �Q���^�e�ubp�^b?��v���0͖�xI��y�3����Ls�_�ԫ0�煌p��
�~�n�u��d����!�K&,">e�5N���9͈��1����.0 ʝp_cb��P �lB��e��.sj.�ma |#R�<��(���+�:ݍX<�|ӯ��Չ���k��%"����Gn!Y�mvA@B�Ls���!�[�ǰC�onRc6�t��"��[��p� . �:r`�8�P�N�������e�A�[^��/�%�_[t8Z$e#���3�/��9Lf��]ͺ���gN�̲�#<�%B�Һ��k_��"������¡<�w\�M�4���j�<.�
��:α��$0�e��m�<�j�	@*x�������fb9����d��Zߝ�H���a�yFhX�x�@���S�]�J`�Տ���>�pi��Z��w��6�e���������r�|�/ڄ<�prH�菣Ѝ��)��F�<�{�Xle�y�E�u�mKe'�nU�6��*�|6L l��90������y����D���>}��8an�<�B�	,�-�-�I������}��G�a�+��&����yڳM�/Ha}�˟������T��B���P> �J�6s�v7C`J^�I~���fe���ss�_�����Aj��?�[�rX��Gzi9�	#�'����6CF��Қ:{��oc3�Ĺ��ڣ�l~عt�F�����ِ�q"��9΄�{RD.�<<-w��R�w�s����9����b��Ӳ�N��W�!ظ��A01$,]��Ď�d��V\�'k�����ll|��;��.kxR�<
[*$�3�=ܻ�HZ�.�:��o|`��Ex����!�Ã%�&����O~<}*N�
wz�
�n���D�P8ѿ�C_���a��[�R����g��'����&�{!�
����DԵQ8�ejVq�d��vg�-V�@a�)��sP�����k�~W�i��h��'	� �R�G��ۇ�Ik�:r�]�� ���颞��>5�ԇ�?�+9)��3F����bY� �	N.u�R���B�����c�J�b�A��]-�8�MH���
'AZ�?�[^UAC���$*c�҇��+��5J�u3 ���P�F�2�MF#R�M����ZS�q��j3�v��vV���!����/�gx� �?�v���ylf����j�Fa/����%�X�=�g�`�W^����O|ܕ�V	VN�%>ՒC�5U�i|
�����J���.<�Lm.����dRd��؏��5�q��ݕE����Y`�=��4%~y	;��s�Y�A��O�t	��-4��8Nr��0�+F�*�T�����u���]�2{� �V��G^*�a��T�J�sv�������^0�.	¿(��Ǽ�b��L\�AcqݥU�</60o �5���:��*O�n I���ǛQ7�c�����4�]t�y����Yjl��a|�����{<�I���%��΍@sY䛗Aon	
[}�}����o��� �����<�����b�;H=[�D(o��1 z��iE�r�z|�U��
\5��̣�Y��s�	���A�P���p��"����s�z\�%��ȶK�Y[��Ň)z�D!�\�2�~�iM_���v���q��*�vJ>Q���h��dO�R� #F.f2S[%%Ȗi������0#��E��7=YyIv6�J#���/^ω�y��Y8����v�Ǐ]����i8���~����\�#:����D. ����L�nJ �� `����(��;6�kQ�����+�P����9=t�DOw�_���jy79��j�̃���(�~ba��620��?�D�^��b@}��ȸq��d��Cw�	{hs���&�W���];H-���w���3��l8�&��b 9~��"�h���g�[r���� �xk��Ɣ,{*�|ȴ1�����qAH�]-�H?���	��zH�F+5R)����Cx�۩�K���1�ɾ�:8M��_��[B��W�S�t%W�N������g���H�I����+�:�᪦mQ
�� �����pK}Go�Ԉs���ϫ���1��M�����ݩL��_B�z�����dJ�7�	�`k��r>E���;���UГv�/�K�9��!�em�iI�0Y�^W��i!��Ka�R�����	.��6�/�òk]K/W"����;���{�0��7-���.�K�<�N,���V�d�3Z�[�:\h(,��lS�ZG�3�+-5֔J���źԂp�,�g�ؠ�?>)74�P��4%������ה`)͛pb�W�ɞ�Ål%��(v���DO�����2Sjp�Ig_���Mpg� #���O5��m��>�%�v�Cū\'ɭ�5��@lW�@��#���rrk �Z.#�0`菸�}���zם��I�]�N�/7~aఄ#0J�񾁩[z>������Qӯ`e�=ŀ�Gb#컸��6�N�{�]��_3+�g���
˾''� A$���ɻ��l�>.j�9g 
J�k����Z�9�Ɔ���՝l�H�x��+��f�g�?��x����{d�F�
�DߴU��W$b@x�i��M�e�^ 3���'ኈ��!%�!�'[ܸ�t.�H�u�gV��Ig��]	� ���� v��%�2n~�-�>�?���h8���{z�X�CZt#�<�A���(S��4�A7#2�V��kx�<�P�a����g�V;�4c�'S͏�I�p��L-��}f[���,&�9i©��F5Y^>��o*���A-�#ˇR�SV�\DX}�&�=��AuƱ?�v(�iGDD���F����CSO��Y�da�r�(C%����t�3>�qI���)b4�.ˢ�e��I�>�d�z�2?�A�d�x����"�is�X��CĚM="�=��
�?�:K�wz���'3��{w��o�8�|�H�yr��܅��^~�=�6V��h��N���۶���t�/~�حMTb룿��
kޙzq�=f�@�Z���+�x��FN�/�s���G��weg�jb��P�bA[p�q`��<E��x���f��ܾ���>42���8w�7�ْ �őz�P�QOe�䮌��e�06��{�^^XڸsO��m�k���(B��xs{�oiTr��pă?;�Xz�MD�~v��[�8m���˚�>(°xo��jy<#H������@���]~��r�p}{���獹���f�9P�9�Gk_������-�sմ?�Yll��Y�X�;~�"�m�k����vxGe���t��A9kb �|��ׇ(X�@h9B{FV�>�$�p�,E��q�M����n ��7�k1[��Y"o�,�7t;H�ĥ����
vn����x$�o;�R�@���7�h�jJ{:j� �E�S���%#����(�eq��C�q-&�i3S��F3�k$����bç��3��Sv�}9~��<~_�(� �G��`D�~ë�U�j�OJ(���>8iҌ�;�[�8GeyhBĬhmM��_ B�*y����;��o�q�9�X	��K�O����X�Le����?���@v���A�D|̜�8��'܀�{Ϛx��D�{$�i�w��R����7����LtLrɯJ������r�v��m�������
�$����h��>l"�Tژ��a0�p���-�|�;�- E6ʻ+�D��^�jt��Ҋ�X�u<�1��e�4y���A��\΍�YM����?�Щko%�Ճ%�W[+B8�Hm��
�Hь��%>_��S�ɰ�"� ���g���>�O9r�Â�5}u�vO1t��uL(��V���[�U9´X�Z?���e��s";�ņ8��h��P`�7<<���#K�?Q'n̕��Xڒ�����(b$	"��U�3+	E��u�EI�Ϡebu����W <���{���3����D�H*-�#1r��U�0 �r�Y�\N��AP<մkV��P��obn%��b���*������E?75&�ydDED]$����ȡ)_���H	���~�b��y&��%}R�*�G6�j�m+h�1r�d�Q.�vj~]pf������?�@��WAY@U����שs� ��x=|���ss2w���N�������-���
��v�qѹ�����)癁�5D��x���n�	��S���h �dIE@�aE�G�߯,RK��n�׹O9<���� �%fV�M�gqsD��s���e�X����]0��+'� K�:BKL�I�3�;���AM��V4�U���m�;�6�&��O�<��ԝc�J㥶n�f�����C_Q���Hl��T7�b�[MFC�Ӻ�+@���I���)�Y�խ�W�(���	�W�/���~���Yf�
��q���a�[ T����o�Ay6�Y�B$�jR>����D��9�#��T�]M���!Û���������:�$�FT~{ǔ��V�E+�y����p��1��I���ӹ�f�%��7�����Y�k,]3���O�T�1\h���\���a��	�����w�
�Q0<�7�����t`��Y0P�$l*76���9i��r�a��u@m���Y�����ei�`$�Dܻ��z������7�����$/�H��-C�����6��Cx��A����t�A��k�^@���Pˈ���~�#A�A~����H	�	^�WM)\�K��b�C-^��#,W,�*R�=���$�)��z�!ҡ'���;�qҋ�z� ����I=}��hb��]���9��h���p	!��iH�J�ɝ]��}���x��4��j�k���
ܡ��Y�mf;�\r�;)���G���LGU���v�u|r�@�j0Au)%^�'0����k"����f���j�$߈c�����J��:?u/ߕ���H�b�<�<��dI1� 
M�mOG�_gy��[F >M�i��Ȳğ���/�ZHB�7���w!_aS� ��Ck��%yB�v�+ܫS�+�N��4yr#@qI�<��<q�w�g�����8Q�t�u�y�8���W��7ٰ1�_��|s|�K+�|�-����@?�T:m��q��SA����X8�(��d\�+�h��%��r2�LSx�\,�۳����D}q�O��5�3��\x�V����T��-r�z��+*3{�^S��Mq�Z/��;�o� 8��mg���P�
<��]��u1�bb�8Q%v�y5��uL���#(����0
��s�^�[��٫#�I�ۙ�;r �X��y��T�L#Q�τ��A��j�(��V�PX�9�Hz��Jw��Ɂ�1��:�.�����|>џ�󪳑�(QI�kP&Z��즰���k2���Sgچs�"�ի�ٖn v"�������̊�T�/��t%sݹsY���v�4�Yg�נ7�<�s��Pq=�:#��fr3Y1j�ʸ���=��aM�_;c�iU))A�G�@u���3:�L�3�K�������T25��͖� �*@���"ƽ�z?l8�g�y�E���xR�1��V�r�Z�K�˝Q�b��<v��q}���z�o����Q�W4ϙvQX
�oh"6�t�����Bզf^�3*��O9�C�])�M��p4c?we�Ş�Pŏ7��I��OY�cj�bUŢ�:^�`Y1� ���3cO��_�O�4�we�������[�SPg����<�Ũ�&�)=��eK@ߋ�Ϟ)��I���S�P�� A�@<���>��q���"Zʝ���`���-��`�JJ���J3u�n�.[��/��={�T#��Y�a7���o6�>q��R�_�˭9yJҮӯ�d%MY��Ϫ����n%Hq��!�C�[�bI�8m#�����R�M�n"�v&z��ef��#Ssl5��o�����=|GT�[w���.u��Y~
֜(Rx7�R���cX�i7x`K��O����V�3=]�s5h��]	L�h(Ƞ#���Rϰ���ٸ���+�|�+�����g،F~���!�NN�\��6yF���*7��9v��<<��%��Qq>�W+-Qn�4���"F��wY�ʲ�i��Q3�zE	+�7٭V81�g�\.�O0?u�qB?v<$���5�J�}?��c��h h8�^~�������TC)�L��3��s��j��|CU��R��@�������!��}<�t������k�-m~�<Wk�о��K�H-�{j6�~��I|��Q=�7U�#�(}6�XJ�p�Mg��i��@j��F�FD2�u���=��/���P�fC��>0���uE�R	��ƏL�R-T���@��K�D
����^^�yj}d�Ѧ`T�t���[��uv�C�W
�q�v�fə{��ѳ0L���+0�}H�������~|Z��=����o��蓘�*(8��~[��nfg�O���gA�|�=։��z���/�"d�?�8�f������wɏ��׍_glh���O��k�);xTʜ!`�0��).Zc�"1�D�J� �n)eկ�]<��W�r��Kf���H�:&�TK������U�4b��|�g���t��>Ga@ ��`�'FFD _⊚�{� `=Z�`�8�Q�?�ίg
)S��UR�6�&��M�u'��K��*�ٕ��,�Ǘer?=�	�/��AU��;�ѯ�@w_�^K\�� Et�^3�Ƅ^($������
U[�dY��䯹ũgI"���1gno�0r�OjFM0���P���6�����f�\8ӜD�b��rV�e� DK<���+�eXBEѷ�>RD'9 !�75��l��m�Ά�`5y�(��;2��~������;��� �NO����_D��aA�R9�e�Y��ӞȞ��c�n�7� VU���w�6�(�Rط��WRr����]8�V�Z����{yC~�~R�MB��k;�M!�F�:��m+ϵ	IL��W�_�5��[��Gz3��H	�4O|"d��F?�8]Mw�r���q�L�����^��wXau�c�w�\Qܝ'��#�u��y;WN�G��X2�}\&�;%��k��?�Q��38ϧ��E�$n1�"��d������c$~g�ڏ��]	�bm���Ln*6QE�m��$8��B�2{ס�1����PҷY]�UXZ���5�#�g��`�|��0�p��*02&�(/��X�5I�eG�	\�9 �f���J&u�\|۩�J�Q�9C�y89�k�#%�LɹnG�w"�1��t�w3��	R����֗*��� -�?]OQ��=�ҏ���g���k�0&�������� �o�_y�D������A܄�[Dߵ�,����aq��+S݁١b��~�k+|2q�+�����<ڃ�j���dt��D�ʣ�DN�<�'P����7��:���s��c�iJS.���&��$��]���HX�&�u:+>O��:���Ke/$M1�,�	�cwa�Eb�DS�<�ɰ����o^H_m���[)�vV�T��II䆨 �K���a�l�#�(�(�͐�`vR�	|��
�$3_��庍c��t�a���H҇�	L��m�������evR1=Mhǯn��*�G�NEK)�i��}BB}{8�� I�Ok+��Mf�\Oq/���SzA�	�ZV���U��|Em*�C|#�����_���'8N��|Z��5n�	�,M/�2j~���V� ��/��OQ!�
��~��Jc��i���YZ�b��)��U����̺��U��:{�[��&���I,�Ե�Hؿ�֋d�������x�6��n��w��k�fM+��r��-N��ՏM,�����\n�N��X���52���E�u��ۺ|����,ɖ~I:U�*�Aա<�ژ�?d�	/�X��n��hL�|Wp�'�o�C����}0��*�o��⪵Ie2��^+:�P�����_��/'["9z�M��Jg\���y��V��+��1ÛC�N����eF��!���9���5�G3T�Df�nܧ�W���Г�4�����*�h�7_��֞h;���x�����jw0Z80����0�J����:�Ծ�tF���H((D�w���+�}-��(x�xOT�r���9�7T�*�p�.ÂLE�$��&2��N�������b���\r!�}�Z����i��������#��x�k)��1C��7���ޔ�<��|P��%W����|@	H���#��՞�F}|x����e�͍	�4ۀH��C&���	ц(� �Ƨ��O"�,�z��KL�2/�H�o���&������)�6�r�s@ϝ�؈�z�d�٪���a�u4mt_;�J��S �q��wa���H9�Ir�VI��^�-"�ڢ7rifM����_QyXA� �R�T4�.0ζ-}�&�.�5��H�o�U8��f���D�A�q������W�HI]w!��E�y�Ҕ�F9����i=��_Q�hw��Z���������f��s��8H�P����sfh����$�W��'��6Z+G=PX�㨇���-��D	2�R����mH0e����ë7>��#]�c!!;2/x߲LWa����{t���B����Ewů��7k-O��+\������T��k5����?��'b�X�ͥ��ᓨ����fr���Y:j�P̄5O
"W+�!��"��03�pZC)�����xV�.�5h�;�LB���wc3x�U�|�E&�2���$5R����� ^g� �'j��r��G���vy�o��NhKH�>ۢ�5��^�
,(�TNO���Ov"E�3_ȱե�.@��H����2�k`k@Җz�$��}���UC�|ps Z���02�얔�)�CJ�������7�8:���GNG�\�
�	dP���1?�꾠�XӖ��	]kψۺ9R�:�����~Ɛ"�Zz�x�>��H���>̞
����a��׳���I�Ӿx[�G7f�&D��d���	#�0BF/�V��*�:i�&�Q��p�(Hf�#�YU엀�����=5�I��
����i��O�[���<�����?P-�р6����'ܝ��,TYs�讷*��F���/f�Bl{�!L�&��]ZA����Y6].I�4-��Zĸ(�:H�@W����* �y��Oܙ�n��?��O"��rD�{���
羻��Ө�PQ�]���w��ja�v���XI�WE����2oi^4'=��u��)n��0�����2Y��Z8#���_zߨ�a�����ѵ*�V�t�q]�U����%zj�����h-@$4-/2ӛ%\фOA"��Lt0p�ɀ0[i4��{#��{'�\��K���)n���)ʋ����٤.�j-��sCİ������H�c=${"GC�m�n��y8{{��-�d�5�Vr���Qw��|�[�.���Us�qN?z�*���0&��U����p����;�u�"���D���k�fp|��U"XȒy��šE�)����|��ܹW&�����U��ע�����q>i/	�����V"�o/������F���vf�NT.y��$�M��T���H&���\9|�|�D9�b�H2-��Po��G�9��N��������]�r�K(� b@
���N~�D��U�����.�ao;~���U\�`f!q �eo�#�����yqʼk�+��=]�p��q��>����7���@(:m�YƔ�q�V�T�5=u���2F�QM�,���O���(O�ڭU�a*r0���<:e�h����}��(��ps`�t��4O��&/1���'t�-l�k�ǩ%�1]�z�t&RQ���=�?A����un��'�<I����U��`��P�h@������Y-�5��DH���U]'���3��G��\���fqEjtgw�OB�6�*:+�6Ζ�F��ޚ�r^Θ���/��;ԙ� �zS[�)s����8?�2����D��l�U4.��ֺ�e��
��qx��"��{%O�j� 	+C��DH?�5�nM[$���>�~�%��q�O3հ"9�}�ɍ��n��!�q ^~(N�}�����mG�=$`�KM3Y��>���M�JU���[�9�B0��#^׺j�W�q��}S���0o�p�|?/D/����E��0T���V�a��{o��lƔ���w$m�
w��]YA&St|���͏n?Q�t�G�c���|V�y�"(,6vNO�����JP�V[`�8���1&4�X�AyiUY�����Ѥ��\���n�D@���V�Y��B]����?�f=�F�׺t	��._fZ�o�P9���$��L�oN$ӟd�9��Nq?�rM��Ŀܵ P��h��^q��w��=����j��~�6��`��m�c�x��
-3xGv�E��![}���7��e��r(m�.~���N���!��|z��ǵ��vCA�vdY'����BUF�6I0�1�ܜ��������2B2'�\)�J��-CH֩���>�'|W}*M�_Dc�u��{�L�(O��w/qP!�� ���A2���R:5�%�F{��2HS�,h�dgg�䫽5 ���ƕ�b`��������a�Tm�	K$��� �p)��]����5ڣ������k($�~�K}&��N�}5S�g�Tz�ǋ������_��C�o���'|5�����1����ѩ8� � @�ͻ޹[&pU-\:��3~�-�U �"~0e��몿8�NW��v$qc�ML���;�K��w)�+�y���.�зC�׷s1����ќ�K�����6kI��1�V����y��hV���jN<��\t�_�����;?a����9�<�~��D�DDGT�:&�(Ι5����N}�~СL�%�9ؔ��)J>@�{�#>��A�os��o��h������Sp�ɜ�<�k��g�����K̐�S�uH<���3� *���.���N��M"��@�;gBy�r���N~�=� �j����q,x�����0�-��Jᖺ�xy�A3��6�z�*#�녱���8�VmA����3#���Կ��*f:}[]��+'�}�9�#FYc�70T������6��B��JM����8��$�3�.`P��4�SL�o���^-���ݏ�$rYJ��M��_�#��L+��u���f@�uAP�c�1�:�l._���5�o⹠x�N.��r0�hJI�B�L������t�n"Q-捴jw3�r;K'�< ���_χ���ʾ1Jt��p��S\!�bro�֪�R�%`μ���k�x��}��	�����W!v��Ƿ��pʅ�mn�Q
�cx��A𣋔'���o�Q�*��T����p�e)�7Iot�ߝv�r�!�2񽐰~]�l��R4�<x����E�4���W�Ii_Ǭq9#I9Qq����wVx���h�O)R�.�g[O�؜��L��&`
_�� ;j:�����M������Z��r�<|�;0ٹ�?�#5���C()���X�3J�	�l1�����X��T���O
#јW�~�W�MT:��	�"��iڙ���M�ҁiz�'4�/�&l�S�-�����i���웱����B��C O�y|����L�/4��u! ��
Z-�^5dN����D�CS���ײ~��U	 �'��������q\7N�fV�W8:��h{��3GY�e�C��M��Ȥ!Q/�i�]�ˠ�]�>�LX��Cب�-��
���nS���H�y�m�ZP%²ƍ�K�o�,$�C�IsTf�ry;c��&8|�TB*�l����\x���u����Ӄug�*�?��^G�+&,=�l���=���R6����6�[�,i�$Kv�@�h��KB�@瘜�2r[$�'l�#&�$o�y������}������>4t��
��g���)
nV�h�Ek�6�ܻ��8�K�"lzV��A�m�]�b�	@`�i>|�-*p��}J�������,�_(X���E�+wɵQ�\ϵ(�&�(&ز��!b���(� ��T�-"Ag�j���S�PI����W}$;P���MVN�g5�t�s�'.2�3��<����4�� ��Rֽܒ�5f98�>Ӎaz��R�D@��W��дC�SmԠwtA�`$��bi%K����6��+�Ɍ[&*g��A^�}���[0�.��y���
<=����IǕ6��B��Jh�Qf5�؀�)���n]M���^5Ս@�8��Y
�)�E�U?n��G�Ua �px�|���$:�To�6��kAȦ}����hPCw[�LͬS�y�����N�Q~�f���O��g�F� �f�J��[ޢ�0�̲�� �r����x�C{"^D� ���²]��wuʦ:O@1�p����@;P�ZU]P��&5=���	$���]lr���x�JH+5-�n�Czi������z|
.7�3e�L(��	;�O_��G&�Vh�du��ë�⌕ )Ã����dƵð��n�$���@�R;���h��<Ù��s9!e��*B�y+��6�f�J�q�P`�+�u��0�I�vL���m�`�%��]�~N�N0^/�D�s�-¹��B,���e�d��_p����~{uK�'�;�~�c��w����q5���zO�E�N]_x��{����.��%{EM�:X��d��y)���Nkj������
]�'�BH�F�L��̉y�$�a���JJv���7�y�{KJ�zi�<��\�}���A\�g�K�cS��쥝0bk����`��e�/A��?�@�3��b�������uf�y���1@H$Oh�L��$٪�q�[EPO��P�$��V�)ffm@{��8q�&�ʻ̫����c���=l��;bJ06*f���@f�<�ۦVF�E��0K��6�w�r�Ε�j%�y]�Zٟi釠V��_;ڼ�L�d�H��r���6��}y�`6"p��lŀQ�Cհ�[�_���k]��&5�9��9�mB=��񵩽�C��P��Z��0��?�U���ƶ��lܔB�a�[�����/?�f�R�"� 8���&&�M�n�����z	����hq��F���w&��ώ�8^��Aw��hs:TU�V�a�ڄ���A��wn���L�O�><K���<��=��?�H�Dx1��;yeӚJT��]�b����#��ɟ�Cߓ�li*��ȲR�����M��!��#!�m2Oة23��[L�B;�ѷ���p�/�5����(PS�Vl��}*�'ik&�~؇w�8�7N��5�2�U"!�º��DH>�$�ES���]t�,�g�2D	�9����/�o�������U�|J?E�������
��i�^�"���|���w�b�b
@J|�B�qY�g����@��N72W�,!a
ȪCC.���ڜ(�����6yR�Q$dڀY�|���P�g�Z8�� ���PK�=S�
��[���Q�G����)��y�7۹����2��Mr����*�4��,�KI}&*؋�F��`E�����͋��/*������5]�75vc���F�,�r�._H�;<���	�8Ǐ��Z�!`���o���~���}�Ծ�^�p�R3^�6���OTB������#hI�����9R�����w���|���[Þ�/}_.ؚL�)_�EM���g+���p��P�l^��C�����A���y��=�{�9/��#v�;�2�l%�Ή�E����:���r��a������vw��ﶩ���9�i��d��9�<+�_Q���8����=�.(3� 6Y�-K;���ߑ�1s�pdL��̖�Rt�WYMļ*��ܥ� Z�q�\>섀&�a>���@���I��"W,wuVk^ߤ�Ş����L,闳�` W�ȰUш[{;�Go�,�-4�f�}�����^�z�5�����g�ut�k���,O�*���%kJƤg+�>w_�i�S.K1G�=�q{?"*J^C`���&ƙ$�䢴��X�Þ+�V3w���͸ě)S%l��&�!b׬�3�a5�V�Ŷ��T�����a��A�:�n�*��=7����W�Ϛ�n���`��������}�X�::����#�|�t%i7�by���1��c�t�P�l�R��?�h�,O��l�H��%#�
�ZQc�4�8>��L���q��Ua��:�l
v_��H�M�K��ΰ�����'���Ű�~��~����m�=��O��G����4�^�i6�@X���L�D�~���*mm,�y�Ļ��(�!�?��	���0	�����i��D�5i�[��:U�z��'���U�����4I��I�9+�&+�[������	!�s���H#�0)��H�����8�(~?�Q<w���?��8�+�&}i>�A��c����'�H��!�q�h�yc�]^rԢ�lC��^7�O�:~և�4�9r����G{(9�H������vqz[o�g{�3�+���ÒK�˿=v�~J�<��1��ctl������Y���G�;�c>݇�B��������;���m�T��N����Ȕ���=�v�vBL�jZ=�B��@��jh���h�7��f8�LC�n�Ј�e3\��H��ҿ�q�~3dJ��mSl�b��lh���5Ļb�$��������{歸<��b�|ـ����l�s���o���xآ���j��1�ȃ ��Q�o�_|yU��^&
��`����@�½��b�[�K�,����ti���:�=Ȭ(��c8�iљ2�'� @�%
�W�g��N&�'μ/Α]��+*��3��<�b��?d�B�q#���.S�æj;�t��0)fBK����5m5����ө���8�(����0�Q���%u�D�BQGפ@�8��W��&�YDe�61��.U���
���v`aIh
��Af�M����$!K�U��p#��/s�p[%eGu�WD}^Ռ$�|�?�E�FcmE�mw@�%D��j�u�`�8w�����'����q�����`��U�K��r�+y���58ӡ���Ddde��)vIf`-b��;�f��[o�X8���&����� �$�/�//��m@����j�ٍ�0�9�(.�w��u��T��׼}:�+��м��!퉥�w� L\��U>�l�t,�Ӧ
��j�Z��/�%��m�q��k�)�p�2\�>{���뎒�k
)�>�!(15
>u�r��X4��d
�X�%R��Ρ�w�;D��jKsk�'��bj�R�m^�+��� �_�U�-a`���0��<���r��׎��0"�ї��)c
��'`�@F3teC��ֶ|��9�%ӳj$Ϟn�Z�k�`�ZނO1}�2ѻE;��2��x*�F��{��$����Y���^��?iQ���T��@��	��YY�#֓�uU�j(iH��#}�����ߠn�+b�;�wsI/�-�`���,��tJ_'�cN���%�j�^hZׇ��!�$�x6b��@G�y_��V�T�f�9H���$�i�z�b��Q6�{(Q�.� �r5���Ѝ��z:�6�L����{��Q�+���Z#�aw��{����Z�W��y��ywɁ�2�`���g��d������Z�w0V�VW�{���KW������×���E��J3O2l*�����4�rc�n��W���������O�� &P���h7�=��(v!��
�m�6�� �6��W	XܥΈ��E�"���_��)�#�fF�B�r+�g���C+�ϳ
=u���a�p�����̒ߜr��My@��+T $l]4#�T�=Uإj�ڳͱ��+K�~�6���[����s�À�-#��j�`�+`����nps�׍f�<҉Cp._6L�)���S���n��e�����9$��܃d��&� �����~+ڳ�@��we�*��N߫������A-qZ�d�eLN+���������I�4������6�m\]���K���%=ӂ֟�ǫ�%#�.rWr>�����z��Ka�N�æ�ء��d�O"̫,ꝒD �u�����>�m�?:�>�鿌���TcI���� !נ"���&�3851�n� ��ݏؙ
�?.���*��q���P�&j�+~{II�d��I���6=��/E�4�3}JF�*������ �K~��cq�������
����
��y���+�=��?� ���³L���] }���!?ˑ��l\P�� �[-�������y��rmqa��	� �;	��Iܛ��ꃵv�����΁�Rs�$��>�p3~G��gղh�qg��"�C#�'9�q[3oX~�:�.�� ��B'��?�gT���Ŭ��7��	ʩ��pq"�H��3i���P�no�L%����,2��'�P���C�����h2����$-?70�_�S����{�|s���ؼ�ro�q�
�G�Bl�*��[�Yѽ�ٞA�dI1*?l�y�؛x�t�=������c��+X[%`��F�zm�v���:Ǘ{o�1���"���]N*`4X�.�o��HX��6�p-���������ʯws�7���N_k���c����y>?j��Vh�y�$*N��M���E-Pa݊�%�-�▷�U�I!�j�ؼ����ZP�ԗ
��=����f8{"��t��Q��)���JyV�6t�y�Q���ߑ�_	3��c����E�B]oүL����蔂D9L���_%��`Xܫ�b3��S���j�N�|�>��<y\Ø!�E��N>50�
H��Ȱ\�DKQἽ�$�^��f��@<�b��7�@#xK����r#�#���J*�?I ���ŹW��{u<����H����h�4� rD���QH�t���7Y h��z�s|�{��ݗKw�P%O��پ�qCA��|��v5��a�*�"g����b�н�a-��6Z/�QK�@'����x�"zMWi:���E\�4�%����zR?Ii����լ�vim<���̘���<|��I�=!6B�����A��rHA����,�$(�4B&���8��g��Hnaly�'|�O�-uD�ѿi�W4�S��Z�Wc�@Kx�8�׾]T���%G�8	�� w�[�@������Nȟ�a���9M"n]�ϋ�gdu:�O�Ȳ�P�U�y�T�o���\�ȍ�c�;?�T���s��� ytܖ�x��W��}��r���E�(��0��%p[\,���6+���2��/.�A���!.
��p�=�!a�q��P�`X�7�:9G�=[�����Y��o텪{ �e�)P�q	��vEh�
c��Jx�����8����&]��yf�5C��+?�S�J��4��i��1�<��e�������e��"P��w�T�׉�!a��'Q �AK@�P�@���)��b�@�K�������n|Ҍdu�Y����=́�����K�|���C�c�$3>l7�ͦEK�*9�ؗ�����޹����)��Ge��@n�E������ C	�M��ѧ0D7f�o+��SZo.�<��+3
H�,�D3��*��^�(b����-;���2�ݲ��������O;]+;Mj�dzo���?=]����)�t�;Fש��G(�sK_ �)v\&Q�\�H;������u縔i4 T�U$ɸ�:1�3�R��g�U����8�B%��$��&��[�&�K���N `m�Ǚ_��H"6��[G�/�kr7�d~e�ˑ=�x����U���7�p]<z�Jl1ĕ�8kwd���W�OFP�ܓ���B���,P�z|q%�9�G�X��r��1��XAh�ݸ�տ��H��l�f̾6���[P�^Q�����t��$Gz�Ka_W��.������	&aX���X7s�h�jțnT��1loOl	�z`Q|6���#�jhk@2���DY��%n���-���%}��sk҅�X�?��U�r�ᐽ��ߡ+P��̉�|Q��&&b�*{��d"~��9�O{���d��5&�Z�x+nȂ��ĭ1��T=y4��{��a�!��>�ގ��6{�M�Y!��c�����O�x��@:K1G�i��
}��Z)z�:��7��Kbnm� h�aW���9��U��-:��}hs|�|F͙���h��Sv�u3Llu�6-���r����Q�3=��9\ v�i�&��Q^L��2U� ��0�k_�#��	Â��������	e3+*eO�S���k�h��UV�$%\��-Y��`)��+���	*������;I�h���d:�>�?��	^�3-Wq8�Og��˃雨/�i�Ԥ
gAxj��;fD�Yui����6���JD��;��C~z�G��۫��g�ʠG�?g��c���!����Z~���!=�y�n�C
���^a���ÆM.C���Uf�w�����=IG>�D�����;C
'��{j�!�S���3����ެ�- C�݋��Yٹe���ߏ�g����H�|i�����(� ���I�d	b�g�ۛ-q�FV{��|N�]�#$�`׶E2D��4?kFsZ �Wǅ�����'sc�-1Ց��2�c�V�����9�4�#�l�G�ߴ��	�cF^� �,/�jZ7iȀ'�55��\^3�.5���@��	ި I�r@'��JhY@�w�3������[��bi��i�6+HM�U��=���e�C=����� ��W���W�oefL-�⅊B�&��?R�k"��[�o}�('�(b�s��.�"�L���~��-Y0+���	A	@�[KAy4i^S���¦a��x��*v��L�eV+���P��%n��-);�<l!mh���\��S�����^�\�[8�׃|	�GOݝ��>�gN�%��y|9)L���Im����J˱�'����%ZE�싆fa��s�����.�tD��r�+��6��]�8��]��J�
�m�Ɂ�a��s��i/���å V$����!A|�?�h�n����E�QfW���{��k~�0a�p����=EJ*Ձ��ɵp�9�˾!(�
�.�>|r'"����a*���f=����.��2^U�K���A��;�|q�s�W��-ݳ�#U��*S\PnGR�X֟��W�5�ي�+�,��*1����
�2'c��ۈ�G�21pg�1|�M��:O��cY��H�i�����ƥ^^nT�s;A�b�{O]�S��1p��?.�s�C��:f�>3��2��ʀ�C+�4=C�f4��=3�1��TYWsx����)l�g�7쎥�tIy}v�P�/�<���N���m�ޢ��2IJ笞�rq���N� �V�+����N\��#�Z�Hp����TZs�$0'��>��+��,:�[!�ÉA�-�U��Wz�*X��p�!b�z�A����;C('�����my�e�!j@��I�$��#��HK	��?� ��Z~�K��}D���$�QTP�� Ŗ5i Sb΋z �K}���-�j��G�Xp�Y'4�ҍ��ބ�${�P2�P>Wb��_�4�OC5����7�|aWR"摨�CL]KZ�ͨcdD��U9�Z�D �� ���yYx�t�EC���b[�?9��_�ask�����^��S
��|)b8�M���v3k��A��k��![���0� <��o���A�5��.o���c��,���5��aOs�ibO�-��Ї���Hq��9Cb/]��*~ێ{��qz�tI�� ��f��"ں���W�5�z�,xF�b)��z>��s��Xk`5�^A��i+:lU�y�Q,��t�����\���B#vv�*������6��G�b��z1���bť�E]=`�Ң��YE�#�T�qy��� ��gj����|E����u!��c$o��@I]�z��}+D�l���6�s���FG��y5�k�W�Cb�b�w��Xx�a6\+��gMߒ�xkw��,^}���T�,��8�������+����3&�0t�����?����5z������!"��(��^�]���F��H�Q��lҮ��R�<M�/��[��D���Q[oܯ"��X��!\^̥{��`|�!Rf��U�/�Â1�� �g@��0]��
�$|�fm:.e�fG��IA+-&�3y阑��V2h�4�`2/F��ׇ� .q�Dh��193))=6�g�벴�qRQ��pQ]@�]-���̟��С���ml-�&�6C��Xt��@��O�N�m��u ��I���8k&������\�����@��� �
|�͉�$�}>D�V|L?l����fX��+ȌB�tz�#�����	q�Р(���H��"�˴SRdQ707�4|{NOk_k��s|oՀ��OWFΤ_�}]+$;�-8\����r�N��2�%1c�������uK̃M�f�E� 
�v����e�W�/4�+���0@S�G���t��ԫ�(��p�z���Mѝ"7_T>]�_��-��j��ԍ�A���er�뜖��7���Q�/v�[�QiaY���q��.8�������v�(�T\��Z%�9��jh�W1A' �>#>�|��� ���\�ʎ�	i��oe2�G���I�2d"�̷Wn����ziA�����9Ce�8;�-�� ����V���,���^k���gaB�A���l�y�y=p�W ����$\��+�O!�+d�@V]�G���0W�~^.Q�䣣����0��r&vzD�2;:��@�c��[&�9��q����\w�
���n�T�fU�S��S���(uv���X����Ɲ,j
�/���-�M4�	��=�ٔ( :FNx�f@�SCېQ�Kោ�����4��m�X�o�4����D�����,t��M-=�#��X��#����I��7��e��u(��&��p]޾b�	g/�5n�����¼�
55�Jc�D�R�+}�G��s��ۻrm�B�;����tI�I��rk�_U�T��T��MT5�8D���HY�+"Ǳ����
���
x�@���)��_�Y����Z��@����1��f�|���B�w�!goout 5zzL8�
��yt�?��waEn�О���j��7�ZN���2VS 0����%�QaD�# oh'g�~,����k�%Զ=XG�/6�<�\� ���h	�Ǡ�K�3���}T,Zx����'O�t��n���-�h�_����oz����iD���Ծ|�<�g��o/���q�h�wܛY��Țd|�T��t7-s���������ǩv���XelUZQ��>�{��
H�2]J`���+5����A��3V���ke���D�q���;�y;�=^w��ް(Eg��F{4��]0�x	$7]�м0'��V��5x�����HOC������/&�\3bE�����R���͂��~�).+dy�|��Q�S1�L���!�w"!f��\$��)]z�ĕ����xzJ��fu�X��h���\�E��Iw2{�I�-����� �t�Te�I(�_��I�:��2�(Rjʂ��@,3����>�1�@��!>��:֫F6`�I�V+��4<<�
�@�I�op�ܭ�À�侞���y�@�0��I�:�X���ð���?'F��r������Yg�9j��k���3�>M4�	��6�;�$5m��O$�	��H�Ʌ�<�Q!isq�ޟ�C�؀��TQ+�ˁ-'�*0E��墋 ��0;��$�k�ǆsi;J�V���D̴d��� e���T�2x�V�>��6�8%�e�=~!�)�٠���φ\ce)Z_U��p��v4��,9L����J�qi���9��Ա"	�Z�@-,\3b�f��)����e|����'ۡT0�_a�Y5x�Y���w`�8�t� )3�t��]sd���8̍�.��F���)�ڢw4=��Ə$32pa ?�!�B!�c)7}i��H�ZT���/�G)8���3�bى9M/��^iB������ġx�I�ׂN�.����{��S5��5Aw�1z��cA�)
	�k0?w���Io}�����'%,��b0P,aԂ�.�A�d2�Me)�z����E�G���ꚃ�ӧ�)*�n?�Y)]�åR���	��q��u1��(r.(`��<��\G1˔"�E��,|XZ��;�� ����{XP��{�- �w�g�QTtj�'п#�c7�J����K�?�\��z�����!t7v�.Q��e��Z t��XR��@]`��x�Y����萼��PƮUx�N�~���<����]�h&'G��I���Н�N��5
{9�����Op��i6@-c�3�ŧ\[n�����r�3�����Ł�͑��`�BX�cQ���Ci��������\���/f�ρ���2J�|Iq�?��t���}dO���(?���X����s�frNo(���	��}#�8$�����{x��l�)�\~���*��"~gj�	DIq4<�{Ă1�����Y,�T7�
�+y:�B呩�OB��wC�)�p�>�	�i9{��x��L*9� ��p7_Վ{*<��${�kn�e9ួ�}�:�j�Zg$�c��	ǡ-�ox�)ӄ"h�J�Kq�$�9�؈`C�6�R�1��Byf&<C�b4^� �9�T���=^,�В?�~���cA���)d*d�|0E��<@E�C�6�K��ѩ�R'�){�ʼ�6�,��ch����s!����
��kT�Z�⢳��%�Ux�Z���h�s`�,&˴'@ɡ���@���ǹ��g�����L�)�C����e��q-���z'�#�B	��8���F6�b������W�0��=���L�Y�R��(�j2����U;D����ae"�x��R�[2����~p�D�]�%2���]j��_����o7���cip`s���r�i3H�xC�����������@
����z�����'�#���h	�C��@f8�	;�5X��>0A�r�,����(�֨�Z��^�aap�%˂�������,핊�I�ER�;�	���O#-��}?��������f^��j�<��/��2cIa�F�'��-�>ӹV��D��`�~�JtE`u
�%�NRJly��+�P5��7��:����f����d��cN7Μ�S�|l����#o�\eeef���n����U�i�����eu��/_K��E�����i-˜ͽ��J�C��P��b��T��gH�E�Cg*^c�8ާ���B)u���ˌ����MT������W��2GW[%�+I�~����2��I���-TZ}�΢�/cf�v	�Dx�C����J�ql8DC?��=�A^����1|̬�u�ȵ���?��]��u+�G�X[7ömƆ�X�����y:�s�ؕ�Ë�Y����l��ue��XT�P.�P�@
���5/p_���,|� (��*��~>k\��}?�ݰT�T����R F
��=}�׾h��O�\�gk�Fm��˩���ad�؂�z�� ]%U9���#ޱ���#���z.��!R��*�A<�fo�6�*�S�g��1 wD��x��0X�j�W�E�H\��6GX�p�W��޷J�\�ݻ�����T�"��ak-8*7�|����X_�̧㆜����H��?�
�h�q��kf�K_R|-�q�vs ��!���"B}��R�p��[ڞ�Z}��X�s$ HN�B"-���4�˃�R���������ꈰ��p	s��zf����} ����� Tf�l7ot��"����(:�6o�[�0\����#�s��l�sb��%�/o��Z�'��*�g��{��Ɠt"8k����S2P7Iv��hpe����(�7����*���i?X�.��	��\�.?��TW�����f��[�w�lSwS��'���M�y�,rN����1��|k�U�����Z'�h̼�m#�J䷿�����M�R���D7���S �4�(m��i� ��#O�sbCU#Y��8 FmشTy�h���k�*��3�~3o�`��q5���	��n�3G��x��r����uw��xӉ�$�c�%A~9޲���J��A 3�a!���&^r�������%�L*�iy����v�wփ�XG1o17��	��Zf;Z��ָ��(��&�F����v�{,��l%ssi��a�a9�XiD��i[D�t���ȁf[?6�S ��\9�ĉ%���yF��a&]�IZF���@�������kS�T�#�q����*�D��	s��*�{�A_�3��|� uP�`��>�1���0���AOKsp��u($���Nd�!�����cE��"^h�xs�z+F��Fs���t�������{)B!��R5�U`1Pu�w�����
�asRK[EZ
�?��
�X�+���n�كy�S(E��>+��!rMJaE�$FƐ(�)�\]�U�j�g�Hs9 ��jKWt�a�qy+��
���Rp�iO�ى�YOH��� 
ۇE�y',���3솠*'/L{f�9�0�	zT�3J��2�?�i�4�J��Q��*~�X�����TR���I��H���B:D����uo��$м��/���n!s����b�C����w~���넉��v%&(���n��s� ����`��Pe�6���Μ���y�]�� �>�T�c�Bbx*��DԵ}t�&���$���Rb8�/�9�l����	��ގE��{~�g������V���T�������<����w1����9��5��в����r]R�t�c������:�_��q|��3l��	S�#Z���]z]6d�t���`	HǫY�ؘ��ҍLX4��+�Q�	�Ey�Eю�n���w����	�([D��]�n�E��Z��7��Z5�ԅ~�,�-��q�4�� ) [a9��f�b��N��'���%�3Q�:U�R����|)?5!όY��)1h���7�\�+�ڄ���-�?���2R��onn/>���K��:X�+g<Α�Yao�2R
\H�@D�����U�<�
Z���L����I�h��(;+<B�eh"�3��Y;;�y�j%���Ih�Ք�4�>�Wd��7uV���o��0���5�P��u���Xt��hԫOُ6�^�6���l��Ylܥ5�����MU�.�/t����Ŏp�fp3���)Z)���d��@
��y�����Bar�C	F��.��	h�&6F*D��s� '�à����Iߘ��$��!�����M�@�k�iR��!>"���@$�q�����﹪�Y��#|W�4�ci1f�����)gָAѿJ=�x���U\IC��{4�}
��h��h������3, ��OA�NGŽBX]?�G�Z�{O�QT3M�c9��^'O�j�`Wy��+VR�B�q��.��"�&S��c����!��6��6B'�-:d��J���~�z���5\���NYQQ]o�$�U#��O�pJSeI����-*��F{"��>+pRݎ�����n���Ϝ�衧oA�<ݽ�㵚@D�i���?7�f@^�U���aҧׁ��{٭%�5�P���<��.��T�R� ����p�޲���Q�9�K	o<�3��Xp!^i����ݘ��zސ�K`��K���LS"E�`��5�ąL���2��0*�5t�,����F&���r!��/a�_E��Չ����fJ=������ġh+�G�w�J?�N����xQT{W,�fv:P�	|\(x�%�i)�(��T�<&�ٯ�2X��"L��H�Y�S��X���*ɥ���@3�&�@�͓E�T�A�7DuA�>���j�b�a �F7��W%S����:��Q+���m��6�*��i�SY��22ĩ8���C���lT�����	g$���nm��1ԇ�4u�.'��)������MK 1xx
��7 ���	�ͽ�}sO��'��@�:��i��(��1a�D���l���8���`�쟄����t���,��]g�}Oc_R<t��7�[!�8�i�*�~p=V���>��)�G�ժtw��c��@��J��D+{��:ðN�T8(�xFc������ϿW�S�W��8w�馢�n����aײ4��u��B	����-y󺩄u�6V^���V^%d�p�9<����2��)�${��Ek��q�����L��[?�&�M
���צ��f��7�@x3���:�س�c� DFr}ͼ[!�"�sP�]O+=�ߩ��v݅�k߶�?VTc F�����'���t����tU�������(+�s5���>E���[����-�������5�CC��i��䠼i����'p�>Ǜ��u)��b0�"����j��@��j�)Z���.[��S�PHژ)���~�ľP�
�ͅT�FB�C��D��.�=�.��V���AO{^��ԉ!d�o�k/(�]��z,��VH���aT��7	�znl��Tƕ<bE�A֢!߀�)��@��0��w����q$~4ֆ�Vh�L��[dj���$����89����fF�Ͷ`�ޘ]�j�l��iVC�tj�0�|l�K�Li��U+kw��}���7��sXS���O����-�(���U.�� A�/��`A��m� 0��t���ٰ��O4�����;]�Y��^�V4�t�%�^D@��'8\�)�zk�J��jP��)Vէv%+������P��#M��������\�8���%��Z��Zo.{ ���[�zR���Մ-�U�&���@���Qg͞�^�ɳ���B�V�|��S������	�As7�|��ek8�f����(D����w�K�5nt�;1�;�S}_C$3ǳ���c�\F����]8_��vd�>�KqkY�_'.c�d�u�̐�cţ�A�6N��?� ާI Q�GR�qȟlO�3Z���?��I��d �6oR���u(��<b��u���G�a���Y~K��D�2gu����i$�b��j�v7ߜ���gCSo�ؗ@G3`���_�P�K��Z�Es7PD��6�Fa*B�3��������ME���y��I�'c<�0Ĺ��r�la�$��{��xo��Ep�t\u�����&9
W��_�^4h�Z�\���M��8�`�5;[/J��ɡ��R��JJ�U&v����!pēӇ;����7�:ry�l��k&�a��O��{� ��td_r�ՠ�<Y����C.C��d]�ݑ|�<��ÿ#����tnu�^4��k��:7F��"
�@�L�!����6�k�!�٤��-,��o���L9�e���K����1�"�ށH_c�eC���|r��Ť)�!:9V́�h��;A�}>���b��YO������u�y��WG��KH\�*��4e��b�G��d��c�f�X�?^B���5�ʘ�P��,M�WF9NX�*_�،�?4N[6���3���A���swVq�V�h���cdbRc[�9���M �#Z8˂c>/�)�+�b��5�P=$!��#��"-��;�[q����9�7TJ��K�O�<�'�x��f?F����*�Vy�<�d��kA̘��.�j?� .dw��&����y�	w �gw
�C��{��H-	]|>�ߺ���������������2Υ+:�1̤^78�e��I������D@ve�AC�%�#��������zW�>�ń�7���M2���v��&A����B�p��9��%[/]~�K|n�a�(��Z���r�0p�E�I�6?�7�\�W�&��V�s#n�p�X�9�r����y�*M>Ud�xv��`�i ��4m8d�<��L���{m����L��k���:rHdJ+�i�6��g��
]��<|+��3^PaǺ����K��z~I��x��<����G�֌	�<�i\؜/Pj�9|/�v�U.����GH���JY@pyC��9���e���G��o���@��y��3�萻���j5
��gB�DVZڏ��"r'�Q�BJ�)*�3�@m�O#��bX������<�` �M�YJ�Me�$X��~ ���̝s��r��B�&��u�=а�g�-��GG�6/E����k�`ڐn�?�{T�Z]�|Ň��I%�h:�}s��?�qm\?x�)"�����`�� �/C㯝�{�*�Q"�����ء�ȸ��?
��T"1؛
,&&��f ��#p�^m��A,�m��Rt�F)��+gs���Myn${{��B[х���m�|�X���J����wi��h��e�K�y������&�8���=8k���Oќ��:�{U�p �}�w�aS3<�n�q�e���b��[��"��bh���YfP\�T�?dT|5%[�)��[�������G���\����"����"�s�t��+D���o"U�ZJ�4�K�jwϡ`�ǅ4���/Q�H�<(������Z��_ZkKV�$s������A�P68�!�F����eӴ�J�Y\��H�($��F$����@�E��w���mW�{v�����g�)o��#U��s���4D���2-
�����"`�	#�Q�N���p؛Jߠ��@(��$4�*Xda�ج�F��k(��ޢ�6���O�,y�S��#��yd��ĵ���IS���MX������	t��R��\�}d���x���U)jX�#?o�L�e���XRX�qa]���4o�	���;1���@B�_h�#2o����y`�9)#o�Rt�W��]�	�q�}�B��������	k�Է���2[`@knU���.�yA#𸙹�LB鯤�mvC��6�\�-q�x?7�!���F�9\���`f��܌-�fU�atˈFQ�������6�a���>��qP���������EDR?������$� \�%}M���i!S�А��a�+*����$ٳ��ǓE���8W��ǣX�=�:���V���:��J��zsykf���5J�M����-W_eLL܇n���L�S	e.~ղ*��%D�Yم>l{���_i�� �؍7��>�Op��!�À�.Ŗ�05���C�W�H�����Pz�9Ά Y��}�-�'�0��@o;�����C�pa2��^x��#�7���v���!E��0M�z6�"�g<��l�_�����W�שHt�/)
nr�v/����$Ga�uf]��,�:əme���P�1���p"̢wU�3P�<�#9�?��m������._�5,�E�p�
ւ�G� �Ī�A��+e�z1��E�Q�]A�9e�w�������;Ÿ��4�����MD�|24]ߔ� �ʵ�kfe�s4��Ќ�rWoZ��%��hTJ0����H�"|+0��uq���{�1�f���PCة���p����@�k/'5G���	�2��Tm	�O�z���ʑă����ٴ��y��}�4��BZ�^V��m2w��,w�QY����=9Y� ��j�J6�y�4���y��zGx��$b`�(g~�R�S���|I����O��#�G�:9�������?��8�r&�k�?��[�4���3��֪�ȥ�	G8���B���9�:�<+�
'$`x~�-ҏ (m��CX����b�H(=:7�<UA{S �]n}�)<�]H�C���yA�����r�=ip2�|��dKߢL�s_n�����g���CO�R4UCD*�sF��ƒ@8EL�^��Qy��3�a�tCQe�~�>Y�9p���x!ɛFAeإ�z��ڔ1�s!߾N_qFܑ[��p�0�,��t�31M�%�]��Ł������.�Du��.��&�%[����R�7Y�<.XԘS��.3�t��ʗ0V"}c(B���ZX-���B&�6g��AX�Pj.f���7|~1��ћB�ʗ��i�κ�;��=�v�n��z�*��Y�����;<�AmֹӐ�F�\�=����a�/�"�B��mE�� k��v��!���ty��u�c�K��Ƥ�\��~�V	{�`��P�RL��ZbFӗRN�����q)@��*�.���  [��r�^l�×>@��Y(�d�{����w�)�B4z�c�gu�7��v�s�{��?�ˑ+6��-�#Lb�oP/���Ɛ;�������0�eP|9-����6I��3�-o�[�+׋7(vV#ݤ�i9]���v+ۗ�=���`�y1c��y����[#<��p��cKE96i��(>����he�\ӝ+�uG�OqS&�q�����Y(��G98)X�8�F��\fl��ð ;����d�'ڝ%!���Yq�9T�v�ItK|�� /�ևT˸jE5�ڝ�uS[t�"���,,�9��9
��f�C��(��9�f���Wr�Z���sG�_�+f�>�	 DF������7k�|����6(����6�~ۙ��g?��sg�v�6]8@Xs���.����9�g��pj�q��>m��T�Q�~�D=àrPO9N���[����9tFT-�ģF6%�[�f2���VxzJҊ���6/��#:��h�ǉ�-+�����{i#)||���m�����Č��0�u���[8��̑ɟ�-8���nnC��֘��b�������D�J�(%'s��z�������L��o�5�Y>NF�	��5L=���4�8k�8�����܅v�+ٕ�-�j��mˡ	x��B�HS�i�5>Ȫ�r�O�8gۼܲ&QS-<+�/qzJ��.EЂ~��(B���|PN�����֊Kg����R�8} ū�+��~�e�`v�DWt�͜����~�㴒
CJ�ʇ�ۦ��I��!_Z���h,�|i��'?GĂ&����7��^ ��l���Z�M��s���`������ -d�p�(�J)5SS);���Ռ���Z8|�`yV��a�wpZ`;zu�������z����<PclS�|ys�4S��j*A��6�(\�K���o|$�e=v���r���I�����t��=�Q�TA(���הm��ˏ�P#'{XDy1?,:�S�Z{���nY��C��)E|`V�1�3����,���/ԄW�& �*�Bz���IK�+rN�D�5Ge��	���9YFx��I���l�w��ˑe�[b�R.l��+�S��3�>�:��R�W�鑄M�F@�΢I$g������<�r�%����W,,eC?��HQWMݣ:��tl,a� ����ScG��q&�^J�s�u(Ԕ��l#wTKWR2ɴv��i���=��'A���
c�R���.�3"	��ѿd0L��k�N����k&L	��p�޴լ��^Z���j��}U�I����9�@�CX��4xq��������u�����}͇���T��w8������������ʙfټ��ch�G���(�D�Fʛ�h�-�]�%~������ �k��ڐ���F�0���$5{m��5Q[��xY�I, q�LQ�U�C=*3�4P�y3~M\�o����C�Mp�B�:����BM�$�$~���hZ"懮���z��>@u�E��$���;M�b�OQ��cg�Q�d�X�m�X�Y��V=t-���/�$MD�������Q�K���M3E�
��/zP~�z�x^&c讅�'CcYGߥ�X�8���s��/B%dA19Z���dњ[,U�ˠ��ꤜt�KH�Dg�_&�š���*]	i��F�K]��7C1���=��A����ڜ���;��{Z�Y���-u��vj#B�wǮ�������w�n�@��T�"=0d��l���J3���w�qc�0��\���>�s�r&�{�H�7�{"�CFɷҒ�a��t��Z��R���DD]����W�9GW�͔��x�s8\�J1�.�0�Ƃ�HpM��i/�k��fLlTa�2i6Q�f
�k^����؋��	MaԄ=�f��"��-���<->>����(����@K�ĭ�Y�2���Y�p*��+
�8�9TȲ�&� �+یl:��z�T��:�i��a���0��N�(G�:���-2�c�&�ȵu1 ����,5�zB?��nVqYPƏ�����،���`�]zc���fA����x�?�9#(����wκH�?�}G�\L'd��k��\}�r������	�:��Y�&]C:}�\�ע��KS��"�U^N�����˟&cv����r��i����U�N8��UDj�ew��yHg�욱9�x��+mD�q���F^23̗�ߚۅC�A�����DO��oq���E�ĸf�pe������4�᎕�vJ��L�����Dԝ�@�g���ULYe)�,Q�"��2����aٛN�tx��@�C���c��o�9���$�E�����E&�5bj��G��l`����AZ�,����@��:�sJ��W����"A�"�&���!#Q2����������{-%�k���_F�B��{�k�hˣ)��qЎ�>u�]n=���BRʹr����}�a'�����v��0+R��v�p�]�b�i�r�%�f�k�����W��y��ȍ���o�Ď�A��@�� �F"��0��T��I��������q�	<ثH$���N�7�[:����S@+���[X�,��b�ƣ��x�4OĞ�F�.����������ݳ}4{�`��cp`��	�Q��K{K�N$�n;�h�[��ԉk�p}��]4W�d��+��Dl(�Ѱ�"t�\�̒�7��U���*Ǔ��rm����@�q�������B*��L.���[�'5��
c�!}�ݛ����,���؄� �_!��ͧiƶ��y��aq�y�!�kB=t�]+�bn/ۢc�m��5���mӗޡ`&��dAa�F�2���Y��8��袜$yL�{Q9xПN�-Vm��=��*"�4�t�
5��V�]�.4�(A�f:c�?�����'l�%��Z�!N���me��At�R�pOL�0k��p7�v&w�j�|�/P�!����P����ԛ�!�"���C�3�h�e��
��-"|E�Dm6����d�t����T-2��(��!)6���RE�0������xJ��s�rt���U�=Օ�G�!���#���t�d��V�BW�%e2�v�fR<<�%���aj�>n?�i�|�KUн잘���b9~
�oR��>~擡���z�� {�1�Q:�Dh�C�k����U(�bva8���3��y!��־�A��ҍ����e.H�逬0��)<��!N���-��<U_#����oZhנ0��2��ܶ�.��.#)�.M��_�tڹ�pԉoH�U���j+?!X��z��?�W�vǇ��x�&��[�B�IJXձ;/y��u]L��4��_L̆�R��W;�/���Pl4�E�;��+6����eA��KT���lP�b���l5���8�=�n1�Z���6�iS����,�Y�]@�>0xuM�Az;ۺ��7.k�����an�_hɶ��"�@E�!\p��܍���`��d��TE-C�PjֶӦ4�y�?,e�;y��|;2���@{���Or̓��)x1�kĜ �KJ17Nê�^�^�����Y�gGc1,E*�2{.�q�Je3����v��H��շn����G������� I����s
AL{�`����Y2�^u��?y��>�k�[�����蝓����K[��j�����8r�t	��Z�o�e^�L��U��-.L���Z;��H�fϽy9��o!����dPo�h(����a�L$L6������N�:�d�s͈�u!�7���ɝ/�t�N6���7[zO�*�s[����^�'�������w$8A���Γ� �PLQ�cu�a� �65��d��lGt�^�ȭbh�Y��;Ih=�#�b�	������R���X�*�|����%�pLղ��գ.������wX�v�����"��&���[�hpB�?5{;r�1����.��. 3��k�����<�ы�&�ga��@�r�e���]��d \]��)�v[�������	e>iG�?�^o�5]�0>�*��Js*dϤ�2�1%ك��Ǧ��:a���T���p�Ǟb��k�9q\�EwX�\�mG<r��{��}e�O&~iBw�y�Q��#
�m��9�z(zg&2'!y_��h�_A����4�U�T��8@X�(�ם9�7�kv�gs�͢$��e��AJ�� �5/I�Iѷvf6P�Xqi���J��L!�3��K�i�_��͢��Sp�ȍ���v
ߔJ�b#,��"S�8V���fi閱� 5JX4�8�_�z}���ke2įWvTm�o��8ܕ.M�&�幛:R���ldC��5�����k���Ҋ`� ��6�y��� I���M<�r�'��#�A�ؒ�h
 �kqh���6���'��E�����$�E��_$@/Y�6o[��Ԡ�g����`U�͒���e�u�w�ɇ��~�N�M������<	_fZ�U:�vG,�����Ia�Bby|��2R,*��Qy�J�_vxo��E�#�p3w6F|y�yW�nm�f5f9���NA�V�Z;&af�L��/`hUO�*eIO؊��t��͈�w���%�<�����l���4��D����a!������8R�P���N�@��Ɨ[�e�������j��F���&�5��s��8�".�ZNY�X:,�y��#u��E����;&���X_��~��#|zaZ�ˀ.D�q�k��|����rmۡ�Q�Ƃ����wVrk5*��(���y��
��!�jC��#DG��Bī��%%��D�z�Y���6�
2ab��71/�D��{YV�ҍ���v���F�����[����s,T)��-ە~Y<�d�_!�R9���L,�����2_l�4b~z��v����8����P�>|j�+����Z�dE�^��]���2$q����`�}~�R����!��v��&)^��Y�zM�.5蚞���]%�X�4���+b/bP�)�S���M=��n'M��MC��J��K���u5�^�f`���[�.�=bƔI^���v�oR�^ܽX��IbO�i��9S;�iP��<._����.1���s��'u�Sw `�Mtҙ���lu�F��%TH��0�D��q�@�h�>|�W�[�~dwJ�)߃9:�ʩ�#c����/ЪMG��Z�г�|*�_�>���ӌ{�7-\�y���N ��6u�$��q_��ʿ�^��2ں
}Ћ���E����t�P��V�TO (4q��C��금�~*���PIA�M��DWKD#n�`�)������
�Q����T%%ވ_~�z^~��F
-���cknǰ��d���0�e�?�޴���b�����|-�'%�����C�Р�S�rQ�L���ޙچ%k��#�G��n��~��.�ɨV�貉�Z��/��s�MȚO`ftqh��3�-�Mx�܇	$>N5�Z�瓙�E�)pP�׊�f��χ욯h��JM��=V{���[F�u����҄+�4�V-�f�=ۡq�G���r
� �He�'�BΎ���ާKO�~��O�
)L���Z���ͥ�X0�y�ٲ��5T�����:���5�֓ɦvښ���bb�^֭��^�������׮@M]rѭ��+g3�Z��?`_P�,'�0�8|'b{w�Zq��[�/*ǚ����G���)t�z͝��,�����O>�N��ҺT�� �N�?��'R����_�׏�񈐅;�� dm>n�n�.��B�ZuТy?�h��0�:��0�����[�}0W�[�R�Iy®K�����F܌�Iй��9?'�pH��B�]!�>�3���U�u]슥�H�Ɗ0�9`�X vV��Q�@�<!z�S:t[�謷D/bzW�D��"/�?��	y���H\݈m�x���|j�>ș�b���1v���0�*W���Y���̂t����v"%��y��e(?�f��M��S��3V�6�N�R ̓�k������D\�l����k��-ϡr��q?��O��?�k�V��W�8�2�
��t;/�chBk�!.�'g��Dw#�t`6�H(CA���t�i�-���{p��C��<)
�BA�ڇ/���]Գ4h�fB�L-p�a�O�W�᯶erԯi����v�P�3PU݌��	bWxs̺�� ЧN�=Uw6�R��ՆQ/WFN�1.���)G�dц@@r(�3�Z F	e�g�$xj���DV�Q���Cij�96'G0�UА(U��gʗ���F��+�-A>΅嬃h1$��/�'�ft��:߳�CV~�n�B�Ǘ���4hݕ"��u,dh.����>�5��E�x��L�	��}p����X60�eZ��4�_��4⥩�aw{�l4������Ĭ;/�`i�x<�˴N/�c���Տ���MD�`0k��&U�sEŔa�C$O�����Rz\�y/-��z��H� ��k���,7k@{�k�K�k��HK
4�]Փ,?�*��m�4�� �S��J���^�V�w�����$�z�	����w11���d��*�����Ҷ���d��氬��4�
Eh��ȟV�6>���{0ȑlW�pIMvB�+1s*��v-1��]�sl�j�k���c@�_���\���Af�Kސ��HNp�\�J,�q��{x|�t!-0��X��-g�iw�Nq4��c(�?*�#6"*HJ �w)�w�U�<�1�-Kwq�� nc��[�E2�LӋ�����Q�nV�e[_dc�v	c�|��VQi�"&}�s������pj�
�6�\�o��z���W��L�pk=��Xh�����`�_����>�@���x�cJF��)1��n>�{��M�5�N��z� �Z�h=�z�f��k��2Ky���z�����3���v�S~B�wo#�
S#�eKC�b�(��=Q�|�̓�i =�x��-f�7|���A�f�����i����1*��?�MN��lEG����#p��̲�g�~�J�@��p� G`y�ϴ��7}!�d}N����Hǯ�¶��i���%�۱G��}R�U�h]T��?ޮ��rBFa�6sb	P}zs�kH���ߚ��&�ٜ`~��#pҷ*l_�?_�����<��}<��繂��*%���	�[�3��N}R=8�x9�_�8!aشx�w'B���S]�!@�K�uq+��<�@��r�ь:`��7�nm�-���ѡإ��<Z���i9*CȤ��X׌1u�Ƌ"�u�#\�f�q��Ƃ�ˆ�J�� �*v1��3��|�H���o��I�����ir@!d��gΜJe���y�LW��QP�/fKS2�ր(�t#���uQ�$���!�����B��R��J2[J}C�_�ٱ�T�6�����=W�H���1{JF�ݮ�}�K��͵�l(���cV/"������l�Ek��)5@���5%q_���q5bb":��
��Q�)��+���h��DGG�+�e������
�@]d÷�i��2�E�'/���X�N"�Ͼj��d� ї-�F�an�"��^��o�Ah1~�Q̆υ&�����8.z�	-�i���Sh
���C*���sW���f��@���z'��i�k5�2�cz�ux��WR))z1��N�s�}9�(cc�6ۉ�+��i��W4gĝ�m�Ә���_@��)���n��»7�?��?����� F\�Ӽ�G�7(ԓ�~�SVN�u�M��a$�Eq� +�v�88�T�]4�ս��K�$�."�U�/}q�����0��������p% ��Yd�j�ښ�X���\����MI��������(�|���'<��P^�
�q�t� %;�m���ή���Gl�'a��P1�V\F��J7}��Ӌ\p<�d�kc	�mk�G꼭m��>����-�U���t����u�f/�>Oc92��m�n��`WΫq�Ռ�&{]�)!��Xt��)���b/ Q�+�����b5��ؐfD��B"�2)}_��e��+�2hcv^U���˿����2�	CX;Ģ|B?��V��_��vVe��n׹���z>YWD��[�j��T�y����⷟��8�O5�yb�ϒ��dn�����R�&+��Wmzf�$�¼É�"[mmllB��s���x��.LL�v�
�-���T7����k�����,�����^����~�Ex*��z���zy\��23��If���Wb��"��Z�z['��ࢾ�O�gB^���� �#��Gҳ[�~ ė� ��c�Sis�H]����M�B��C"�o�R����	��~���|��YC�|�%��D�ki�`c��j�����X8�����ԯ��Bf�U�4�
p����� �|Пjl�rnđ�� ��՘kK-�N�wDCL��tt A��Z�*�Z����,e<Q�)R����O|��dۆ�U�nC�"Td�|��˄޿�`Z�D�A:�W���T�a���H��o6$���tE���.�Nm��~?��H��y� ��� �����e+���8�:.ޑ�rKF(�;x8e�B�9������Y�+��k�vp�|���r�sMhR/�j0:H��}p�ўC>�e�Z1X�S!���4L�V��^斱Z�����#h�!P����0��W�P�:����#-�Կj����+���Ye%�ߕo�H�G�w��/*���̛s���\_aۖ��ּ�ź_}���N��$]�W�oI#̠mA���T��)w�!�e��5Z�]]0���C��y|u1F��Mf����9�)��n���8�v'�C�2����bc('j���OW���0��`�m�g��3�v�6qzKvwW4q����=��H,�}���Q�_00!BD��&�EI�K95@�x#PD�J�;��Wq��Uq�OLJt�ݯ]
�r&���x\E_��z+���q�)��_�F� ��m�����E7�$�l�� �,�t���Su	o�����u3��DH�c��lf��Ԅe�� �e�{n��Rd��
&Ɇ���s��$��RQ�xr��Qm,�7��u�]:"�i2��F;�I���Eor�T��np0�E&%ܟ�~����jl�u����|� �Ւ��z(��O����l}���
R�؄�3P�a9�"i&ד��n�uhڴ�C��u�T!?l�3g��)6�J1���
0���mfq��%K��c8�.�J��Cm��Qd�?�S�EY �_�'�?Z���8TeY A�-^�Ff2T��=Q<_\�����J��O p��w�2�
�(v��4H٣$'Gp�Ժ�fv����	�A��ּ�^�^��}��Ǎ�}�wW�X����Px����}���i�X���2\%>>���2��;�x�ܾ�;RZx�ܻ��V��o��&1�#}�v�g@A��52l6�X��3��|`�, /+�q�^��&[����������Wӛ|�V��~z��D�&=�]��~zT%�hx�&�����%\��EnBnQL�[��DZ�ɑ޷0	�|4�H:�����w5����b���fn.��=��P������g���[����l���;;�6�D`#�U�R���G���٨!Y6<�4��d�f~���߱(?R�jؕɮ����Vu� �D@��b�^Ke
�ޠ�1ė����ډPt�_���z��~�!��_\T�yd9�鬃�v9����_a�908�Dd�%*�>qd�|�x��`��H���Wk1���t*Y���-w6�ͽz�rCI�gnI�G�hJ�?�2�Z�b��ݵ�l�(1G�����֖�nT*����Cp�$��=�����VÍq�Z���مʟ0(xQ��f���1m=z�����;m�AI�?���#�d��h�Ar��և�����e��i���<V<�n���l�W�W���'��X-e�^J��>d���f�T��d!�O8�iZ��o{�y�6��v��3^Dq4ڻ��A�/VB�"�-xl��Ж���2�cӗă@������g�����]-�5�I�G6�)w�;x��fo/K�;��7�=~;U@�@�U�B��_���>]he�Hbe}�m"I;�x�]���~.�/��ȝ�~�������T/�p��8hn'�>
�Թ�����C#��л�ĄQ�b��x!˿5����n�M˳NW�����FY�![T̅FC�F��J9i�.I�O�/��W6��HVE����SN��ਖ਼��d�ؿ��'Y����X2�C_�n&����v�گ�����M�L�)�p=Ay_�{��ŕ$��n����v���!��o���"�"}����*�$y׏HC7�p4Ϯ��������+f�S���K[��Ja��Xq��)�z�\^�M�P:�� 1�j��6/V���Q�8���.:���U���C\�b���6b��V��>�4D~c}���Q�Ǿ�匾�ɞn\}���f�*v��W@�6�>R}(�@X*!_�m��n���)#֤�ѭ��)v4�����c��fd�{�8�gRb! W%��	l��/U_cմ����t�$����c3:�d���r��Ί�,�F�M���QJ~��P*ك?c�<:���[J���}���/�iU���֯�P5��}����31q�Lj��B�4���.5�~+�i��CՂ�j��]�oDQ���娌�VX�DR�,�W��N��:l��Q�������~j��j/;��Fe7�L���/�p�&��<��|)��f����D�cK�&�W��Za�*�fœ��5�e-��Z>L�@�ܔ�f�k
����o!��i'�$�V�]f��+|�_s�WZ��ꊿvQ1�L\S�'G_�df���m