library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE ieee.std_logic_unsigned.all;

ENTITY LAB2PART1 IS 
GENERIC(N:INTEGER:=8;
		  K:INTEGER:=20);
PORT(
RESET:IN STD_LOGIC;
		CLOCK: IN STD_LOGIC;
		TERMINAL_COUNT:OUT STD_LOGIC;
		Q: OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
		);
END ENTITY LAB2PART1;

ARCHITECTURE BEHAVIOURAL OF LAB2PART1 IS

BEGIN

PROCESS(RESET, CLOCK)
VARIABLE COUNT: STD_LOGIC_VECTOR(N-1 DOWNTO 0):=(OTHERS=>'0');
BEGIN

IF(RESET='1') THEN
COUNT:=(OTHERS=>'0');

ELSIF (RISING_EDGE(CLOCK)) THEN
TERMINAL_COUNT<='0';
IF((COUNT) = (K-1)) THEN
COUNT:=(OTHERS=>'0');

ELSE
COUNT:=COUNT+1;
END IF;

IF(COUNT = K-1) THEN
TERMINAL_COUNT<='1';
END IF;

END IF;
Q<=COUNT;
END PROCESS;
END BEHAVIOURAL;

