��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#��m�4���v����\ϺLO�g�"�g%�a�^�S�@(X#�a���T��R�Z��W�$����"�|Ԧq�ݾ(�?S�T֤uy����h��
�Ƅ7 ��+�щֱ��8oq��B9X��ʸ�J��*�ږ1�$���N�E�"�,���xv0v�%�i��&w:O��N���z"��8l�VG	�����_����L�Y_�$�('�X�׹	aH	�X,+����,uԺ���>Q.��
����s��z�)�9,�D=���/���x��ܗ҇Y���n���i���@�N�G�
9i�7"��v-��̩�^y`q���F ({�9C�7�nl===�x��h��Ă����-�D����U�>�i�Di�<�y�M,��c.���{��pLe�E�-d��̙яﰣ���3��\�K_�+1��}��-@�o���c=n@%��İ	u=��F����fZs�@��,�S7Fe�������ku0�|S|W���.{����za����'��Pj������Zl������%Z.�6{��(�s�o��nH�ߨ6E�co+�ܛ�; w=ߘ{�E�1yz��ڥ�GR��۩�-��k��c;�ܱj&k�ˬ+Tft�shMU_ra�e�|��.�eĠ��xs������������o< �6�zvw0ky�tNI��u�.��1��� ~�N���_$�J�˔K��1��Gy��������(`r4�%�|�2w��W e)������4:`���q�T��զ�ޠ�$G�0*W"KG�L�S_P
�&]�������'W�$Cg`=a����A,�l"��}�>���~kzE�[���G^&$�ZbY�Hʑ�������2#Z��bnq�ٴ�4�Dgs���B�UCa˕B?�3��yO����"�Nم�r<@��zǳF�� �rZ�?�y"����w�-�"�4%�r��,��V��^\�0���8@-����aAe�{�K*\j�"�$���+�/����C�s��9"DyI�{;���E0�zE�m'��A��4����O��հ�_�)/�;,<�Hn�p8��yŊ[�����τ鰫x�Ԏ>�:�JM���i�YN x�b{��0�vB�Ʈ4�4&*�(�Gq�M�u����*+����z���&�4<�j��[O|�j�1�<�������R�f��ڂ�xԧ�\\)iPU5��!��v��7��zR��u��E�Z�k�9@�u|��>��_�bs���~�)�'�-�����"��q�\�ݦ������i<�b	^=�A�v�q���x����4<H!xb6(C���lv1�F�ߪkO��W�T�"g�"�y$�U?Y��IΡlT���u��
���8��mGԬ�h�L��M~��9���`���?�	�%�8��9MO���VQ$ :���v�ɯ��yQ�����A�)��9*�cK�E.�f��(0��}qf�6�{�u��`�4_�a2����g��-��]^\3�f����HPxi�YBG+t���u��A��;�QP�4Oo�`�:tF:��^N8$��dU�'
���"�0���e����}x��K)�w�~$��=��c"�Y�� ���E7 ��x���5 ��6�A�c4����F��%�N��̑_h�=�Ѹ?��cg~����]/l">r�t��OӍX.y�s4��5� ���tUJ^-��nX_��&�����Y9��O�Av�g+93�x�y��FMo�Jx�� ��W�e�R�[�՚Ƞ�B�d�ω�2@�]�H/W����S3�JZ)�I�a}�1���J-0���������(�l�.'��u��FR��Tm��ARf,�,\߼Ӆ���(vf�hO����gP!Fg4T�R��M���`����� �������(���p4Z��L���rC������Y�QԐ�z3c��jb��"�G+�j@!����'fl���΃�1�����DtIw��w�ɽ8}�_��mO�K(�!��qT��?�ʄ��	��LY�3��o���,�bH�|�����U��7�(?���z@g�o�1�#M�-Tc��.#9��ؿ�����_k��9m0��e>�
2��7]�l�<|��]�!x�y��^5�4\ø ZIoL2	M s�H���yl�D�P�C7�X"f��GoNd�>�a��E���ƗYf���tc���U�jsl��w2$�6��j�*:|�yMb���.֦H������~��Y����F.�sDg�O�T�^��;!=d:��Q�J��Wџ*X��y�k 	=ș��@�ظ��NN�U����.�TSi��C�����M��-�	ߠ*z�����H/�ߝv�p��c� £�.7�E6�C����,YϺ��|����Z��\w���l��o�I�A��ѹ�z�_��3'l���ݔr�y��N�.NL�D��^UPǮm6iw�A� ��k�aZ����/ϧW/e�uqF��~�#lw�>_�R)}mK����O�� ��]؞�������2�ߘ��M�!��gS�nۈw�Y�*�� %|K��pš�r���E4�fH��E-���:� 宏�SEG��#p"DZu%�#��pvv2&�N0cr�]�~������E�����O�c��:��F�����a�Z�|�5�>�جKb�2��@E6�.N�U�^��q�TMXLho1�[Y~�=�ǲ�j������=�+�� R�b�f�Z�Zxk)����Ce10_Jg������U$��=�I����un�x@��e-h��ut3��L���1����+g�i��#Szx��o/q�P �X�8i4���J ��q�>�[��
N�C%S_���T�W�S�s�O-��[@=�#-�e ϴ�DR���C�w0�����A(�H&�{���|F�@I>&,MD^���DV,���Q�P��\�≷'�!����;�)�eo�_�{��.�b��J{Ԁ�t8H ��,>s2��?�m={��i���s������ A��W�1@���\�u$ˌ �
{(k8���'r������{��ڭ��M�\5/�9�&#��\h�|īR�zc�����ܓ��2�ׄF<��v`�Q���g���=+᫻�Q�M�R����z�,de�J�ۡ��c1#��$_tm��r��O�#�����p9$5�s^�����'�%^!��7f�<��]�;�6d]\��v%o�ۜ�d7���+>D	��eY��u�o�����48Y-էu^Qa$��1v9>Ϸ����摈��ƘO�p�b��xy�E2�#Y2�(���8��O�'�-K��Fp����W7�;hᅎNm��/�P$��H|�?�Ӹ"���ei*���@��B�8�3��ީ�(w��LJN�h�]���k[9��3CA�����>d�S5�H>T�vS�Ñ�M%�jj����G���%�}��ȑ(nőV�e~��|��v���Zn 4��أ�2���I��'�dO�Q��c6��� ��3/�����2��j�A@5�ބ���gVX�L崐���;�3��)Ϩ��p��[8�7�Fo��:cC�2M�����B8��Be@.����形�art�Z���"�Tђe��+��).k/K�ϛ$Q�a���S�biFɌϏ���q��[p�Ɵi\��3�ӛg���� �+ãP_N�5�9��f�:U~1���+����,��H�vO��ӱ�?9�����%
�x��� K���F��������Js�mQ�S�����\���oR�<�(x^��OQ�G�����m��F.{�&0:6>��[���Tۏ��6~E�L�CYbH�B=kI�4��umnǘ^��Ʌ��b��H�l=�����`H��'O; �u�-5��l�1f��r�̱gR�/!X�I���r�<��ʓd�_��<��mU"�t#�4ޥ�W�5�e��T��cåG�MA�������I'��#�w	����x�
����C��\$�x/A�}�m2�Xך$nX�bpVŧ,op}�{k�ŮSũ�D�7�蚁�h�u�9��������@Sv�d�I���t�gN�k�����A%N���hb����$�0�>4��#����UfTzsi%չdr�cg��"@l4@�����ŵj�<5�r�h~�Y:�r~��qpN����X���J�h�Ќ��)+{�s��_����X���uY�S#I��U�ӡ�7Bi��`|��k*���L�n�W�u�&��:cc1~0=�Ӥ�-c|�3��6�~�B7;�VM�������M�A�ك
ډ���}�]�Cѹ�[�|��U7샵_�o`dN`��׬S��F͐2���k���}au�vdo�N*+U��r�X��Z�2�_a���Y5�-�a��/�mO�݋����6��g0�0͡��1�Qp��	;B9�e��4H�!�yGN�[�٭o4�t�Z�" c��
�4����#�e�{NN�x�t�J@��Mʮ�@�.��r$���#>?�	s(���[��㏾�J����?�I��6|�����}�KLt��`��+����i�p��Ac_~��Qβ�~�{:�i�dP}�0��j�F"�R�8;�21�R��>�DÏ;�Z�ĺ��;�\r��d�7�,+`!+V4R�Z9��nBt���D�D:�[�~<�M�g���\��$D8$�J�d٤�W�1 ����0E��n���_�?�GH� �ғ�1�n^��=Q1�`���}mnr�70�!�F���JaƇe֛�|�o�܏��>�>�tڵ���� � Ld�+�$���Z���r�H���/� pCW.Km��m=n,hs�0�0�h�۸Q9�ʍU�A���3o����p�B�;0#h�{F>��R!+��+ɉ�,wO̊�!�J���8��rK�-�y�~ՙCͼ?#�U�^���:cކ�n�w
�= D��'�X��@$F�M1�?�L���Z���0�CdB�v���:�t�ܘ^��)��i�.%��-�/6�?���°Tu���ic���j�9�҈W�f֨Uʹ)�v���I�Ε�tb����1�tH>�L[N��7����H;|�c�+=�lf�<�\]6!��k�`f4�zL(���-�R�&�u	�B�<1���q���=z�-�]8�ƈ$Y�0H�I�U��3�G�Z\S"*�5nBr��c����k�M5qb�4|W΢����#�p�t�X�J����D���d��b*u���ړ"8�[�!*PWK��q�"lH��WjI�?����d5"��e��}?�/�^��|�جOa��2������gR��%��ë�"PI=���)��̗Y�^��d2��c�;�x7E�C��M��peMV�UW�����%/���֔��_U���TS⯨Młs��=q���ɿ�ϭO�Fخr�Jp��n�p{�0�����'��eil��a�l�z��?�Pj�|��M͈�ZeJ�B�(|މJ��D�T�OtpTiƲ�r ~�[��� ݃���!oG"��c<Y��l�d�&n ������
�M���:��8��R�z���e��s�18C��>n�X��s��mhǗ���G�?ll�5�B�/�M�C�,j���W�����r傛�"Mѐ���Rw@.
;�D�B���e0?��j1�� T"���oA@�qv�+p�8,zi�P�%����у��zl��k�����<o]�:��T�Q����VXg�ί]W�W�@f:��%.����Fo	|%�~���:�
�%�����.�:7�.�?�A	��7s�N	+�cwG�����N���4򃫮�.Rz��E?c�~�M��#!��kUndғ&�F�\I3��Z��Ze�7��2\)Cu�q7��I5����7m�d�GIA@�J;?F�Tw؄��<���*J�q���z�6X0�g�����ǔ�Y��T�KD��U�lB,e(֐�4�L�[1
8�[��j��G]"��Y�����������`+����M�G���&+�T^giH�K���������)X�G��͍���8��Ю�!ȥ�w	tv�kzsM�[+^!xq�@yy��M��qL��u�#�/��@� �������Sq��G��57x	v&�MH�#M�Y�f����ݠ0\�]�36F��⍴�tX֬Ex���-1���{�6H�8�	��h��ǥ�nh�����+AR��I����e���Md!���r�|$�r�L�]��Cta1ypUd6��s�+��ʞu�&��3��S�O���
{t�,��ɗ[�ö�]}v�M��쩞��Qz�5!HN�/�x����D�ɺ�@�s���2k��o�@/�5���L� �ɔ�V~�Xs���Wz�JH���g���)��V�y�uZ�8�Wn�\�(Y��@rS�)9#�=��q3?͡���`q�S?(�X�>:S���%Y�|mAM/���b&Q���|��%�mg��9������B���hݔP��[�A&^2�������`n�ă�{R����F�`�>��&,NY�*�ݠ9d���Zl�<i:mk~p�ET��y�o���OЦ+M�3!o*�\�ٕ��f�,n��33U߻�3︁3(��6~�M����I2�Z��g�\����|���;R��B�i�%��<��ph�;pq�sX^(�P`��7MfTx����Ҵ$��vsd�w���� �86���A~�?��߽�	��7�I��,_�Z��A�!B������KJ}����:Ow5-��R�UJ��ލv< �k���h+e@�b��%�%^F�^6����0C�^�k�g0V�����������!S�"}(K�y��{e��@�[T%0�҂������'ZȱR�A;�>�)��E^�F>r?V��҅�$đ�-�z��w}�n