��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2��@l$�Ndy>e�p���,� ��%�x`�4�W��!��:���������uH?-L����,A��iFR�!�ê2���1��";Ɯ�p�6�3�����n���۱$t��\MR�Kr�{Yc-б�{g.�����K�!+��<���)_f�Y�H�{t�E���-�?����o�\�g�Eѣ�T��ד�*��I2�N���!~�u��g[���|S!]j���Q���N(���i+�X(��z��@-6��!�PIVZ::�u��ډ��G$�!U$D����ӕ&m��JK���͖�.���N�'������5�4^&��L�JZz���*k����I3��_��(��.[�}�ϯ�K�h��axA�n�Kr��';�'vp]hT�I���bb�a�0�y#�1 ��8����w���^T�Lu����W�6�͚E�E������� `�{L�F����Ƅ6����$��7G$�9�� �mt��۲�������+��Ywy��ڞ2� ���V�;adx>��!�8H��X9��5�����k�eJ6iW_��q��ͽf�2��ɂ-NQ�g���L�n&z�Ht�\�L�������Y;�/:KqWW�X-^�&�G�����\D�RA��G"G�����BF�������V��!�_0�	ۣ�}۲I0�ܕR��A�Z�؂*	m�4yk�Zƈyh� ?S�/��#!���������iE������
������4p��%�Rf��~+ȇ��+�y?Xi��n׾��Qԓ���┝��+Q�E���'���-bl*��2DYra�/F���P�r�	��������FU�-�2	ג ڷ�,&>j?:P?�Y,I�r��g�B��!�~��}!7�z�:����J�Ƌ���P��쓱#6hF�E:B+�D�1�,���cX�O�[H!=d�6�����R������P��6X���[��f�5�'W�ᴓ��_�?0W��|�7W8���֢��Ϙ�(�ћf�X`Mۘ1*�62� ���0�x��_���6k�g��7�A"4������4�{M��ўq����Kg�O���!15)�+"��Ф���|��9�m(]J�qYd_�`M11"�I�L9�ck�g�Cci:]2��YT�Bh��>�~  �;zƾ���+C�8d����	֖�1�g��̱�Eb`^)v�?�v���k6�3���춧#_9�pJ.�*�HlO���MQ#��ro(綆�9��RG�����=����ʯh ��*��g����øH�_�Æ��6�r�$}��"��}�����&il �e�O�N�����S��jb�-Q^�	��j�*h��̮
�=��~�G)� c�X��������bt Lln�ҥAc��`��!�TV�����S@�(�3��*�Q�Q�F ��*��"��}C���1˺Pu��S��n�V(�3z+J�l*��E=)>�@�͜���Z��f�}��3N4/��D�[����q�<�tʹ�\�5�d�i�0Ƅ���/�+�#]����U�D`�-��eo��&��T�c�`	J
_[76Uu`�aU
o��mO�w'�2c)Z�,�-/s*���{Hr��o��V��̴A[���"ĀF*��i�ܟ�͏̄�P�V�� �\9��#���?���CB�~:�LQ5��ͅ����P�ز��2�{x����
E�$s��3��/�Oa!%:(s%��)�y�p챁�ݚ�r �:o~W�r��M����@��������8�������C�E��`��ր��!���j�k`�zX7B�x�M� /Y��P>x�0��S%���_����uw�HM�v�3	������*NSt�o���~*T�ǧ�H�"q�w7���wR����3��)}鉣Jӭ2�z|5�$��;��5o�������v�A�u���t�o���I�"D+�/�B�7������U�t��*uLi��>����.§a'5���d��ס�<�bv�Sճ��6��F�iS��Vk�0�{��<��W+�|t(��k�^4̤��O�,a.W�U]u�q"A�^ʷ*�K
��r�$}mFR�i��ס��z$�^�\���
ٱ� ����4�zu|Il$��y�tU/B�J�g�N�	�_#�I�a�/����*쾦W��v-t(��P�b�po�F���^.C�h�E㆛I�#�0�aJK?F��O�E��0_ή m�Vq���lw�?*_	0�Ʒ~.O��U��`£	�j�vM˷Q댱��K,#�xaB�Ta�2��筺���?*p<]J5$�U�lBs�{��;��]�.��-z�V��A�;�6�q����<��8\(-����{�?�d��.(��'i	1��l�ۯ���o�۬�T�P�v�x�X���+����j�����i��=�Ew
]�{w�RwG��К�:w���hZ��F�#}HGiK�;�(��ރ�8��D�,��ޫG�_Gy.������56ɔ�$�b�u���ԍbZ>�v�d)��XEOu�@2sZ�HO_NP
�&1^'���%L~��TzIE)P�����#y ujo�ŉ ��h��V�w �[~����$-
ܼ�9���E�?,��8�\I�f�d��d�,{x��@���I�;���M�z�%��"���nņ��y�D!�9o�<ٓ@+�W�0�n�'}�9����O��4Rz��r�@� ~��&�3�9̋�g2���i�ݞ��=&`tO.d,�~G`Ơf���Ս˦zR���z��J�y#gl[G9og�P^/WZ�¯$�6o�0��_���d�nY�Yhu>�JoRbU	�3U�x"�U��Qӳ������u#�D�S�E���&"6�����4�u�a.�L�_j91e��"�
pXaF����m������J�@���];��|N��ᤒ�_���B�W�^�������A� z��׆���\)^q����<h�c�bEm{��֢b?5*h[e%pl�e�'�M����M~��,���v	̝t� �����0l���U���s��� ���4��zpϯ�F��Hĸ���bCi\�X�:��[���.4���/�bőR�7;Z�,����<t̐�5�>�%�3Ƌ$5�5� ��3*��̎p�M����z�����SQzv�琨zt��qP��r���*��4k~|��KK�3�8��{���'�4%G�G���u"E���n`�u�/ݸ���g♥b�H��q(DfG��J �3z�`A9@>�f}V���́�jc�X=<9`��@_6�#��	b�"q�]�30p�6[�4JW��CY#����B+�9.��
Z�̄8KDܫ\����%'cAC4� ��b��T�jC��w��4�<�m�h����RZ<q��^@oXN�ѳ`�<[7���o~����ܡ>� K�8`��d���paY��dʎU�ZF��q��-����WXUm��|5�'�AZ� L�Jk_�6����l�J�
k���Cb���X���댁���ܦ��#�x[;�Dbv�@�zm��Ņ��.��5q�q��D�n}�IZ�����x�]���,aގ^cʬMN��N��F?=��c�F���ˋVg�I��Xl��`&>�����H���;�/rU��.��MOsV��aĺJ<m���M�"�tv���ċې�]C�)El���i_����薼�ꉼ�_��v@)ʰzm ��8:M���X�l�"�k�*#,jQ���B�x8۷uc"��8wB/^.�2�U��X2�?��ග����,<$��ȩ���d�GV��*Ɂ4�PT_ݿtO&�sǫT��,�6=��&�ي]��X��&��(�_ ��5,7bX3d]��tz�`{|.(��}cy��<F��S��c����Du܌z�x,L�����?$w�����8���(}jyڠ0��:[�S=�r�d9f�t�����Ԅ�[��1	h�5��kTf:�N=(�'���Z���W�Xt��9��L�z�0
���+�Y�{.R�ƚh��5Q����۰::��Ԭ?�Lqz��H��搃����|���*�t��=�Y;F�G���y	p�))\X�*�, ���}`���1H;^�6���Wd�Ǘ�k֑����>���G�{�����P�1�cL�h���jP#�3�%�A�d\4N_��w��g�*��LN���S
}�<��fݘR�}�h"Ґ����h"�-����"�2N�NgE�}`��ԅ~ɚє�>�����5���'%L!�8���(���� vfH94fE�>S�`�H��9g.��sA>iɷ`<�ːz���d@�q�2F)�PU�u�YkFji�0+�`�б\K5P�߿_!�q"�3i;���Zo��si���kg�y��D����=o%�E/��-KMGU�H�a�v
P����
�t�U�� ����m���A�0�i�?Jo�sg�㈍�a����.{�t;)�����G��SW~�D/}o6	�")�<�=pKP�lS癕���'xT��j��H'A��7d@1�W��Ab�y�uD��c�RC K�CQ��C�1�t��K��yeK�u�7�Z\�O,㨐�>v�S��ӑ�{�!ƺ@$�D�`r��4�b�|ɓ�(%��4�r��A�d"��,��1��Z��u*j�&�
���?q��M|�|,w�"���@��=,���B�A^z��u6X�:�Z��^e3�#C�ǹp�f�+���M�w��>�G_,�9 �-��?���,�-XS�?����Y�r��}<�M�V�e�68��:�Ă�!�A`�A���B֍�Oh��C�a��vN�q �}�?�!�g���#�U�E��Pļ��@��6f������|���d	�,����s}ѣ�79v� U�>]Y=	i����g�h����%�yE��J��E��4Q:\��E�Xߑ�a`$.lt�_�%�_L�o��N�
�K}�3�?�IOu	U�.���]&o���NT�Y�����-I��#C���>����p�w� ���Ñ��:�ec(.qi��1��\u��-K[+&�x/.`�3<x@��Eo��?a(!�}61��]*WE�E�����g��N3�x�Q��aά��bGWk���l�S���_���-�"�qi�l1��z]��PC�o�����C7&���(Mz������R�� G�P8����p��1�2�DS�n|�����ֆ���]�ǽ��<��d�m�C+�F��ST�~�*^��sqLxw^Gvs4�fJ�R�`��a}Μ�V�в�ĲZկd͓��)��<�:����s�p �qc�Ǟ{x[�3F�3�CnU��~h+C���ӻǽ�6_ʵ,� x�ŰJ��#�s���יBhg�!C�;a�^�݂��aS�&�S��!vj�3ݢ�'�H�̢rR%���[�)�=�ѝ�1i���bX[d9"e5�EX�G[���m�g-�K)\�,�s܉��~��B�S�0�uS㜙4"ɦ�yb������5B]糼��(Jm��_m�|X�=o��d�% �fɌYNgv���w�_��T{�\�^ ��<l�M���� �?�Bh)�$�!]�&��s-U��! bP��N��b��ݢ� %rQ�Fh���O����gM��қ�ŧT��>��B�s�-f�U����K�����lҰ/`�&ooRU�rU�"S��HS��~�Ƥ��zi;*:q��L�ΐ4A��)V�#�'y�?�����8SC�%<=$�s��hb��-��r��Qg+-�EkPh������
�^b(������h�kk+���OgMӿ`�
���.�N�Tr.�7���@<��F����e����s�|uT�w�30�!#e�\�W�a.
�'@Z�5ma?���R�0JkԳN`?4�!�	"ՖjRx($�&��%y�M~r���>�����.F������?���#��ZW]I�(�d���+�����N1��SU��> *h?5(�צ�-���'i��Wr�0�g*.?wU�?�.����v;�������?��s���{�M��<p]���/�z]Է1V�M��iш�0��<&�1ɕ�R��	a�M�Z�����I�A7�vGJ�F�:�cƶ���]�!�� -JA��:�Sc�9\(�1,?�^p O-����P��+@��o�ۍ��+U��Z#�'�L)�-�~���1TY�,��IʣZ���k�M�!A�]P���ݗ*y!XQ�9�e'bKJc:�eIy�µ�H�zsJ% �CZsU�9�c��Ŀ���ˁw�,W�k�BȉV�|�bh��|m�k�f����g��*���oj�E���b���D��Gm(�s/�b�N`<DY��~��pк	@�����45v�m_5H{��T���9�ol���v�0��3�4(������X��Y���.�H�R_������\]Ĩ|��r~[P�=D�9��u�dU�Zd(�|�D�X�m��:Mk!�o̹Nn��g�c�����֙o�E���([��V)�8�����(���|j���Q$a��h����ͣ�ap�Z/�햙~ۈ� �F9zy������tH��i��?o���Q����y�NF�}��̕��;�kz����"o�<Á��C�ΝJ��!G����7Hz���F1�a��6�|��/~�ܱl�jRfhF Ӧ�2`r�'��4���䰓kk�s�c5Dt�4�`Ѷ��U>���s!�����i��'(�46���Z'�⎣Olܾ!������y�e �.�ֲ�w��DR�w����O��ۿ��:���Y��=��Y<���韉
�-܉~=l�01���߾�g���B�"B��]ԫ)�q�Q�o�O}��n�:z���:D��2ls�JbV2�e>���ߘ��`�֍�įe	�c��Q��� 2	ѱJ� ճ.�%��a1��������4Ð��7!3'���YW;2YT��W�U�mK�=.%�^�<��b�{����P~���J
�~sbdX�4�58���%U�fug�ҦE;(��C�R�a�vvk8/�ŽblZ�n2�%&����O��p��@��X�Tr���_J�?��h�q�x�ʏ���8?�r=�Z�Z�>:�j�l^��>ѽ+����� 9�M�~�k,1���e���4��`{=b��?��g�R���Y*0p��[��jvV�d�r��\Iw%���r�Q ��E/�9��H똡z��3�$�QR�m�N��r�8j(���-�K���D�W�nM��Im�%�MH+�C�o"|�hX�9�	|�_2��7�*@���i{va����2Vp�����ƱO�ON��aWZ�+�?|$w<�]f���>+f�s�?��!��#� ���n��v.�e�L��k�;o�S��c{<�ՐJ�jǾ�J���&(A_]KNJ�d�s����(�^�4��n�> [A�81(6�%��(����Z"�&n+ �)��k�+޼��";�f��R������gS҄xR����	�!\�<"J�_�CN'�����$i�|��J�!M�q�9��07M䴔8*�NS�����5C$�������R�����2�Qj�#�^6��Gк�{����&ݶ�� �0(Z�Z��֫6��%}��h�Q0�B ����4 I���C!m�?�.bB����_��Z��s�a^�MpB�ⱀ�"qi#k�\��I�c���z���7e�t�uP?C�kFGb@u��n"�D��AF6�dOm�>,Ic��@dK����o�4����df��~a��F�Am��ҫ������t���f�]�1@�Hc��S�?!�Ѕ��B���<!������qyId��h{&t��6:��43�E� Z�?u����Ζ�q\?{�w�<�
?+B��&�!�8�#�<�:����lM���0�7J�7��!��#J}��}r�V�)����z�c�J?�^H:Μ�x���P���1h��ۚ'>�:!��b��Tȃ�:�=CeUO�搫֞�����Y��L*V�_6,�Ѿ�vg�rBXS���:�3s�G�к(�֦�T��������a�s�"�?/b2V�]��1v)é&U�}'R%k|8,ּb�V�5B%�{:�5��P�n>��ErLH%/�Z��p�n� {t����Tt�O��%��X_� F��W�v�N$=
���+�g��<�I��%;:�n�!d"��\Y|�bI�[8�i��穗���z=�:���wM�)��l�~P;��> ��`^[�`��k�����u����	=�	��SҎ�|��%����G��	H����]�X#t
aȡ�)5*�S���6v�H/f;/����� l�`��b�Z�U�ȳ�x�{iX������`.\H`#���|R�'�W��S���n�w��7�<�i*/m˼[U
XU�<�N�-<\t���q u0v��I�4��p��a@�˒*��d�jث�Q"I�/V�Pj�٪�:ב
A�U��5(�1�����8M�&���p���H*xGN���_S�8��0�`�*�]���o��M/8�_o\ 5/��e�QLCJ���������� u2Ǒ�_�SS��net2<���W�&q.��s����@�L��2���#��t�fO}�� �[L(x���{�q���䏟�W%q�R��R-+ϫ��T�����/��M��d���C�ۻ7��)-��j����z�:���$�Uܦ3�I��أ��-Uѣ�M�o���A��p���x����&�XC�p�ƥ, ��� 5��?\�*@xha�Q[v�d�ߥX��r[*���4��N��si��2Z~��c����3Z �zͪ����.��}]_��}�g���e�y����*|5Sz��}��5|Lo,�!�Aa��KZ�B�S��G��6q�n��=�%���צ�u1$�T.-:cZ����ݨ���	��N��L:C�Q\0G����a�)��\R:7��>���70{��t={<� C�r>ū,k-:��V�:�˟�	t[�#;b˜�= ���j}6r��+�\����%�-I*������5�f�� �-��/� ����[��e(�E�f�Trq�wq���sf:ٷ�k�E}�~ �.�3W�O/f��f���9*
Q����b�?�Ċ�p#ӿ#i7?����vhf��"��(j�[G�I�2������G�*�	�GjV��]�<�TC1V�^�m�a��r��ã�,�3��K�?�c$jV��/x�Q��{���xs���ȵ����?Z�U�*R�l2���H��P�v�&��˹� �9�2%v�W�c)�8-�Z\�2��Ǉ3I)�LS�
h��[E�5�++���r�*)NJr}��"b�}y�N��2@�Mu7����k��<+��@�����۠x�����wC�-��w�˨�����e:��_��!4@x���y�X��B�3���ib�HO�C^W�!Q!��\�4F%�bH�[Z3N��q.C���aw��	�;�����g��R�2�Y�"s��V?'��T'�b��p�l��3	[fm�]p(񂎫Ԣ������=�{���.�W�HL��G�1
N#����`*jÊ��V��ɣb�w�;�͟#kvgi�{O�Ƴ�0��?�%d�d2t
�Qe�k�Nue��!���Uwz<�/�qϛDVd��$���ō�@Q�0�.Ig�v�=����د�N�3���Պ�W
>�\��j��d�pq��֮r�S�-9�'Et�2���<E+����]T�ش�'�>U2�[ɿ<�D���{i9w�+D�^��>}��d�=r�QA*#���/�t����\4�S����6�1['R"�Rg�x2<�]����/��,���3Rb+`Й�����Mp�D�7�W�I�p��D�*] ��y�;�GE��<.ɨ)]��Qj�Ǭ����/����#�=d>�Ar������+VƼK�o�����ʦ:ȳM�!��8t͞<ߐ
��dwY���m��۱��!�)��D!�1Q)1���ܛM���]K�9�XW��v7 ��m28ݘ�)��&+#��v��1�r�
U*Hl~s�Z�_ho=����!�{û����=vYv��g��(I.w�\�A�|��#mUQ�OqC��5�0�VŁV��_E��6�R�K�h���^��=m5�E�����y�I�F,���S�)Bq �*�-r8�j|_���"5�����@;P��Ŕ]|HT�����ƸUi1/�T���?�N�����f�P�1���\`�Q�?�n�Q�|�U�U��w�.k4���Ӻ��o �;��P[B~ɅR�f>���w_Ӛ�� ���ULN��%����y�J��!��D�lo��(�0��I���d��#��qW���|u;!�Ak�x �^�V�'#�����;71]v���"�ٝ�=K�)��N��)mS;�.��v�V�i����j{�2B���]=��I���z�lD�4p�	�<��Z!X�GwrI^:���l��wr�/w�c�5'�����y?I9���b`�uBUA^����UMg�ѣ /������t�I}����B�M��q��N��<Q*����[Y�c��6��L��&ǁ �pJ6���
z���D���ՆO����A��g�E�~d�%�F-��t�+j�G�z,<=�i~$,0�J�ba��e�͉�� i��X���e��j�DT�,W�4�6�{��w�~�a��_cW���Eh�	*��~]^Xb�Y$���+��ѧ�Y'�uuN�����	�Ӵ6b�w_u[�5ڪ��m'>đ�`�]�y؂ �:(����R��&`�i��-2�Y�O#U�~!5}���!�DmY휒�x��0��>K����2�mʀ�����<���;��ʥ_)�NO8��ˍ��>ym��y���X�B��EM�V��ߚS�Y7?����_-[�7jS��;��U�5k 	L�Dd'Mo��d��^�)"S��\p�g��p�Bcv1]�!(QqT�tփ�~ �E���u~������ 
�4�(0i�U59#|Ը�1��R�s��~�9C�~�)���X�zb�Umf}^�n�n����LS�����րi����2j�c�<�Ph,X�"z��W�.L�dV?R{^;ށ���]��5;����Ư�7 �BB4.�\��Ў�kE��p��n�
�T�����W��˪,C<�F��|���4��M=9ϥM"F����."ae~�ȗ\F��G�C���-
�����<�3J�j��隭R��[�`�bY$���^0�F�3��w���RԠ��g:Ē���/��
b�Õ��1V�}����y�3 r�/��]xNj0E����TF��g���g�ދ���5s9|��y͍Xc$�D�t���u+:1���Ź'o��*�i��1	�����+$ɒh���5�����`�47�j�hԳ�{;׆C�fܳ��`������4�}w]�]��镥f��T�'seZV톫%`Z�f�D��<W��׭��seפ�]<ޑ��z�6�b-F5�y.�TϹqG�G+� ̜B�4?�~����H��Ѱۙ����91R�k�D�)g��ME����~��0�4~��a;Q�;�52��,���3	�"�J��S6=[x!��x>/Tmgb�嫀Sm�3�*� �4RV��Ȏ��N�6�ߧ"D���$���S�<�F��Y�ɵgAjX?N�R2�f�ԯ��6@I�����x���I�4�ѡM�9
|�k� �=Ȕ�T�	�)�Ȣ�v1�,;������z{�;&��,��N�e5x��!O���I����Ɲ�O�av�G�+(����6��O��U��^�STAw`�q6N�U�g���E��^vnlU��r��2�����B� ���g�B,;�}S� |�y�X��N�"#j@
l����`����Pzw��}~#!N�����K˫_��������m�5Ť ���5��QGZ�"�Q���d���(�4
��|׻k���3����������k ��6�k���p�ޛ��N:�����iO<P��K.A���p��]�ZC�\cU���J�[�\���Ky���=3�a�A^��ͼ��pz��,���aG%��fy�X�̷������d�	 N0�"D���&UqS����'�m0�x4�	ؙ-��,�c^�[��ͯu��+�UV�N�Z��/��{!��j3qX6$\/9��t6�Ħ���-y�%�αW~"5?�<��퐊B6�?�� y� #��a�� �'�%GA���d�C��⩮��k2�&���yM��ei{�����j����t�0Y�pbA�R�xtw�ڃ+V��~��Z4���U1��) 㵾t@0�z�����2����췈�=l;�<���o�8y7�N��?@ԓAKXÇ>6Ͽ��C�2Ƕ:���V��	d��k`���#E�G���ޚ�0R��#F_'wn�YEB�@f�P�*S�|h実���	�=	t	�(�HU���4�Ɛ��GL���"
}�g�f�5�sl��:�i���L{�oo�!��ւ�Y|���\�����2��CJ�����+�@Ƥ�'PVOAϯ��Z �V|2�
��8c��^оj��4�O���U
Y�c���_����%ep���Z���^;%�/��y�{�4��]5�S�[$���J�ߚљH��:�q�"�vA
��t �˘�Kߓ�F���#m6�q�IXx�����t�7�_�͕0��P=7��5 �)a�ARq�؛����w�;�������)9��G�f���v������xr���}�i\X�Q�h��2 �tR�~F�2��j�W�֪B�y$����w:�u5�t������/|�>�[�?�@5t��T��EA/r����Œ�V��ZqӅ=1b�X�fp�t��
5xNAs�S�ZM9YH:~�����������
�1I�<@��>u|�>[S'���)�%9R�lg4�F
�{���0pw�i��q%<�����6����	D"�˓�\pA;��u?����
"��`��c�C���MgG>�w��K���sĿa�y��im�xn\Sԋ�(�,VyǡeCθ���T�c��ѝ�Z��5�#�߭�:_�y)
��7uʙ������=Y߲K1�h�(�dX��v>I��G�D۰�X\�2�K�#��
� tN��yEWi��`FVB"��K|tz���e7X0?'�BX�h! ��з"2���=��X�fvw�[Ƚ�/]3?�{���7ݺ�iq��vo�q~)�A�Ha��㵆Ѥ�7�lg;��U�r\w������V~Qn�,xMq<�3jy��vti�߁���æ�p��yX�,R���*t������l�3��I�%�R�_��],/�B�Dq��'�sL݁8$ܒ'�̊�N5nIe�ʼAi��������O�O�ߌ\��lJo�<��N���x=�ϰ����Rr�������j���`��zXDO��,�����Dj�y2���-��1����a�)z#�Z��-�[�a��euK���j�of8N��s�`�H[�/Q��L=�݁l8�=L���c�~y��Ȥg��$�J���#����N>YWt�9��:y4?����G�Z�x18C�*��\'����/cx՘3��������TsI��ϫ��ҫ��^�6�����h�� �9��;W��,	k�ɒ$NQYA�_�5�s�zq�O^%���'��e����E2!�}���;�VZ�-��� ��>�ـ��S��@>b���ַ��d%%�D���J�`k@ݡ�c��*��Ѽ��YF�7G2)oޱ1_t0+�s�,bbB^O���l좋#��@��aT�[b�S��������̵Щs`�2/u�W�Ur*a��g�2ƞ
K���1O�VbQ�22R�p�������j}d�%%���Ae:4��~-�+�If���#`|�[4�-���,����*�L,[n�?�,쑛�r5�EE]�OF����t�c�+uc��9��@gjtB�	��״���e�K�0��DJ��K.��l [o����&<��$�����r��2�Z���[�)>�L��}K7ڲ3!�st!l9���RJZ9�*���]~��%���%	��A'3��Rղ'X.��L�Ɂ8>��X��.l?G���! ��뉶g�4.N�������C�[��%��/��&�iQ#r����
��Q���2R��y�����X��`YB�'�j$�n����n�*C�*�'B�W&V����*�\�!f�{S�74��SȄ7�J���DZ|�űR98s:f9]���a$���P�~���>y��'A��P����ꓟc-}�
,$�IG�A����=�<V��睮>��_DͦIn��D�>��Le��"���oɠvq�N%�c0EԂ���/.\z��r|,8���&�:Q�缦���F�/D��=>���4n�/����I*]�"��F������B1� e�a�7кA;SPlnˤ�@6t��;s�z�����3<z���Tꡉk����K 	\=I���I���j���VGj��>�?��|ޖ���cXYq}���o��îi��GZ��k�y�5o�3j�d<�#��n$�̾˖N.r����<,s�QSz��Y�Q��":"��	}�1���4�	A�g�j76�Y���X-�VH�#n��|�Yk{5;̲}��_�l#>L�K6Ƶ4���Y?ި�*�"C�ƶ�ΰ��U�����
�9�y���5»tw?ɺ�����{������pI�L�"#�#f5h��A�!����˞̦�*����I�~�|��}��V]w�udz�����_�]���T(��
��}�v�������Ѽǽ�q)����5w�`]h��D>5����.2���5_g���\���x���D���H �#t'������m��g\�w��ʘջpi#��?;ɜ��=����U\e�.(�q����o������1�]���d�?�J��K-,�D�M�)��A*Q<JE
|�jr<�f��k�tD�fP-4s	|�8=Ȋ�x���y=�j�k���4���ۆB�M��JUk�����X�ES�u�O��ʑ�@8��bN-g����>ڻn���ng�\���l��g��M���cAz���C�rv=򃳿�'���zZ
���؋Ug%�bR�=�u>�����{��s�����m�+��ۏ�P���t�����/�Ί(7��)/ª:�ý7�fC���ZB^|M�p��x��.2Lc%L���ِ?�F�)/�!l�j	 ��ԅL�g`:�}ŋ�r�O��3J�m��P��ZvB��ϥP���R!?�oj��AC\�ٻTw��?��^�ķ�FTT�<�7ʴ�R�e�|���^+FP�0㻀`i< l��̊zv��I��}9�dDJ4�(�EE�ȅ8H��<��hR(�tf� ����3�6Ƕ���@.��D�!i��������4�"�Ma,��8����������Ձ5,rr^�MHИ֋1��M�Ȩְ���g��/��8;[�\猳�lK��c��.)d�����JZaq˺P*jHq�:zM5�I�iJ����V�`e=,����jVB��o�kM�ׂ���.�f�&EGj=�%:�P>¢�R#S�r�WN���O�ڙ����%bl#�N%�6gl�?��O�����{;�W�QG�;�3t�5U{�vk��Y�)Eh
��]�ѽT9'@ͺ�{*��W�I^��V������3�5E����<_�է	C�ɂ����mluە} /��b?�"��_DL�:��5�F�ηuJ��)�f�� [D�s�*V^�D�|E�(�-�Ri��w!�5�(P�{��
��Ύ�2��wI�S��aI���F4���>�Oe��`G4�C���+^dp�y���#��Wo�x�:&���>l�![Ӎ����ݱ������k��쿰G�ED,��K�n��dvl�e���v���4"����5u9��F�M''N`ļ��$T��zѾ��ylY���f�$�4\�`>��i}��W��Y�J</�C@�����!�aa��}Ii4��Cx�a�|O���)yFwL՟��hO׏*&V�c�{ |���G���hYw[�r&(up���]�>]R��.���Ĭ�=���Gey#�<�O-v���� �����"{�jl��k1�h᳻d��Ի��[Lw�l�ƢA�G��U���t��eI��7�� �;�_y �����l7e�M���x���_т���ه���N�]c#My��f��G�o@՗n[�]�����/+�ڵW�-ϧS�,�z
F��e�GiZwq&�XCD�˝�7Y^��:��!EA%�*jh�ޞ�_9X�(P�)E���t�oGd�zt������Wha�����;�7�u>-�7m�.��ڛ$���"���<�;0ޅ�9��t=�(�ڡǀ�,��Q�ⵦ^c�կ�������,��X�~��2ʴ���lY`�x剑������OI�?��-&��qsc,��T��ҕ~��U��f�+