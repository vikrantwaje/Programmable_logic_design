��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2�ǣ_4�^ZB�}� ��1��g�	�Զ�Z�;?h���4O%��	��J��2ө<��������sn�،�˧���}�;5�y/._dvv�C+����;�v�� ���dk��h����Lw�y��\��n5X�t�#���<��Z9�;lH�w̎=��	���� �p��ĳ`[������ ,�gޏ��Wհ-�6v�5�$��Χ_����_!�rp3�'e�퉦�B��Q�p]>���ܾ+�
��h�ο]�X���t�@M+�5�p[-h<�"�V����%D�u=�,�@�'��m@��t�P�0d���B���٘\�m	���S��,��p��Khљ��W��g�f$�#�+�<����[���B�cݽs�Dj1�>O���<�k�E��(� �����dd]����wG�8uJv�i��ho_O��"��Cg�L�0��1������GS?$�a��`er�Kɷg,}Ey/���h#ǰ'�=E�l����(yH��NJC�Y�2��+u�kdx�@m��`��D�ݰٌ�c@$_lu�ă�Sb)w��&j;�G��9y�܊T�������{|F�\[yyͬ����� �P(�x(>�9��
��$�w��sƖ�����Ď^P9�VI�	%b�VV�?�|���\R.�����ؚ�b-r��GL�f֭R��V�t4�7���WDn(<��F��]�|o���=�_��o6�K�m:�噛(�&�>��;��d�ϒ�N���`����FAc�b�(wKxD��*�S��ֈ��T�-G�ƨ�=�*1��h�xU����� tAZԴ�25JB9���>80�t��#�sl����h1��ɍ�m^5��
��y��rC�L&�������M�����}W�|���
2/�^�J�1Ny�S���Jr�U�@���duu;����G�����M�}�^����FB��ma�g5��܍#�u~��r�v� �;��+��X~n�PN�P�et��WV���������]��;�R���BMY�[<��B0�e��+@H�Ol�� ub�q�O%��=�ڵ��X��3?�^O
%����(�33�)�;8�%D� 5��
.vȳ�m��6�e�f�����25��}��n��Z���jP����8�po�rƉ���X
�C;ĤJiѦ������]I#��%	�: ȓU�	�@#�@=�lp[�2�m��?�Ѯ`�{��r ���u:���d4{��q.0m�F[k�"�=Ǳ���G�I��IJ�ᤎbt	�at�Q�J]\�"�e%D�������j��J�@�f���>"{Dn^��JB�۷ݴ�Mk.���&^b��Qj�̢� j�����lv�g@�P��\7n�d��ѷ�&�6���!�,�U��%!ȟ�s�i�_�F&K����C��5&�y��}�sI�1�Ji��̴,�`@�����j�"���E.�j�r6s�>���3��$�RH1$�j�C�6���\��0��7��.ǡ��h�!��(̵щ>�޲� T{��̗^/���Dl��J���"4ҕ�$�Ę�����R0:C��� e��Gv�V|��v��>)���`h���Tt]�Xl)mfz9~�S̃ɚ�6 9���r%�cDb&���"�}��z.����i��M�� 0���5���e%�\o�����ڿ'���#	������_F�̖���~i���l�Q�Z��VbI̰��3`�$4�q�[+C� 	[*ҹ�f����&�;H��g?x�.�8bH!~*�I�c�װ�zf6�=+��`Eg�83��}�߻ق2[�	�e�B��c�����j��V���]�6��W��c*J���+�(?�ضd�/�u�l�]��S$����C$A,boYV%�E���u�Yo�ho���o�t)U�Nn9�S	_J�w�w ��H0�3}2J�j��2��LתxoӶ!��f��\BG��ӄk1�Ә!FAx{��D��ds�������X��`�{����ZT�AZ��h\���LyՑv�sM�+َo�CN��M�Ei�����������,=p�
8?��</Y6�TqQ69�t��V��oL�[�{(� կGlϲ�P/�]>Ԡ����BC X��՜%�I/�ƎH���ea�����uY�Af:�F8�3�4�n ��.a�{Lf'Ʀ�S�ܝ�����t���-\_j�0{�Ǹ9�߂ ��hp�p� $���p��7��d��b�V�Zf&�/���x!ڂ*Q;S~��j����n?-r�m�EA�t��d��~q]
��k�D�4���1Ci-
(Jy,�1zyMn������MV�R3� �r�@p��?��0�H����D��P����81�қ�=�����1�F�Ģ@�����U���u���(]]�}q�1�D���i����g����Ȃ��G���ja&