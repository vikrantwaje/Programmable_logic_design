��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�nU%��l�F�y��7�R9e7���}��3�)Nп?�j?+ t2���|��T�Y����Ũ����Mp$����Q�3əxq:��/�He��h�8�fT�H2���[Թ�0c
z�9E$���Q�](��P�!л_ gݽ&b%}Vd�$�O �����FX�Ofb	 ���5��G��r>��T�CF�I�&������y�C�)��QNF����4��'Qj�x_`�'օͰ�x\�����~�;��˄lB����8�Ѳ�RNrB&���uS���o��w�!|
:ϻ��G'S��.��Hk��+*��Y�wsuGF@�˜����C�|_�������;��懓ˑ�7f0����D��(�.x����J���<��϶^1��ac��A�~YoȾ������r�Xl_V�ٜ_��1tڰ�"[�Q�`sպ@?�: ]�!c��k3�f�����!ȭ��p���<n�2�N}�o;�u�+��S�:�nHw�1C#l�.�j<Ϙ�'�jKø�ZH;��_��t�l� >FD�d�_���,���ح;�;��ǯ�"����ebe'�/���Z$��Hk�?=ŉZ;KZC(j ��9�	��v���~�o�yc��J0%��� �j�J���B��K�?[�m���5~J�oc6χ�WO�(t�Y�X׆��O�c��t�炲3p�"�� X0�8£�?e\v,���t�i&�~N���'����79#� �9�]��5z�ܣ�'_}k������:މK�E���,�M������ab'�\�L�ă�>��z�?ׂ��������C����R�;�lo�6�PX��b��y;S!�8��"N��S���R�U{���`�1��?E4:�X������R} z[�'(H��J_I�����S$�W��qz��8m��V<.W04�Y9$p���Y2�
����V>�ni²��{�|sǟ�7!��E�`a��V({	ա�4�i���IEJ�bY��}��sYS�X��%F��F���z�	G�Q��T�7�:ԸU4:(�����Ky�*{V�ʈkH� +)٩����%�@�E��z��y�U`Ѱl$��Ch���r)~|,��!J3�=-�YzA���=)�ރO��)�xR�����!T�ȸGݱ+fΎ���u�쌭P}T�Xc��n�y�;�AϦcx��;�n�J���8���F���:���GU�d� ��/��t�j��盥�K�^o5J �p����l��zm�%��ö����6��,���V���,*(;�Fg�e��1����C�xcF�(�.�G����S������r�?K����Gr	�F!)�jDW2�T�!��26����i|I�(��%�A�E.@�_f�?�J���U��(%�������ܦE<n��wJF��C����gu���޺���/��O���=ߕ(B~���U�a$�w���
�i:�0��]�*4j5��X�ͯb��T\��~�@p�� 
�a������lG���MUq�fM����I�A�q�n2x�C�-�_���v��ǳ�=���d!f���}0@5�X/��]���_O5���V|�S1��Հ����]��\a@R���V���)M�^8L���ͼ/��3�_�s����{���Bx�+s��I%܄˺��	��t�G�B�ԙf�ݬ1�����O<��1�����(��7�!�!�y�^��`��<�t�ō���%�ؤT����A�Xk>l���R�3!Z�yaEfZa�i�=��6\Q�:J�l��LQ�dyo�6�M5�Q�F���GU7����y��=� ��L���4sPZ�A���e�"�mRa�I�)�L5<:���zV�`$-�(�`�G�	"��yh$�����y���N�"ƛ���.��	��׋gTF��FI�5���@>�W�3�Gj>�
b��Lش?�*�pdZ��D��&+�އI�9"�kL�\�-H��:}���X��=)�I��>P�Ճ/���n0+��d4);-lv���;�a-����yX���$�&YǾ�W%[<btLK:��[��@�f�@Ļ������1���\����w��0�!x��$w8�UmD_$�/��]��L<͝D�6l�hEb[�D�pN��c�z�0y%q�slp��X/�o6���Q��
�N���%ӡܲa��)�'�In`ȾA�<�Rf�Ƚ~t�k�F�M;���qG�2��X��rI5@��kG�GDm��� �9F�n}P�E��(x��j�k�0�m�P���5~o��R�@�����K��@ɒ��:7Q��w���"�2�?��Փ6�$+���~�w�;�B�[n"l��Zo����_�Dz��a⤌�7ρ�
EG�Ҹ�Px���۳��~"¥�?4�a�;���'�+Ȝ�h��z/�<����`����Λ#���;�V�A@
��nEn��A��:�X0�8oE_���,����Ar�:!M�+1��Uw*�m�D~n�|%a���c78�ƌ_M����6���X�\����GcB�}���#��Yƿ�B^(��$�)���I��Թ��n�|'��Z�Λ�JF�ʤ��Y��G��h�S��?�W?.��8z�z@ݼJZ����)RTD3
%5ໞ����=��i���,��U���
j��vP�_d&�7����π� <g&6ޙ�Wѱ��@־_!4=�}�k��|���U��ז�B'�V_�ǥ4�ʷ�)K	�A��/�R{���*TH� �T��՝nQ�xq�2���1�O`��	)�8g�z-6}�)2�u�p^)�D,P�Ʉ.���H65z��=z$�� 0��ȩ1C�%V����Q��5�Z,M�@���I���8@(E���X���g���s��vl�g�b�����.�=�w�Y��g%LSo%�����W�7J���SY���b�DD��7u�}�,x��y�h$�w�-@�Hq
����9�4���<f��V<������,�-��J,�]J�rN�V��ǶB=N�~��R����?T˼K:g+��@2�fC�
Z��5/"��AϵG���F���'�$��,�/~��4�ᜍ�g��#��P���&A��;,�fJj��˞35Zϊ	�M����s&��b��}�c��d|�5�d����BѫșA��]��h�m�k��~w�Q�G��|A0��橫�1�Ӆ��(�lEs��&Ȏ�R-�&z{ACE�wx���2�%��=�P`�H�]!���R	�)(e��J��Qb9���f��ev6^�g�<5b�'�򇇠���p����������#���a����Bq�|UryОs��q��0E0}C����V� u�sH���Ղh�K_cm��ّ�����M��5x����3~�* �T0aK�����G�A�w��������%K`�&؋��y֯��U�ۥ��uL�#+��v�Y�{^����ڻ����wb@ [n.b}T�Q��}H�%�1��n;����eXa�I��N�(H�l�}�e�S$#�~�͋O\��	
,�����X��ۂ��H��τ�mU���86�%��2�d���g�g�q[�� �0!uO����h���֛(��A��Y&���F�!���/��m���r��S�N����G2n�ʸN��]\*�#>��S��eg�T���^3"�R�أ8Ӳ�gvIm�7����1��ļ�z"�( }��I�z��0qF�q���ɇO�E��^���.Asg�o�i杨���oA���Ӑ�����`CPIm��pl>��v#!4��A	�G�O���_�	w��Lx�Y�(�_r�z{�����Zr���䑊���6�h7���a��O�d���Q܁�n�@�C|�AR��e�'�}�Ϲ��Ч�
!�oM(���蚐.׆�`k�آ򋀙�Z���w�ݵ�U��5�a�Xn����c$�*v��K23{�k?B/\�de���l�ׇ�ʅ&|�녾���v�/^�<|M�xy���Ge9o�yD#�zdT�=�'��e�p��X�B.�	�`$1@Nj���lͼ��v���%0�]8��>R�?�1��į�^���gsm�Z+ƅ4��Z%�^;S+��D�<eڰ
��{і%<Ȋ��m�v	��"ƋmZ��{Ug M؊�qyT�1%�Ŷ��7/��x���<u:���k���6����R�!�ES����[��!��yC>���&ráG�S �e���9�����rI�m�m
	8Q��Q�c=*�G�M�d�Rm2s[��o����� 8F��V����Ʌvʚ����NWhL�뙵Wh-��_�|��;�L��K�wJ5�y3���A��2��d������`� �J*<똣���|eꆥ))r��z�������s<�N�2��Q�0��k�G�?�驢���In�� ��4~o�y���Ψ
-M�/?��̞�ǰ�In׌0��G�:jZ������/_Wۥ�E��Z�&p���PK�h���V�ݰ�.�l8R]�Fsƒd�����KO�y�=F�)��भ��o�;|M�c= Mfܵ�rF+��!�&´��x�-R�d�|�~�X]���<����!��GҪ7���IVV�t6q�Ho���g y�NI��Wo}�ݔ�#�]��Kr���[=�Gh�
fۧ�/7�m_��6��K}N,��r9��wl%�L��ɤ�iM�Iv.�+.�Ԙ�W%�Q�0;AV�eΫ�4v��{Tt�2~b-M7>���Ǫϱ�__���@r����eڦ-9e��ɺ�*�[�֚hy�.��wC(�Ïc�ڳ��Qg��6�K�$$��kMU�q���^�Z>9Jw���v��lD|�n�>������L��F��%Tk��{�,���k18�?����/��ń��:G'ji�y||+�
L�U;X�����,�1E�$��|׫�)�+_.1�_���f䉈�¡Ag�������B��![�Z��i�6)1D+GX_/�:�b���ճ�i�J�{�
W8�B�tG�}�\#0�=,�ˤ<�Q���Uc/��2��,�����iĕ
<���`�6����[$�U��Ir6g�r�Mo��Z�����AY���''`�&�q���xb����a�C�@����'J����igE�m�6���ܛ�����V�2�M�R5s�ƞ,H�$q�hT��l��\���
L��N�ܓ�v�1������U�L����T;{��"I%�ªz���;xO.���|�G�2(Y1�n�-���(������5Zx�M��"�۹m#��l��|�	�߱YM7,^���RD��F�_%큞$hsj_lUfC]��Hs|��Ƕb�#2a�j���[G99��s�`ì��W�S�Bǒ�ARO%R\$������X�u��	\��J�&��M>������uu�?�J�G|/HU�a��`���UnZ���1O�o� �n��(�7lީ�b��I7���l���A&��g�.e��a6���;TQ��D���J�aI]��x���a�F	�u��K^G1��"�N�%��O��,j�A�Ƥ��ǫ�k@�`
` �_M*��ė	��"��bp`r2�����q�k囥j��j SCn��m!)o���.�w@b)�h��t�k<�D�r�R"���MF(�c����(7:��Ͳ��+�ኸ�X�������O���X��4䔣���}"�ۡ@9�� ��M��,���x��Z���!�Ԝ����B��E����my�	�=7�����p�p����U�����Qq_�vF�p�@�=ۃ�[�=�Rs����ш�i�iLԹ�⑱��1�%������,9���.y"D8o�S��'mp�?'f����R;�������~:Q���3�Q٨	�1&"x�F1���~����D���q?��k���ec`]Hdkk
�</Y?��v���j7S�Y��f?�*�2�	M�)�'�����a�/�0������Ta>,�}�lSf|���N��)\�q�x�W�!��7HxJ��@0}�C�A}M;��z|�>��pG����I�IW�ؼ��mQ)���ˏ��B���x�	��k�ڽ��e����uO�0�O��V�1qV�|���>�;�x�&-��(�J~3��xP��c%[L6}]����f���\��o"�a�̼��]E��@��P�R�a&Ra��~��Y_�t	�a-Qs�h�iTn�g��p�I�8�Bq�L�R�k�d�\{@uq��5\/)}�ƾC_
rM����I�J$��,.�N�����'@�}۸�(BtyH�Z�R
v�~��qo�40*� 8�<�zƃͰ�z���m�CI�>���Ġ��3D+K+h���P�~=c�����b/i�����q<�.���Z���Go#r!O�i_//�*���뫛"�9���y�B�-�&Uh�ﰒ�Q���K7!�>�d�=r�k��FH�a��}�(|�9/�)��r�U\��
nB���TfO�@YCn�AD^�=�&в�%��i��1�K#l��M:���x�y���Wr�E�p/WR?	S K����{�w
p`��(L@���M+f��a�(X��F�$3�3%��O�k�	���=I�}��,-V���w����444ǣU�b�bK�,��Ӳ�9�e�aK'hQp�`��)�:R���3ͅ����U�i�L>	��<_�����PP���_�8I���ϯ\�\�qz>�P�F�9�R2�����<�=M
�Btr*̄�ʀ�2s�|�}H�c�6��<�4�1�ߥᢰFz2`��)��1r  ���s��͈���n�� �ǐ���>�Eۣ��������$�f�'�H�3۰�2kX�3��Ş�"*�sroׇ/���f^�T���xNlsf�� �HXeLI�&yo$-���G�ؕȎ��RD�u��\0����%�����@z�˫���Y��M���ƨ  8h�yx�T��xR��x2��^~�y5D�ئ� x�����������%��{��x	$*�s5��&E	*�=��:�
�i�!얋��}�p�߫B��A�DA������649R��iK��:�w����<#���]0ȃ����Q*���88ؠ?�M�;g��:�J�	YF��ȫu{iȰ�\`sFA�:c�fC�*�?i�ٜ�a+YZ����d����ա>::�I�$��ܐx�L�S�g��1�ng޸��#����΅O.Ё�*P,]�����<�,)u�oa&b��3
GA�b�:�a*g��#}%�4�Y��,�T����6�" ^��L�"�A�~���]�k���d^9-��}���g�Ɗ~���I�'(��x�Y"^9��%LL���)��4�l���f���YG����+�{w�[�Q�!���>s���
�}��-z/a�cO��-���u|�ɢO]D`���[�PJ`��V�v�\f��ãp��b����.f�l̲
\Yp�FM��a�\8Գ��<�G5���#�( � �w�"La���c%�~�}�:�Q�NF��Fۅ�� ��,��k#a�R�������kLO���E����|{,m�����FJ&��U�obNL�%؉�6�'0f5��.\!�I�_3�
@$�����T��u���?3�
�	;�����_K������� d��m�x���?�B��r�k�4�6$a��9$#2Gk��`1�Mz��l|�6f�՗��-Ϛ<?�|�[�.�U�eM���_M�� ��qkv*{W�7�(�6�}����nD�t&�;�+8�i�ֻ�۳�	�<l�k˱�U+�u�u��8d��O���=���&�(,뎭��/�ţ�&o��������|3p�ܶ}�U�Z�#�zQz��R
����_�����8J���uQ��	��?��1�c��i�.�
I���z�E���X
L��:��^�y#^���Wֺ�h�AN��n��D�NQ��S 2��֟r�ZB�"#؎��C_��
�l5��Z�o�ν����qLsL�GQ�2�x}E��:�sϓ~�L�"�;��x-�x���Pm2)�>fl�n�pѾ.��!�3�
�5�����(6&;f��TB{e�\��Xw�hX���2�u�I�������1^�c�@�[)�;h������&��/\�	��e�S����bi������ꄶ�
'����:P�?�ٺ�	� ��F|����<��*�%ه�%7����%�v����o�?E�&Q�7f��C���/7	@��Y��G�g���:[z�a?T�ɗ *5�Qx�Q�%u�p�.�l3����@�+8�Vb�k�Z�}'y�
`�=Y>�'��]o am���w�D߁ݡku�$��BN�X3\�6�Z��8kK��#t��=�zߌ�B�-~O��>�eZ0;u+����w��2�+?�uor�����*���9k!�ߏA�^���8�8��������u1o��N��xST��K7�.)��;t)�8�N�j��}�o�3y' �|�Std����;Џ���L����pJ���z��b�2�6��|�&��|(��D��o�wZxk�`�L	�#g;Y��V ~��_�Y*���uS��l���r��>��*9dy�;���]W�FA�a��B^�d5�,�Ҍ��J�T^.���lZB�̡�k���:F~)��7��ٌ�[nsŽ	ݸ���(R������4�G�Ή7������B�eS�s[j��k����/ǆJ��(^,ð���(06L$�+j����4�,-�~L5��Tt��]�:0���i�,v2�~��d�)gmVv�/{EXIl�4
D~W}��nL}���.Z\��� lhA�P�+&��B,[#}��$!<
fͮ�{�d��T�Ra���$�̣���V�Y�Z)A�>3��9���9re�K�FKc�:��1�"�'K+^`}<a�WX��\�k�����#�?�M�
f���?��9%��P+�'��0g�ӼM4��Ԅ����sdQR�����C��5��Ӹ�����J��r�q�Rb�0����Vp���"� ���ۍ�k�E�*�B"�i�������e�ѠŇ4���|�-=.sj��(���t�p� ��X�MHO�h��������y��� +�߉7PTp���jJD�(q1�����/�2�#c*��F���!	Vi�,6uZ�������c;,g6�}���{ɾ����7]��Y9>��Ŵ�>�c@)0��>�ｨ�
���"tV��Vԍ��R�#/���:|K�RSd��b��N���,�������B����̰:R\Y�kwnȚGS����D^�	�R��Ѻ��S�\��9�T3sqD���o/`n������ڡZ�[2������
�D,k+`���B.�Ty��p���y�$h��xݹR`DjL�|���a2|⼥��|Xm�E��m�RY�����F�Ѷ������"�*R��zN�>���MM�������qp���U+B��H �[[ٺM��*�+cߵ�vÿ�e�)�����]m����;AvR�*�Po��VE��_��v���O������� �y�,�W�g�c&���.K`K��f�jY4wR�]�3:��6��|���S�����)��9�TS��iq�ǌh;��_��J)L�	��"0�3e��ag�M��v[r"�ibHM�	���~?z��<X��7�A����@Vk��_T"t*y���Y�盀%Ї�^�����:�U�I����V��I0��jͫ_�۾��_l%}�cn�OS�1p��U�~ad�Se_�z����i�C���E��\Ta���@Z��[�uI���	�v��&��z��8޻"g=>��Z��om��؜3��٠0��y�R���A�/�T�U�V&�s��o��/���-�M�����jH��{���"�Z�l��Q���Z$<j����XY� ��PN8�e������v�+}Cn����C���4�tҎ��5�1�$p9�E雯�ai�����@�1͖�%�-Ć����S3�܍>��M)�AH�8�LӖ��WIii��>�IM���/�-bمK[j}�c�Á��8@�x٦i�6c�9����+��K����z�('{<3�А^H��F(�9��JF�7E<ٻI��<�<x�U�:�s�\\ޏ	�^�c�.l=@I��
f��ĕ:*�K��Bk"���Z��7Ф�TB�����H{�N�V]*m�[nj��c@E�=�q�����ε�l;=Ε�Ŗ3�6HM)��-��gn�QȀ��'�\ӄ�ҀC���6@])���/�\@� 8@P�՞*Pp`tR5��3��C���w��%���ődWC%A�lrec��"Z-�3�v�V�&��k��HɤBNTH��� ]%�%�Fչ���?d�Z�8����I����l�)4'�B/v�.7A��MC�t��E�G�gLkX�B�l���zE��)A�����"�FV���Q��Ԩ�7� �P�����Or��λK3u�Fo�+�/f���wa���d��9lb]�6Q�1b�OJ����)�Yr��4��zW��U���
}j��;Qn]��b����{m�p�xqRp�����
�|�ȼ$��D��Q*M�">�@��*�z�e��b��+;�\�B���s��J��A# ;�"���^��7�1Za�m"�4N0oARI�{^� �3�y��,�)�i8��+/��!_V���K�E��Ri��Ka��n�� ۳RSʳ6)K�n7f�j�`�\�yT��28��a�w&�fU��nt��$�@t�����@���~�D�@�u�4�>
A�JDa��O�}8�,�ls���A&����2m����/�[1z��w�$���>+�8A_�Z�V���F��=�̖u����p!��� ��uq�@����v]�9T	q҃���#�6ieLu���*���d/�j��.�᠀�ǔ���cW4�%�������ݤ� w��@ Na�s]�]������?P�MҦ��NoϾ�ȝ!QH���2�?k�g�멣u�Q��N�`��E����9�̵. ��2�aw�FJa�c�,?XN/Vr�LMm�2{�/��NQ	�%���Vs����?�4_�$����}Cޮ+͒�����w�Q��|:�n�s{�\o����J�;b�dE�#ʸl )Xu6p�f�o豇?E�T#L�]�ᥪ�;ruB*V.�v��=^_a��$�Fݽ�o�Ә�/�����\�RuC��;���#K�s&V��+rk���So��DBca�[��\Y]�!��#B��k��j<M�&���ڇcWmd����^���dMہ�Og���yW��]�=�ׁ��1��'>[�r��ݖ�xh�? �mƽX[�Fb4��r� %wC��9dF�蛀4L��Ӝm[ʀ-(X@@� @� �ᴘr՛@�T@��e����-��-�r�]��P�v h�뮉�,Q<�2�=;����-���e�pFkUk�B&cw����5�h�V(�[j}A�W?g�I��A^[�˸�{��+ܗ1v ����ĩ�����\lz<a���akw3�ӫ�S�>�&i���e��� �y��ϰ�o������̭!i���GhU�h7\��#D)�u�F�Pr��ɣ��V:�M�̇o�4Ɉ��F��_�̖�ٰ�����J�x���sH�_��-��B��K��:@eW$�q��"g0���hAO�ڜI=Ċ�w��Z���gw`�rʬe���u���������ZZy:%m�Ђؒ-W�&qs�))VXtc�k76�^���o��|��8#��O�p!���D?����4S�l�1�0l݅\� e�H�>%O]4DWQU?3�ZR�^x��7����/�iF�.��X����s|�R���u�*�e��I뤶��M�٩7�8�=��BV��wU��-�9�S[����9PҎ���LjZ2P��@򂩼/oDq�;k'�I��%�d�N��f��t��l�L��F�D֝���AU������X�W�+�(��K�������h.{K�&�7�M�^3�'s`�N��&�I�\#잔���Ki�mT�j@�S-W�&��n��A��Ϲ��,�z3�'e�����Yw��6���"(p\Ԧ������7۔�G�T^�eMf�������,n0VwAi/�GO	"}8S�g_q��d��ya��P��՚�� MD���ǅG�G%��3�F�{`V�ec���ߔ��@q��G ���rX�Y��O'2����&�]m�h�<s�mJL���;/@J/�>%� ���FGԒ����C��'H��N&�1��;P���`F�Vv�S�%�4{�+ ��怵��Nm�P�r�S�;C���w;��<�;��r>fA�����Ϫ�P)��ʓ@�f!�mb����I�q/�W�OҢ!5�C@����-�� ;R�4���ꖭ��u�⑎��n�cu�9i�h���H�R�{,ZdA����FH�Q�2���zG�|K}�)梽;��+M�w)#n�^�id��FdV��R�o�rRaγ8�RPف����2u2n��Np齧e�T�tFo< gq-�j� �
�f��CB�sw��Z����	i�x|nHCj/0=%~�K��`���\O%ƀe]�����_	Zr\.��0���D��&�Wʸ��(H���Y�jRC�E�����Rp���T�a&�&0XPL�������`�/u&y'$ةPι�(c}���
fh�$��}�rWc�Sc�Eb��>֓et܆"i�1S����.�6Y��5�^3/Gn�p@�ՙ�\��x���4���]���gn��N����th�����ԩ�	��S&x�z~��|�Y���ѱS���z�➞������0����t�"�������q�h�lY���2ZH@��z��0D����I+���RZ����h~��3P9�����k�18����"ک���}9g����d���07ì�m9@{�k��ey�}��dyW��?@<ν���ρ`�5�Eؔ�5��Z�w6Lb#�|���6J�i����q�M���	KBx6�Q�QFO�S�;��e7�[`栞�Y1��)�x�y�7[c�?��Im����uE.m�C;Je1��OF2���AL��1�J׋s�%���"���3*�l�[Ȋ��JvX�e��: 3���8؂��S������&�>��3C�	�tO<3�[H��:���gz�yj�dؼA���I#8d�,^���VE�=�Mx�J�]�F����b=J>V�}�%iͶ�fɮ\/�;)c��������P��{u��c�2ڰڇټ��l�p��&�X���͐x�!���-���j�C8�����}�������\d���D �Hs�_kiY�q��F�F�J������92�/h^p�����y�<�vE�)u�\�p�W�	=��Bhr�l�nlth��a�_�5d�݈��<��ؒ���t��
$���X���tI��K���?z�9�
������j`�����8��Z��b@�_P?��E�	'4K�}1��P�K7�,߬���_?|��l�����r���"���q�qV��!?��7�����ư�b����L�%B��cbR^�9��voZ互��Q]O��	��-}t�4U_�C��Q����x�y���Ұb�U���<���:mtyQqi��oG�v�^����c�N*0_�o8�H�L��.�hQ���K��f���/ʗ��}����?></�0��̺�c�9��� h�'E��ռ�Qù��'���p�cQ�.��d��n���e��O�{R�5N�@2�_V���Y_��]1���)�_@�/s��EUuj�����l��c˗؇#,Y�-�Ǎ=�����
��3��MB��Z���S�9�g=���pd�W�߾ncT~q�U���"���2 p=�Z{��N�䁼!=��'��DK|;u��q��K���d#䀫46��&[#N��lz�QW�� ���Wz$�+MnC"�=�� �9П����JT%�X�
.��-� �c���N?��ܲ���&@�a�G�y�]է����񪑤pc?	&��8Ê4	nI�����4I�Cй�D���'s����-D���x�'��,�|xg��-�f�鱆aWf�Oh�q���>�2:a��80�h��Gn�����R��4�n(�"����3�kՒ���D.�,	���	ˈ����,U�2y��<f'�X��t��`��Ӧ.�.L#2�����̓��Jz��[�4�";�$b���LP�xf!
#A��^'102�j����}�;��2�_�,u�$�e��p�m��̛?�mu'���m�E�'#��cc�:ndUo�R��:�~QcP�P���)��S|<|	���|Ji]	V�%����՟EN"(�<�	jթ����+�p���F�/�U-Cߋ�3��&�4L�G��Y���yBuu(qD� ZN��g��[�!�i�[kKM�����>��ltt�c�d�n43J�'�1K���B�!�ﬥȄa}^��6�o8����^���'E��s�_m��	�E<�bs��(ó�k��+P��(�?*�%Mq|�.a=�E��^�����f{�3�f��:�@�9]�5�5�V��6�E���M�e;	v��v�X��$}�$�^x3-�91�:���?w��U��[�yD�"��x?8e�F��4����_aS�o�V�TP� x�;p_<�	m�a8��L��P��Jζ��
 =C��z���C�	~�FK�d�,��u#!����	�Y������+�ࠣ�:t��b���=�|�	Y��,E��	q�o�2%@O�Xh���D���Ǒ~=�l�L`$fαDw��G߽����x&x"3T#?2(��&���r�H�)�e���4��?�� �j}�'
�w�vN`��ewmk��:������x��^���ɲ@(T���T�k/��S�5����B9�"��
H��ԩY�Շ�	�ߒ�<�tm�������G���S_���n�QsH������au<D[銣@�c3=���H㻓&���oX?:�h���X��|�!��`z�+�<��3��^� �=�2yC3B�u�p(D&�<Z����⣺?3����
p&�=~B�P����� s��d 0R��Pb�D����bO򻮈�m����(2��S�!��H�fu8��%	��R�������<��?������b�}�zɿ�L��-L�%m����~K(�h�¸�
s��M��Li��R-@�)Pp����)*B��s]��F�+�8�8�E�@�69Q˛n?pBv�7jJ-"�ϗ�����j������v0v+��%[����?�п��_���y�Ђ�׌Y/�
��:I�n�?`\v��2�xM��
ڝ/$��
��!+nA'0o�ϦS0T�<6A�Z�#�Y.E ��d ��1Ӽ����;u������������������1r魳��Ie�oD��U���B�$7={��������S��hn�O�Y#hkS���
�V�A����s�x���ٹ�~�gȾ��$����}
�!�suB�l��sgN�l1xDk`�vG|p6����\��A�X�ɱ���lr�d��B������j�ؖ�p�D��0<�r���:>���'CU-S���߷ǒ�"��o����m'M�!�95��Ml�
�^4�$(�?����=,|p���T�ڐ}!�Y+LB��p )Ʌ�1��u�ط,�p]/7�м�uf� $+7l�F��'H��')B|������l���O�ΰ2�[�gשZ���n�X�Pr��rVI���3^M�^�}[Gů�Z|7�%���q���JbzcUn4�����2 D�M�tf��.��x�9��H0�0�������3���c��� W�9CG �x��&Wgy�̀���X�H�̂������ES87�Ι�ʛ��[�����|e;���<;7�f��ꋰ��}�q���@�;����&
�0\�j��򺂁rL�IP&���	�h�����V�qq�`�<��N�T��,P5/����V�����{R�/~�M���@t��Kp�+X 慏�D�.��8Z'����k��k��&��ȞA��up�&vy�"F��G�;�+�m6OoMf.��:r0~·�'�Dq��[\��L� }��з��}a�9�|��8"�X>?��Z�����̔�堐��A;���i�
��30��u�N	����<������T7�I��1������H�<�q��"��+�Q��W\g�)������0�����1Eo���U#��d���ұ�br��p�u��-�V����w�c�^-A�����%Mϕ��j�ré�����a��GQ�����ࣕ�h�g�����l�O��]dZTǐk\�L�\�AfA$'+�s��CT�y���'������9�ʿ��u-A|��"ws�32�uӂx�au�q���p7Z�/�+��<$����m�cfx0���4�4��7Wt���?O`ܩi@*O:K����ՉF����(XTgHěc�����Z�2­������(NdI�T8��c���q�Q��h�7#Uԕ8Zd���uEO�l��*9���1?��fr�f5n}zd�������}��,5���: ���8tF�q�����{>wٚ4"���&�N��� UZr�*���SU����@��˘�����{��r�)���h\�q�����ݪ-^��n-��/_���z-Im4���jq�[!��#�v�C�39��_i��6�`�M�9�&��^�6�~�8m�G� LQ�`�Xm�yѨn�tl�{��H^{��(��O�����:f��Q��n��Y� ��X�![��ʌwT3����l��L�L� ҙvV�v'�]��]<��v�F��<�5L�O�]���B#=B@a�@6Y��%p#�[��S�N��8��}�m����b� ���R�$+�V`F<�����M�6�B�6��#����d��J5�,�H�,�+�S�xW�YfF+-����U��:[������"i:���>�4�i7{�%sC��qa���qn{��X� ��a����~��r1�y���I�6�!=�N�'���b���z�AU������M�\��f8r�+oP� %F�� .�G���@-h?Vڂ��檎�Ċ��	u6�0^E�_�JX~�`�[���mhvμ�7� �Z����gkG/���f۲��>�&��*�X��J��C3�*E�?��&���<��£�`���d=��X&]��bt(F�P���>�XK�m�C�$��bfZ�E5�wΘ�G9�c�N^^r;َ�XK�؏z{&MZJ�I��J��VHN0$��6�`rf���w��9x�_�վF�ZMV�-RT�2�~"F��]{�X2{�#�u3}�iE`4խmϜj�(;g�E�h�Yh;����2r!y�!$��n�	����������:o��%>c���g�WF��Ĩ(�}����v��޲N<kD�t������A�\eV5��KlO��DV]/�Ve����a�̢���Q����bf`��VVr��4���KNU-�����
2άRY4ޟ�6��cCV�i��p���D�v��5)
�S��6X�<'~N� �ߺı���/+�0��Q�Ę~mw-�gh�T�>'l��D���x���K��D���gw`J:77I;�D�ӻ�1.p�uס�����Hv�����T��p�dc�}��'�_c4�ΰ��Zc��"�@7.��'f���5�*k���ǫ[.]�/�����q47���E_�
����������!4�T^UH2�ȅ��ݣ+d�WM��N���hwe��H�^���ע��Iw�C���
�0�M9_3�}g�d�I/�7�� i�b�l2�S�E;'��Jo�zٳ���a�C�hyV_%�N�X�6NX/\h�6e�n���h���W�&Ӷ�ci���${�jm�8+��5��J����MM|�x�((B�T�%b����&e �����c4B�Z�VR�TwK�:'o^z�K�5W E���}�Z�k�Hv��c/�g񋇲�L��V�g����z3�g��i�kCP�Q�abo�����
���Bc�8�B~�{+��p��5棪�P\s���E���g��� ���oOK����l���'�S��1MdH'7�_����]^�����3������fb^����L���'ϧ�4�Nu$t+]�4P��dQ��Y���Ȍn�3�"uu�@#V�Μ�J|c�?E�_�V�V���$�jz��`(�7��C��{{��)n�'�R$5�a�*��ի���u#����S���b?Ȏ�״,k��3I���4#�zֻb�vw�4��>��[hs�JX���/�� ڙN�����w%�T9w���u��v\m3��r�� �4��=K��E�����Q�Sl�4j&@���k��4�s��ɤ�{�ͯ�1��\Q���O<GJW^H*����u��Ʉ�Bu2��5���� �윿>-bi��!G��-s���Z�3S�Z�����p��S#�����4:x�P�!��c��"7�uGjR�o�a��j3/�=`of��x.W���� �T���~�U��N�Iİ�ɉ6����t��D�ёͭ�'���@�%Z���H_n(��)�z3&H#�1F݌�m%ު��١ s��R�������u�(�0;Rj%�Pp�� ���T�B����"��~��`�Ƞ�X�����0�A0��`)���C��/l5�=�E�_a�0��&^�	�p�>g/3eۻ$�R����<ӖW0�R��|�d��
���37�����wc�Ë�n2-�PHi�/�1}��5����^���ż��B��۔���(P
sʡ�B�ڥ�m���YX�^���/��-�ֲ��ɍ���f�LI+b��p���HS����8#��AD�ΈO�8��۠<Q	}�p��������}9њ������1Y�Q��w�o4��b��9��
�f�lv�傊��V=B�t��n�y����jq�5���x�ʜ˿���x�h���5`�)-[A=/�:_�ٔ��`�w'��?���?_��0zk�����c ����^1a'�i%PU�P̉UG���@��:����{	�L����/[B�iv)}X�]`������C�����a�o�<6Y��3I��<��T6xD�W�j˓����{�Wý�&��9;�"�4��o������<V��/��{2�[��.������1PI�+�@w�3ۮ�l80�;�X���>�8�����Z!⼨�����j���0��5ʮ�ze�v�7�e�@�U~j��Q�a��2��O�)�]�I��a�f�S��	�}�AR�R��J�p!8s����].'�?w#�����t3%<��S�Q��j���%��g�^��v�	(k[����W���C���!��^�H^lü��J�ɻ�+\���d2����f�v���v�_������Ԡ���4��7-�b���c���	����+7�C�3��Xi_���W��y��B�y����5W���3 �ޥy�N/��5��;7�u�>�I�V:՚����0���8.�گ�ͦb����m�L�������"��2~@��(a�_�Lqz��B�sW7ŭ���j�l<I��yM/�ىʜm�X�J��)���Z~��c���.�@��2�ȁ;�r��/�SʤON4��&�$��1�lW	��r�5k;Z�kA��4�V���������rD�Zb��m�B��P*JW�/}�µ�g����N�"+��;Q[��'�P��fv���-�m���!�|�`��恮ֻ���>w�!�ptu��^"��I,�x@A�}��V�I��4	wE$��k0-T����f�|��n�{j��\y '���=�ȂnA������*��[n/2b���φʬ\������|lZh�O�� �F#` ��g�HӀ�(����
~� W-�+�e��.�*�� a�x���f��f�"ku�̩�T92B���䫓FT�Py�8��%x�VB���g��܃{[h&�/q�\lx�c�y��U��6��|HV�P�깑�Q'��p�8]\�4�
�L�פ�8����k k
�(�x��I�X*1�o�]X/��͚����{�Յ�h�8����`QD��J�%�7���'�jG�{Ƙ��ܱ�7�<�'�2NS��W�{猍_Z����`Iٲ����G�8g���A�7�϶ݵB4������	\�a|z}-�9��?��C�w�Ь�:�^ڥ�ys;?��f�+\�����jr��ӮF*`�.�����|,F-���k����{������!h�H���R"�b�pȎ,�p��FÓ�q����?A�%Җ~e����^����n�*��N����hj:w��p��I�B��T}4 ����jv� �3z�����)[;͓�Ġ��zL�zr0C�n����@��~�?k#(Q�1�)p��ŵs�A����:'ж���#�BA6Pm��X P�q��ɪE��A@x����$p��l���}v_wvVk�S����g�����e�%E�}Ρ)�9��V��T�E��rq�b�kЂN�[{�s�=p�Q���{�@i��$�RQ.B�o�*_"�;e�� W7yw;��*���o1Ov)B
|/�J��z�9�I��u��õ�H��{(��O��	W<�-v'�}8����Rºv � ���ۗ��l����@ ,#J�(�Ak�c�,=4�/��H���Px�K�B%om�����h�Z�3yn r�M����q������L6|���5ai�Ά.ce>˫���ۉ�ѢY$18�Jkn�~3_%uH��d/��p��H�Q�|#m��#S+?��L#Y�r+
@����1��p��%%�.__��k'�|��,����]�`Kv~T����.�c%�􈣍؟��.��M��If ƭ�&ND.��j���^�Q3�����:�������q�)h^~�y�`:Z���өd��.9���/�MPv��m�YT����=�*kalE�gr8%Q��>gL�Zj -��i�{pUH~�<�Sr���0v�I�؇�N:�(@Lچh�A�y��'�[Gj=���C�Cb�H3�QW\�fS�;�򨢞o(��v��� ���-�&]�xaY1�tX�Ns\������^M���w�P�Xs�q��M�K�ܴY<,��/�Gn4*�{��E��??i~��G[a�E����Q��lمz��'+�)j{J�ԩ�F��}-%���p9e��OF��r�O�$M���WV4��VA��G��B�z}�8IW1��5"��Wc�{E�92�(C?��5���
���4�a�h\�����i$v9��|�0�q�E~!����h��L�t�WN@)���Dރ�!��k�K�Z`@�\д�Oyz#��&�=�PMu\����Y�3e[P8Q�=X͂�(E�=t@8`�������q-�ط�P��c{�>�߭eh�J]� y�"��n�m��U�*�Q�q/���?3Q��ͯ�����h����n��2�Q�M��VۘQ^�R����ENc�f�Y�|,��E���	\=Y~��g&Xz��âs�J�T��ת~�&�z �"U2e�p�!�wKcE��]��}�4���VS��\S�\a�UE#�d��"�$\?��f`�q���0��(m��lqM�	p�$Q"��P����K��>�q`���t�r����'�~��z=��m�W$��|�Z������"��`�d�Ѓ�+q�3���y���=b/e�g�E�.g�	r�ӫ�;h�'�џ���)v���sy#�Q��L�^�e��ΩA��pq5���G�ڶs���(���:�o ހA�� ���m�#�Xz�To$Ҷhص�~ERm�օ�篬-��lBU��g�	_>�8ǈ��vJ`9V�#�D=@O�0�EHvY3JԿ�������YUw�)oy9�ԁw�/�⚮�C��W��x>��S(��������S<耐#�]���ʏn�4��x�`������v��Zt=t�1]�S���x�y�=��m�m+6��b�v���;9 ��xX�ه�����i���>�]�mZ���6|HcW�\�?�u�b'��Ћ_(b�R������Sn�=�� ���{�R8yMXZ�����+YR ����9�=nW��T:��B�NbK�E�d�4i�����J��� ׉ՓR(fv�A9O�f2�y���������-�􀥤�Ϧ1��~ps9�$��OƈXo���	|E�k|�{mg�F��faMO,`���}2y�2&5/�%cSt)���'��i�V>�Ĉ��Gܒ�o�V��ha)hNm��:d�B!����sP9�r�x��<K&F�+�����Y��/��EVA&��c�>B8�m�JSEPU�ٲV�o��ÇL��<f)IDt3�ῤ��a����F�V|��\�0S N��	c�n�XЍ�8��+o{�����+���.�1��^�
�Ou�V�ť��5��^�k�3�%oǼKio�|a��zv��ņ�)��d�������-F˷B
r�=�g$���8���4C5���������V��W��f$&�W�\��% ��Q�+���1�i��/�9XƼ�D���SB%<�
8�E�J�9�Yv�a�����,E!����1z���\�w�DN��7j�=�
��d��O7 3�5xr�|�����% |��GC�P��c$�~A?�*yOUD]4bO�>�,7���c��>V�:�6�4�� �3cH	���(�4
������7#�fWb�f��Ǩ���T�Cw��Ǣ��+l-<��f�3��������f��BL*Qo?��?s�����c���#iz�R�	�q@l��F.7@�����y���P= {/�;R:+����3���I����dbe��/.^������m����ƁtH��Y8����
�Z�c���2�!g(Y�R0O�����a%��q�wg�t��ٝ8=e�:�4P��kt.wቻ{������n킌���1���P+�9%I��0Z�`jf����C$�x�>/�gW�!�]���A�|�Fw�A<�搾�y���6�,ˬ�a@��]�����Ud���=B�9:T&�Q���OOby�y�F����6踄�'�;o�����ڑ��G�T�(���@;��~P?J�7�R�nz�� [��:�]�S�-J�ג
Y�2�~�2�}W��vG��S����)r&=HM�pXf��R+^�\��qy�1"��e�]�	n���|Ǚ?	�m@m���˃�|#�_}9���C/�`5�P�ՙ�#l}R=�^F%��h�?�f�=���r���)����GKei���7���@�Q���M<���W���SB�%�_
��ΰ�qa�G5QhN���zZ%#�}�?��C|cԟfDb�PL�$P)�eg��9Eimn�|s�U���~����� ��c��)((b_�mA�u�Tf߫�s�H�{'L<<����H0G��밲6�z?��P�~��S��F��c;Eh�
�,���5�S�1P���O���{�CClؗ)��o)h�ڣUD)�	�ۜ|w���e�@�(,�p��ͦ�������m��
��}��3���G%�M�k-&��5�М���(s�c-.���J�$�Q�_�W���@�'���#	Cx�-[�Bק!��A0k3Y�/����ɭ2�Zu(js�E��f�I;B9�\�S3�t0�'�R�B`�U�s�穣�g���D��k�;$�hj�y��8���:������&M��T�(��M�������i��8���i�@��y�L�JoQ۞��>��1,v�3�[�W��"����$d�j��H�%+�{�.C�7�9˄)��<CK�A�����yHҰ/a�KmP�8Əq��o�,-fhlãF� ���(+�X̰���X�ܰ��M�[�`�TF{�+����(�t�s_u�|a �Si��n����4Q���cQ�Ā�:+�	Óe��1,�"x��km�I�+0Vp������$�,�3��48�/�(��z��ȋ��:��lT�� ��>l\b�"U������ex�3_8��^��Y�
�>oOk��.���t���5���=S�2$y����P6�qWTL��\����G�g��ɓ�"�G��w T��Jx��NH# �h�{�t�1�������I�*K���r*��X��yO�X ��(�89]-�yx>W7���X8H���3$1�Vt�sId�ٚ��9��<��so�r�O��`×{�{�l�y�~��~;�J~�t�M�Č�GJ�Wy�Wp��LLU�	�	�+������+�$��J��T'�U�O�P�ڮ0E�"�<1g�|wY�_����̭�.��"<[�}��Y.A��=��W�"k�Iuo���+���l+���{�a^��+y�b1�v�h�%]�v������~jN [^�����㖰�8S���� ����z�s���L������'q+w��B�&'�F6�H�?� '+��h����WIh�/�:�����_9!8[��3�gض#���x��bk���M\������u�=Tt��B0�u�"����R,?MZ%��l����V����Y#�R���Y���[g0/����]�O$��#Rk���,x�/�6\���--�7m^}��."_-�DCt׍��"e�V��öڶ{p���( ��_�U�����t���h�'��=D�ү��ٸҖ�����Y��㹳&����a<Ԟ�����
�O���D���k�&�Ȯ<r-���3Y�|K��b�~5%ۖ){�������S5�XF[���f�<��[�D�ɠi걊�������$nU�r{{|>��c���='��l�`M!5;tX�&`�8�\��p3#��|�5���I�ʀ ,�1.���0o��Q˝M"&��]��'\<�7�/�awS�%���-��*��u�Ae�{��z��8����r��󠻬ӬF!lc����(�i����ȥ�\k;�3�+�kʉ�ڎ���	}h5���Kak;�MGY~��������g�D����:��b�p����Ҟ �[E=��.�r�?��	�`�EI=O����e�e�;�c����a`�(��=�(�og�a�8x��Pn��~��=���1��!aw9��3��6������}*G��U�@T7}��d��p��dj��o��r��处�l�B8��"�v
&�"�p��� ~��~��h�U�+S�J3�}�K_�س�T���F��@l\��O�@&5Q3�&��0�Ppf58��s��C�I������r?�LS@�1�n|]-?k�9ힿ�y���-W\��^�O�ms�Tw����_�L]Z3{�9-[E50u
����Iߊ]�Һ��J��P(8$��>%'6��$7�Fd���������Ԇq��<�b# w�AG:��7v���qg����<�.�/Q��?)�H��2����!m�f�:��]p^��s���C�鷁�us��c���zۘ
5��R� n��i85����h ��q������a��o{�d;�Cv�!��˲�}k����~�	`1�Mj�A��S�����#� �ע���p���m�L�zSv�=/���$��%�vs��-4@�#"�Y������B~��.�����N\x�ƀѲ��P����Z�u9`$ST��T5Jߩ�y���'��0��#/��,�X���L��%��������)�eZV��s+q��eޛ��l�Y����7�7����%Q����q�NNu�o����eE��n��)����tj��9|��"� /_@�2�3�)9�!�~V��W�V�|����K�v�(�vu��Y@�_� T�{ߺ���:���ԏiϙ�ǹ��� �u�����;�]�~s2�Vj���/	�N�"�ۿZ�eBr�KG��}-^�A�ڹ9��Dz�����L.a2P��x�;G�3�d⣌]���6����,]/��i�Bg��3�\�s�"��x�L�ǐ�p�?�O�&ܝk�0V��y<�3�X1�l����~� 0�X���T=R$X���6I7ێ��g��&@�z<5~����g��+�J/[�{���*mw�����K���`������}��Ǻ�g�7���=���po����2��$,��&pk:��wk��4W���i�$�������I�:E���Z� q�`�*_�a�@�l�oբ�.q�&��6�=�Q^v}ũ���&��s��U�|fm���i�l���I{�����,J��!�=yOg��E[2��R�k&p�һ��r�k�3 ک���
ָ,X��w8�S �z-YSAR^��&�W�O%�ԣ��[�����뇬�L�BrK=��bսn�l���蕕��#*t�����k������#H�¥W<7Q��1u+
?�����T�ae1�U	�2.�Ӱ,nu͚�A=o��0�4Pa:���0SN�(7",�a,K�k�um�<U����� 1�d�¸%���f��r����o<n��˺��lEi�Y�d�G��q�EJ����#�Y��Vρ�]6�)3�Tg^����&��[K�4u�<לI�VT%��2�ըKe!08�N��%�j����
�ΰ+iS�ft`Ll�i�zᐮ�ΔڊM��m[Vw��d��:3�]gGXp�������N�BB��������K|G�j�>:�����h��E�k=V��k��B��c�/�l��5��'xj��̹[�#f ��*�{@}�x�Eo�K�7��SK���鶊�B�g���<�_�M�mBV���j��c~5��q���j5��V�w��,�{�|�L8�͚�g$"`�!�Y�O�E�Pǒ���T��Ӽ���|sA��ki�И �-U��o98ό�Xx[ԂbVZ���v>�Ti��6��a���,f�������V�^��uÖO����j���;�A$zC�^M�.�+I7!�G��	6#�Y5����	&2�tpO�{QX13�1�'����b�i���'GT��Y4������������>l�m52W��Q�.�,���.���_�a�yb�pF��;��Lk�;��g!4�F��Y�LJ���|0ZZ�"z�d�zx����
������?wI�a���?�y1'�1�3��	.}*ԛ����i�Q��@�t�H�#9�,N	�
7�juUPS�n�+/���'r(�˜���[���f�(��z��b�⣄��ށj���
��$m����y�귇��)8�~Lf�����q'�o�5��}�80�˘�+F2Cg �=���SW���W�N�Kcs�Rfrg.��ͱ�W�N1=WcF����/`����1^�5��!̱�L�G�����"��0�$��-�y�_/���`�h��^i�����k[I�O�
�����.�H�9P������XKl����V\�=toh��"U�9u�#{�b�}!!�̈́��=�~lv7Gڲ�9��"Cx��æ�l��/!ZY�gK�W�F��`9@�~e U��H���`÷�V��T�q�3y�%�V�m�qy5��j�d�Ҵ�{D���-�����FB�`����.�H��G2T��$�^f��ݵ0|�^$f|y 9�\&�BW7�_Mn�J�b�9�QeK�k� ���V����k.�  B%�%����fN:;�2>Hꔁ��T~W����c�lo�����B�ю�XULKT�aI=�R�x�eń��\uٌb�4,W�����4�0:���釜h���at?Ls�&8�+����稗��_$6���c��!����t֫򝥏c.$-g�)^MA�TB`�J
�OڻL�V��i�YfY�O'=��r/���I'#j�&�Y���v�R��td�֞J�И ����9z��~6f���E��/i(����>�9�f�֌��
]R8�;%2�e�}�T"�aČ(��	=�J�Q���i���7Tn���"��S������}��Gʕ���0���s2����r�!4��W��O8�˭���s3|������^C,�0q)>�L�Dk���f��iI�#���������_�*�>��Z�A�� ����O"�dXQ/4�WaUA
N�)�	f�G-p���ػL�[<!�L����/	2٭0�s�9<��Vm�b���s�C�zD�k�+ �!g)�(���խ ���M�\C�Ӝ�;'�zOCR��Y`�Q�v<���9��̉����h��aN���ѭ��%���Ga�Q�xgZ�6h^��*��eԱ��	�z�=�z�ת����ߟdS��|��xW��ݦ�la؎��	��o�h�c:�aY�&� v�7��M*���M��m̨Q��B\��<ô�u��t>���8rh�69lt�!�7�=���u�|4�n�;�4�DM��4b��H���@ ͮ�6\�����,�9O1��q�t��-�bdϪ�yw�4��$�J����Ǥ��ʈU��n��l|2>��
� (� ������
�Ò`~x�
��w�Ŀ�;��M65�
W RT�7?�-}Z�՚&�gFu������J_߮��TtA���R%����ӯ�g#�!�W�f��������D�6�y^�{`�$���D]˘���R���m(���S;#�b�6�R�ʲX��-E2̟�Ř�XZ�ל��*���r�(�O�{�5�u���yR�'Gd�� ��4���K�T�6��40�V��a��Ю@��^��S_����(V���%�3��D%��#�u"fj^L<�_�f��?����*t�r�)��`ǣ4���D�>8wq�3��]=o�q_`z�X��h�,FU������%呏T��O#�H�ia�N��,ģ��L��p	��O����4��[����ny(�aV�̑���L$�x-4Ԟ'�J~q46����$��*<�h��ظ�T'�����Ff��o%�Sʹ�1��y��yY�x���~��w��vf����:y-�q��Í�Z~�#�!���ǁ8n�m��=�%���rC�W>��¨���9qy�H���t��E]s$�Y}���]��ESr�
��"���SNZyl�ko���qx�f��Hm�}_'�W��6��=��+����(,�h���Z�m�������ÎC/B>U�R��k%�)�G�:z.��c��v'k����S�m�P*�?���JL��~c�gp�O'����_w-7�(�Z�B�b��=z|�at�mWq:��zܲ�����3�'�T;^2M� �Ť��ny�|(������n�H7Ϛ��C��
E0�uQ�R,ǫ�H|7r���'�>oUܷ�ʨ�i��'�$3f��)��ӷ{��L�;�=�{֓Ed&=��s�c0��j8-z:㰶O�(C��<o��gFy�T���|ڡ/`E��ɨ~آIJ���f�J�m=�M�&�i�)���@�B�����sS�I9�:�,�WD�?���D��BLZ�	^E�i�eڞi	2�s����������$.��
D���ޘ�i��0���1���C{DN�o
Zu�ܶ�F���@�6��>�:o��ԣ��J�H���}��Y�GJo����n��ө�&��MƧ�D���1�%�����n+�� �����jQ�Rٽ@C�)|K:a��m��sPK!K�,;5���=Q?���9���'"\�:N�=Ɔ�i��v�e��[9?�1��1���&�)�lF��^��@��A�����@��8���q�Z�� Jɸ�p7.�J�b�������Yx�[c���J�+[Z��`8z\��Cq�][i��� ��H���]dr=���(�3�-�2m�R]E����ƥϸCX;�W�&��x���������ӈ�LДh�b�f���� j����0x�C-�n�hc�*���. �l(�4�4����r�<�
��.UȞE�緁Y�B��@�7!8����{�>͎sv����w�m��hXS��z�k`k+c�F�-���+���󱭇(\6��uya���-*!kQA ��j�qJV��n0�S����B��C��L�@uJs�ݮ��N�=����}�]?�u�Zy���S��8*U�Ϡ�B�M���2u�jÙ�j>�hl�lP�d�M�:���*4��4��n)7�Uދ%���`N۵��˴զ�j�$W��I�Yϖ>O4�0^�oτ��r�A��o�
I�����i�� f�}Ag��jo�V���L5xt���M�Ӫ=���j�iS���R;���{fR�jt��O2/N!e\+�������Z&�k���l�;�r��}P�,������3ZzO���P���#��z����'gMTQ�R�Q����p�f���a��)��Q~#)[~?��LG���&AK�Q�L�8%3�ѭ�lР��:�KU�9<��6_��z%[i�s9�4
���L5S���{�\=R���O����e������n����s��ãA9�H��ϲ_������@w~�M?��%Hǀ�i��f�/�̩_����w�d�8����������60�,O�:���Ph,_X/�N8�����#���v��878��T]�A�m�ce�nn.�@Jv�'<��7��$��U�r�l-%$�ZRl�OU���u�'�G��ٍAǟ��*F3�/dB��q.�M�jβ�I�rA!�".	��?�v�RE,*Lp]�6��r*[���$d�	�X@�C���>S�}�5���^=kĢ���wm��U�4��%uV~�� A�j�gF�������pj���(G�þs�ƶ0�ʧ��5��Ĺ�Z������#���:ᙦ(�p;eq��uA=�y_�f^���--*�k%3$u
��"U��!j�iZ�_B>p�I�B?��g{�v�ۚ���V�ڜ;RW¼�E~�}�X���,?<eO81ɷK���=�\�4yJ�'��
*�W�! J����:?{�-y��A�BB��7��֡�x�5�L�`�6+d�Qs�9`�F��w�"��s�5�Γ�8~*��ҡ���(�)E�C��ʐp��p0|�?��"��6z����,;x�W1�/�*En�.i�A]��fH�o��I���q��_�8�r��=9��ƧX�_p��G���eE�vpf�kә�rs�?s���h/c8�w��y`⯁���֠�,h5��K�q�u�� �^��������w��e(A��3�]U���p�?_�,��tꄭͣZ�V���g��S��V7���ZC��߉�P�{R�YM~���1�������A�/(�]�sz�6��G�����=0�����ů���J�+�|����B]G�+& "���^�Q5�%e[�o�>E{�Klc8���	Xj=�>ѓ���ɔUuf�ǋL���>��*�[\�Pe��ٚѝ /�}_�C=��� T���X�sWrI�g�~�0i�
"юg���Y��L\��,;vD.���h��K�>�q�H.�v
LX�7��k���(�oE[�N0��8ʢͻ�c?�$�Wk�*���+$�껵��p��s4��P%g��3,pv'��"?�ް��zř�shC5h-iƙ�>l`�*��(�T�c-��J�j�$�hZ��cX���� 8O
:a�]�M�x%O�?����s~����0�k��F,I��RX����#�k���8&�{��9B���a#�ч���Y/_����S�*fr��6�=����Y'��ᛴޒ�1��m	\�����>��Wu���Qf�!L<跌��"o���xh�ƒ��� ҝQc�ˁ����o�?M����r�8��1������_�	����O���$8���=`Rv���:bp��:���W۰'rl 9���j\������-��(7&���Qe=U;5�LO�^��a��t�{�Z[���_+�֬n�O�5o!]g�.b�MF`v �}d�/�^GS�\>�>L�H��9c��_����V,q}|\z�����(|2�k�]j,6��T��p1~�p^�|�,�d�D�5jZEH�߲g��lg.���]l]H�ثl�-.ۤ(��9q]���h�OFa2Y���EY��T�#_��)���Z7��.�g!�BJ2�z�T���������0c2�ǱB3���9r֣ [B孑I�5�/�pVs��Ww�^i*�/�3Y2���Ŧ��?c�#���*��	��%�s��g�%���,3�Lie��SK��^H�*ĺc�TD���ڥ�{�1φY�x()�������^9]�*V����	�_�,t��-<�ml�*��4u�g�)�Qg�IY�Vڝ�Ui�_-Rn>��eV �-2H,��q8��LX��_p;�>�̓�ZNS/�UJ>.�|CT�q�'�7yS}s핶�A9	Pl�Yj�SB�V����Osl�}%�Xܶp
�
Y��I��/���M��^�dOΑ�4���Y
�{+�kd�N�f���^ e���#=�v���Ji7ߋ�q70�l�֍Hc��}_��rĽĔ�}��'�n�)6���Ld�#y>9��{׉�3�L��D��"�r})�8�[?��T�1m�w�����W�~�J�d��D���D�̟O�ɇ��8D(5´��v�;�F	��&��DY�5���Z*�S��/�sF���[�x7Ŷ�*ug�@d��<��3C��^�C�=���vK�NG\ ��#�
��/L���c��g� ���ʇ�_�/)wD�P'i2�ɉ]p $��чM��h	ӱL�<|3�+���B�ŷ�j��²��Q���U��6áY��ﯞ'؄_M�!Kܔ�u�M���7HŖ��C�Q^⿰x���
pIԶo 	q_3��r�����@��yNi�؎y4��믘 PE�y�]b\���/w��lG	��y	�㓕ԛЊ�5N[a�?c��E�Fd�?iA���O)�
���s�&eU�0'}��7|Fi������_m>e�5o^	�F�1�o�98mn��\38P�P�e��Rj���:+	�sK�"R�<S��4�p��Jا(�E��8֦{�7 ӿ+8��>��`vt�(�_H���M���w��W��X{��9��!2������m��Cp$�pA������K�x;�_�E�ˊ���0ClЇ+�Wv�	0>I�_�Ks ��۬�ڐ��&y`�f�bR���>�Z����C�X� ��g|;3�@Ut���>��el�*���&��T`�ܬb[>��.�����4��6a���[<j���a;�方�[$ �0`f�1��o����hCUuX��x���5$?\?����a�{1<Ņ�uƵ�ԣo��e�.��W����� ���T!\�����B���;�	YNw+�@\�z�'+�4��� ��M���ra�5	�v��~��l�������Q�B^"�j�X����G5���W���^5^? �vF<@�0\��֬��ױ����Q��(��KK�X����t_jǟ��Ǻ<2q��c�XR��M�������1F�6B����xބ�*9T�T��v1��CUmVCy'��&=!4�I�� 	��9<lb'/-��g/��w�SsWI�ɉMh�J�QD��F%&^%R�(撂8���� �@*v�Vё�`m����^_���RgA1��-����*K�%��� z�!0TK�{��]�}5��6�\t��V���D��\�����
L��D�|�?��pY=ҕ"E�%@lY��Y��Ի��l�ۊe����9� `O���bC�3��+��&��M"Gᐱt���Z�r��5T���gt�\�{���w�<��gj̈���=��ܟj�1��6�B�
�W2rЦ��Ok8)Q�L���8%uD��t�1�C�.s��e� Q�L��}�l���R�l,��n7�-A�zG{�x.�R�[��=���+PO�ޥk�RN�<I[aҚZd�j�>�~������������K"!���Ay�0��ۙ��H����`�?�M��@<��ɗ�k��a��ޏ�n�̀�y\�{��i��ljy�2%(aI��v�Es��Щ����S��8�Y�%���?-�?7}yj!��*0�@��FD&3����25�	�qX�i��B\�Y�8��Qo����.�sJ��ݶ�S���o��dD
sPx0�$J�	d�c&��1�WY�x�䦮8i���O�@�4�������X����`�ЎN`!zl��
��\��*R�օA�F/�#�_,-��!��\����AZ曕7Y��<s��RЎ�i(�v'`i��Hw�AP�B=m�%'����{�6v�T�+tCp���Q��ڀ	����Ϙ�5_���rƳ�;a`�P������?���僞r
�6�[l���I�18/߸nW�rR)t���!�P1F���.n��ŁcV8�y6��j|�x�(-� 
���![K�}�p�{-�"G�x�Y������J~��h	&���`^u�_�����ɭ25����Y�q�qdt~��̃�"�`B��S3�'~���@�'18X�*��1�W��i���m}��%�	�`ݖ&Y��w�B�.n���%���%�_����͝�������3�Oo���kžɺ Fnc����n�?�c�5C78�7��440:o��ԃ��1��K�`���ٛ�jK�|�3m:�-�J%���+,ն�)>}�'W2i��}��d�~���B&
z_�x�)i+�w<ᕹ�qO���PbN��w�g��8{�濐SP��_��Xe4��Ǖ>�[_H��i�9S�B"u�$t����>:�5,�TB�P��вm��SF(�CB3N>��s|�%QT�5��2�#bz>���%	�N*�}�,�����ɀ� �Pq�p�����D�U,	�Oa�R�Z�^D���ӏCX�8*��#�j�ᖲ�d�H�N Tr�uw��}���a�t����<��g5�4H�`[�P?"�y��t}2L�DAh�K�r�r~m��+ٕ�Ra�q����ൡ6��}iDN��?f�dR��[/���ʞW�����tH*�,�i��>!�6�~��1P>���M�P8I��H�@�Ȇ�?��T��/�/���<�3���>��ܰ�t������	=<���?A��/TU%lL�/����+�Vr��p$�Y��T�^Q�E�v��1-�G˸2�s�,̈́��=V���X`_�ϝ��m��Ķ* ��� �k(���h�UC�Ý�ZA��"�B"�
Q��!0Yy�&w.�DZzz�pQ��q�ƿ^�jc��L�m�O?f^���ðuΖ��%L���s�:UҺ�[���ŉ�V��}^��"g�q=��P��(Zv�@��f��Q;u�����c�=���$k�K ����@���M�����y@��^�7�$�+�95%��F�s���պ�	���
i�P��V� +��G�`w�ҕ��<���A���f<�'���t�^��� ��Z�s���-����
�gYi�u:�����"�6�*��jt/�t�����ԜY�����*��
��Rw}-��O�O����G&=Rɴ9��^�Ǩz-l��O�`2�/�'�r��Ч�9i���,d�rP����<n6�:5{p�V��2�o�?P��Qk��0N�BI7�>ٜ��=T��Ⲹ�u�r�'��.iэTL�0�YS���]�V09�GoL>�0�$�8eUD���L��'�'w�`��j���S�b=����t,c�?Á�[j)���42�� �Pc�$��Q7�P��~d��S
�$��2�T&`_�Yy���!UG�ea�k��t��&���緻22��I��Q�t㿷yE��"[ⓧ��5�&��}m4'�)`W A3����
c2�}B8�kx��;�;��N�F?�e��}�QP�$}o�e�lq	�u�݂p�|J��Z���a>mii�9e�,a)޳*��3��?�����mG���e
fO�6��@삇�!��>3�SI���$�i���7E�3���<�F�Vv�Ƨ�M=��5����$�P�c������y���ć��E)����'=X�݁@�aGͱ8C�:��മ�؂��!�j�^�K�}[���i���44�J8@h��]b��Z���%z�h�Pr�Ud��eB�{�E�0=����<�2j�X�n ��,��r:O�u�X���$kcq	t8�XV��)�9ӖOa�Bkvūc�Mư�S���`̛F7s�G���F-��Z^�>��#G>f�@�\_"��U�M5ǼSx�
r���{	�F���v=�X/����A�����m����Ҋ{n��c���d�$�l��a�S�"c���8e �B�#9����h� a(�����E����1	$~�0l��\��/�ڼ�ŠE:e�ԜF�_���P<�N^.2/[�4>���ˣ��gcrb�'�aT{d.׬i)-��2rrwP�R�˟�1�I!2,�'�z�o�>��x;H�2+nI�]@�U���c°Aݕx>�N3�ە��� ,���h|���d�Gn���	�r�[�T�������ɛ�'�@L.����K���9��s��}WQv|כj)P��	Q?����媓\��o���E$^��,�ĵ>�&$����3jAlP��l��z�"QA�ĻlB���/�l�?�G��	�f��>%#2��Ȁ�9L���\��V���gsKI����E�"�Pm�ϳ#" Ã�)�z�L�����>�g�-E������G�MI75H���L���s��&�Oge���Y�G؋���kY,�0Z]y����9�ʌ���Q+�gdӡ�7�͏/=ù� ;:���k�X���k�,���11� y����#���UM��XN��c�1&���`x�.��iBM����Ҝ���'@Y�ثN��zJ�Y����Ѧ��U�?����𕊅�INƙ��`����7Ɲ��_(�u��g���=	�J�[H��Ӿ��F���)����|�ILf��)q��;t�����S|#1�'d����6wy<;M���[J1g��� z՟P�sf�ޙ�w����9:Se ��"G;�������:�!�әC�9D;��	���mry]t6��Nk�H�H)�QMd�MRs7��ПC��詙)�b�v��AܪA���z�<�H�f� �-�W��u�1��d��Ĉ���t�Ԩ	#����eeBH�7����I+*����Y���-�i�*�#n�e�zL��-s	�DZ6���2�zZ%g��cm�ѵ�O{�9j�e�>�7C#��{���Y�� ����.���H��g_O�S>H�gkn▸�T��?�DZ#�Q_�&v�iN�v�'Z�����T��)R���U���"3/{�(�"quy��"o{l�a�$�{��e�7��������#1�! \]��R�~4�df��}��E:��Sh�C_C��Gz����&�(��VF࿷~3З�BUb*%�u�ў0�:e~��ݥ��:Ԩ�aܲK�?#�Ҋ��*?�}�H['��I��5�Fى����t�����W9�f�.�V	OJ,��m�G�Zt� K�h�aJ��=$D7%(O���X�8�u�_�>b�J��3�p=`
M���#�\�j~y3��V��:}��2t����%0��Ki�OU�Kt��[,]��\).+ͱ�����kO�=?�;�����,��G�n_�Lqn��v�����t�c�,�D�8'>�Yr�^�������"s4������y�˦~b6%R)76���Tz��� =
x�k��1�-w�fwNm����SH�
����Z��]om/��`���[[)��t+=�ΐ��<
3�#Tr�s��5�F�9�}��Xg9T���'%'x�G��C%���7��v˫�W�5x�`��f��J�Nm�p�f,�m�qa��?�����F�|����هY�[]U-g�*L�i�^�Vm>��V��ø���������`!�'d��Z� �)��a�&��Sǻ��~ >fk� j_ny	)��}�cN�;픟r���RJ8	��f=��>Q���[�Z��}?ƣ5�����4�e���p�v���-�F
_��\�⿪�#܃$��-�7&���)/����l���8��f�#{|�NEta�6��$�"�����q]:�澌��Q0':��?o*W�Z��Q3�L��EG��������CC�!��{ђ��;_���	��2͎�N�����۸8zE���2'FĿ	#)��lm�\�#|5���ڂ.��:y���;z��Zl��I@��X�L�����Mqj��A�8��mٌ�+������^�&�N�*�l����m�oc�*-��Av$dZM�.C<�d`�³�- �0��������F��ST���Y��"���5\d��)��e���*[Jn)"�7=��H���Q���lx��L5�{�/4��O�S���hd:�U0�U�^@w���V��ߣ����T6�㸗�FTԎ�� *U����CG��xc�>�9rm�I�86��B*�s�=���A����0�_�Z�:�T�7ͿP�����4���
�u.�Z���f�+��HK-K���A��@�';��g���a���œ�iA�j�X�oq���y4��,z��p)�L�\�X�Ź��{�!���/��\eţw�`޼��Ɖ�s~r �zL�g�*0��|;�,�����}z�� �JG�\{��z�c"�Բi�&�+�:js~M�.���s���LX��
�5�`̡�Zlk���'W�%��>�N�Ķ��>1!P�E�O��h��{�NI��fz�X���V	b1����,�f�!�I�������e�}�7Z;sХ�Q���H��]�/O�֛շ���0x������ש%
��Bl3IPW��e0��8K�9t��Ȼ��ԑ�=�\(d��ag'�ǴKw]渕8� 3��%5�,�[��i>���e��%��Pvm��ݚMdz^<��>�1�,�d_[q�y�#�%9����F x�P�K]�GW�o��?�%��1�~����$ ˓.�ԘPn�?�|%K�>�摁���<N�~¥I�������í܋���b��٤Z�&���q��{��®Da$!�E�հ�$�[P82����rL�A���|!��?m�`!*�x�F��>�pd�ܗ�z�g�^���[(Ƭ$!9��<X���-�����b�79�������eQ0��2=PgQn��1h�����K٪���@��4�X^^��0�i�{���!��X��cY��<�)�sUr\��o�jϪadA��� ��迴�=uU���[^��(=�T
���oM�xm����>Y����x�r�B䢦�|�r7�2m�r&X�W8f���|�|�1Nd�1!R����uw�x�AY��<���i���ߑ���eϲW���q ��JƸc�w�U�
ΎM�\��������w��=(\I����^���ʌ=S!T��☏B}�٪XN��{7}u���.���G��=u~��(Z߇�?-���ԽE�fqj��I$%V��X�[�X S�����đk!}���DX/�"H���z�&l���(�8[��P�7l��t9���ͩ�0$�zo=�>�[B���vf�匷�kss/G����H�R���GC30U������ec�>
��Xѧ �;L�A�A�i�I�${�k�&���N^��'��Î�*���z
V	��D�m���q��݋���-`A&/ٚ��ܐ��&ؿnvǞ�s�:� D�S��"u���AUZ�r�V;�� �iq��L�)�����v:�P�*o���o�v �Xu�ͧr�Ӽ��'W�<�Ap3U�W�Ñ���{M�w��1��k�
"vbdyd��'1y~'3!��R(�d�P�o*m����+����o�<ѐxo��?�Z}j���7���Y=�fy<8�L��@���>��@e:'��ζ6�*���_�<u�J�A3��@����į-�*˙�$�+i������)�4������#��;+d2;�u��o�����Ta@��@¨�^�T��3��(��~�>��?:��.��k��0��*�X�:C�#�ȸ��O˧B��Tsܥ��F�r�hY�v�<�U����e�Y�����$����Vd�+�����o��m�w�R���T�G�7�LRC�PwR#_|�]GD8+��w�W�{*���n{X�^ad�T$�"�����#)c^C7ᰉ�a}X@Ti��Jt�8�z
�f���`�,�m��P��yF��0�.�ڵ�?����D~����¼�<<h�s�0P�$�*����r�t9�h�[����=�:\s��pT�����S�ӣ1hP�Ù�a֪vǽ��<g�9@oq�bZ��Mźi.�A�\�dؠ?���^
~S~��i�;�W�C|�>&t>�1��m���*�9.?F�u�q�q#]�RCT����&� �u>Z�v0w�eM��)��oR�1�bF�)=�X:��O`��1�0�.f��"�f0�ۥH[��(�(�tJt-��k�" I��aU!?@}���@3Ӱ�d`���ւs�+�N�� ������rRo�ft�h8��4Xo���7�i��J��tLȣ�Cz���ζ����:ջ�G��dc��%щ?���3@���0`f�)r�4t��d~��kP���#�بT**'��	+W��"�Aqའ����y�,ZZv��pL��0��2���e=�T$q����y�����m��/�y�gS�C�}3x1ό�w�6g�r(t�����2�<ș�C����G���7JWN��|n�g{�=q�B��5�`�씑z��	I�<���8 �T�])˽��)�)���G�h�ɑI���7<.��\��p>!����fW�G�8����z�����w��Չ[��H�Ƒ����T:��,qum�����	����Z��>��,����a¡r�23>'KZ�rĝ�ܢ-H%z�#���5-�ҿ�> �T����Q�)ҽwY&c��9�5UZs��L*b�$���/�^��^vs�<�l��J�r)�'��}4iZ=������$>F��;���"A̍�-ܼʡgy�_	���!58�oמ��`���sY�#��Y>)�������8]���ZD;���:8��U�1~��V��S�P��e,���*���n:K}*���Y��L�q�D��`N��6A#S���j<2A�SF;&T1�N���
��R�e��bH�ֈ�קྲ=C*+&��^ƾ�~��I�w���谶 �u	�`g$��[�3PG\ie=��Uޞ��wVu8��R�PG���#�ۏҎ״�B�3�W�Yc�L���69t�N\e%r��l{0���=}�1(Ѯf��w{����Kv�V��4\FN�L���r�c�u�sd��W��C��x���]�
�MS�|���w�M�b �b���f�����*��rc1vn��Y�۲�$�O�56�D)T�v'Jo�3i�Qm���q�6*�h��%|�_�g�ل�K͝W �)�6(�v�,��z6��2���{(��I��m���^�O 8i��[�*�[v!S\�xY��e�v��z�W箪�D��Afڬ�j�)���܍��)����PMg_�~(~3��+f�Yt��;��j��o~	�ŷ�ڠ1)۩���]�;J��l���=jq@��k1ws b%{�����0v!Z���}�v���OC�uc: ���'��9Fջ�l��yW�i��5��M�6�w5ю�LP�fZ���$p=3���'�.������	A��s�x0#��+�g��H'Hi�  ΀>,�CY��0����b�yO�3b��F�Qt�㪨�gJ{�5�*g���~�}���|N�ZXma�`�(�JT8n���m,�V���}s����j)��l1�Y/�I�;3D�SĔRaD`����nz3BN��;3	9ly<��h>/1�����kd}8N�c5�42��EW�ˌ�Z�ī���Z�y&q���-ǽ�Uh��G�F�=��E��of��\�kث��_@̙�͉>�Z�xT?�}��'ܻ��D�)�`D���`۶��i$�A��_:p��^=����P�"�����2.�SrT���X�H�6���P�sO�q����XJ$�5�I��˧�?��"*���B����1�G�>�O[v�m�q��,�WlT�c�]���_
T8���a��,�|4Lut.@�O3�w��P��K�q?Q5�7�7��]��?S�rNB���g0{^��h��X7�J���Ύ���3M�����Q�dY�~��%#L��;6��v:v����C���=E��9\m�n@��/��Ԁi�?S��2�Jrm�uQ�_^��v[\��>�C�M{���V���PG0�g���K�_�����A���>ȴd{66��OSe�LA�uw����CQN�-��Ī ��%�>�شp��Ʉ��%m�`�8��;��m7��7'�j�*��#��gi^�瘀+q��QW�N_Y�1�N�� �x(�Ϊ7Y����/"�t��뼎)��Mr�ԩ m�U���f�_$��"HC(��%V��#R5ZAT��:Kɔ��^r�d^����Y����9�
�9�tJ~��3=]_�^"����(��zB�T*��;R��F\�����r���J�a�(Tm8I gKyXN^�6�h1�H+k�0�?�p��q��Y���z���#�I�)�`t9N�wZ}��Wk� �!�~�G3GLm3�N�5���k�C��é��xw��TL%�t�����-�"!��|��� �&RG��"��e��8^���C��D����������i�9����H���s�կ Y!Q1):�F����2�-SQHh�Ӄ�1�T<g��i���]�hti�Uug��Co�X�s��S�!3����k;,�R���Z�Y��$�R�����KF�I$wG��?w5�	ʺ�<�r"�m�������Q�(�^s���[gb6,)⺜�G���R����Dbm�U����R�Qn�ц�[B>1�h���2��}���[J(�|�=Jk����$F���[P �wE��Du
[4<���H�P	y�*�x٩����#`�4����Բ��<�1X~�o��
j�'�$H�g��ҮC�[��Ws:����$L!���/�.�I�D9���^}���a?�5���I��J~p�!xz4�u��\��;��Q�FwR������3l{�f��?�at����~\%�N|S�l�ԝ��!�o�-Nв�ow��p!�sR�)=I��-(I��Ġ���7����[W^�|r[d����RNP����-u��Uc|P.E���h_����W��y����'D�zk��-�v�&���M��$]�5���.l+�'�/q�2�֭2F�Q�DG(I�U�8M���Ix�~�Yu�DR�Z �3�^�J"���~(X@�yZ���6Z�`M9nYXz�|���D������x�v�����6�禿C�F`�^�W���~ZR̾��kJ�V�Y���Ƅ�A����m�=y���H�p��◰WQ��c�`X46����t�����}���&3@�����[A��]Bv6-��f؋4vμn��_Ќ��u�JC$�7+��҅C�-���oS\�"���h�>��n�����z��'��gl�_���{��ώ3\�9�a��N���e��UP���tCR(�|#���]��I.�e,ўf;݉� ����Xb��G��rA!�G'3.7��q	�b(/���� ~,	p���A_;q����풒kb���T�w
�*�QI�w� !�y\�I��e�lM��y�Պ`�����J�;��
����� b60'�#���l�]�?��$k���wr�Rm��]|o�K�C>(J��a���o�9d�	̗�fq��L��/�,�����9U������>������U;��ͬ�%�V@j��+ìeD��5����%�a�$�����c|���o��8#��y������f#�#�W���
X������D�g�	P���^M)�i���(�;��5�/ؤOvR�� -#�/�����#�b��z�Xy%/&lԎ��f�Nn��~/�?E�dUJ�܄���0~D��>�؊��m�f����<�I`<�r����ѲݨA�LO�\,V�����ރ�;����>%MAa�:�`�,�8[��QE�m��gQԤA&1�_Xb�6L��-�7�Ln��	9�M���/Y!&�B_N;�)�>ۥa�"$��J�*�X�P�h7r�ER��� �N��^�t؋'�rZ�t׻XR�;��_�L���+;�8��`�����8X�n��&���{\��|S\v0M�dx<U����T��l������6�m�JL��&���i��o��
����ڳMÚ��T��3����P���,Ё9.�DX~�-��U�0��+ 0{�k�O�f����k�|���U8/��.6�==���8�i��!��8�Y]����� �� d��� ���x	�4<X���QJIp��W�������3�#Ľ'�w$��������kMr9�>H߼��k{�|&Y�[e��{������]4q�c����C����ʒ�ȋx�I�c������-�w�����ճ���������D��u����ɀ�4�:�\(7P[�{<2	luH�]�h{��>C��,�_�F�k&�R�1�Hh9dϯk��X~��R�<�\�ѫ*�,�b����(��	g./W��U@V%gY*���������3Q,[,���_�h�7��x�b�(��$B��P4��aEvS����]M榄H�POa|Ӂr��fm���?|=n�!�8EF�⨈ڇ}���+����
N`�Uj��"$iHuӒ�-�B=��h}��a��5�'�����y{v�g�͈�y�M��և��L`�|���Ą�0U���T)/�p�LW�L��\?x~{	iH�_� !{�*����|k!�;"6h�����j����-"�=֖ΥW�z��մ.�b4�$b�����M���7���$0�M��|,�Yl�;�"�Ʋ�0z�o�~%�,ً�aC�
A���/wU@��n���p-2֧`���0}y\{�$(:��蛪�w	W��>�g�jlPz l���ԝ�d��2��C�%.��QJ�~]wx��u�d��)l5���r�z���D��'�薝��N��lYa`+�]��_�]U�N�Z����TI#��9�����S&���-C�c9U���K�O��{)�{�U+�t����S���Lsw��� #b�m���XL��/�-�.�(�x2�8N��{��%�z��c˴�~��bʀo#��;k���o�f=�3����s�(Tq�9c��A(J�a�	�f6��O&�4-ݭS�pF�Y��j�t�}��Y�s�_��C<�Ϛ��`�LP�tR.!�X��q+�CVR���ާX�pi�8�b}���E��"1��"���6@��m�A��Z1����^�Ѳ�����_/���7k�
�/;"�#���I\i��9�����&�$����9f�� +�K&r�a�b��x�_Mv���P�/��fg2�Fo�Ƀ��4�́<�@�t�����k����Ϊ�4� �H~d%Z��v�ǟs�NրM9!�N
��^>���G�.��W0M%��k�&c�|QI~3�*�^b�.�[��;�8���������Ra�tU��)�4Yf�x&U=50�$�WM\��yH*��E��qC�:dX�mo�|�����r���-�G�.�Ot�V�^ݫ�e4XU%T�C�ɺ��7�8�1yu�[�J^! �Y�9׀=�9������2���|D�(j��*ܒ����t��,�,)�eB*��0�H�J��D��H�|��h7O����0�@#O���#�u�v*�k
���u�h�]�}"?Ц~�w�����ԛ�P~c4
 vZO�P%~XYp��Pn�^䠨�Ͱx���SȲ-Q3F�V��J����Qe�%�=�q6g�h�y�5N��&�ډ%��'��f�\gq��t��c���e�ؙJ��"�m�|��6P)������4�j`�+}jҾ%��΍QH
))�7s���ϼ�#o4�|9�c����bԚ*�J��**��q��c�]-�;���.�O���`�}��zjj4�	���H����"�cQ$Gȷǂ�e��V�c;a�d�sb�b���ś��I�pm�n�yh�W��X�ݥ{�t[]��z�G]n����" `*�I".(<�w�ܔVjN���v.��ZuE��B���W�9ޮ�X�b�5޿�_p�U*n|b����p�>�k�m�8��"nzw�,X���O^����� ��������`L�8��>�r4KM�{O{y�i�yz�sؼ��d{��Х�i<_��`+b� �=�[`7M3;���(.�!���V���9�]^��d#�o���N��h����x�"�zb�!�M=UxY���([j��>�t���
�!�Q��	r	P������q�f���*ӛ�Ų��gY�<�2��z�%��N<}~���E�lʠH��
��ֵ? )��8����sΡuv�6�D�Q��\�׍� �F�>����x�f��r	���	�:ye׼FIh[��=D�=C�e��@�8��E�T}KB?���81�q�(���U��=èbӕ�e%��0�`�Q"|G�;���:,ްQ����4��Ղ�P��9����Ƴ��y/���S�Ůkn�07Y7uN�ۂw��a�`x�a�CfI�!���6���!�q���hp����\��/@���4�P#D�*R�kAd�dƆZV�g1ʮ��Y�U�����%Ų�_ ,��	�k2�m��g���ǝ0�Pn��r��=ebu�`��ZMC���L�c�v�Nx�q�t���UĄ�хKP���w!#+p��T|�B��0���#����P�"a��}��A���UA�C�	X�M�
d�\%�{��;���AW6}C�#�R���xP4����;,~5RAӍ�Ple0���q[���`R |u��yv���D�����JH���T	���2��;��Q�M�N�k�_��L?�*�imߺ���*j.ٛXG*�VƦ1������,}��vn?vgo}Ul�a��W�a�u�� ��RS�"�/�n���	�#��H<p�u8�ɜ�d�"�KQ/T(��xiլ{G��9a?VU-R�x�?��()���ɧ��-<�HX��t4�]|-f6cރ�T'>���8<ҷI�o�R�@*>�0&`���Po�W���v�K�1�~_�zE0��8��}��=����x]jE�	��Ki]Q�.i�
�2a|�M��~��=�ͤ�T�$���[����pL�����
��H��^"�Y�Ҥ��(n=xAq��21��?�8gU�x��p2����<bV��Y����7!�����|�^#���ެj�b�:Z:��-R���(��������JL17�Ӆߎ�h8�U���B���mg�BE?-t����z݌H]��� ��I������0m��h�����7�Z
c���8��M�[w�i�<F5֝M������b�t�|��6�.���D~�x;�d ��-�^�5��d���D�k4
���Cu�FM���7����Ȝm[E�ly'�3�X��R'U������AX(�y_�~@�v��	�V�u�L�0���?^�U��㯫� ,����zD�"	�k�$�O>Nq��m[V�����d&��NF5U��4��h�:�B�)����vb ƌ s�;9M`�؛�L10�~���`�Ml�\0�J]�W޸Ae�!����qwfh����D��G᫓@4?��~RoI=�C�xtc��ё���ۊ�R����[��8&��T_�9�U����'�M	/x�Y2c�X�&u��`�zs.���4W�Z��*�;#o�q��So���)ݠ�d�݀#$��ou�:��qN��F��)�N�¾����Y�Ň��>&ڛ�|�ƫo����g7��8S������U���O���V���=�WzuK����hH�1h�� �'Gr�ci��*�����FJ�J�=Yk�����8�ţ˶[�TV�B$o�3J��3�^B���lյ,�׭��R�|���0��<JyU6��f�����z�&��h�h�I�6�%�J>��̬$Ԉ<��rʏ,��:1y䒰�,�y��
�M�f�<�WbG�P�� �q2��Ӑ��`)���2�ƢG����rBXb��"\�!�	�Ls���@��A�7}��HU��g�jl�vҐLl�/�6�9�ν�]2Y]�Z�2��rB)i�C��%ݛ<V���"�E�7����pF#��ڟQ?Y�
S������+_xO��T������o���c�bԘ%3Q����	u	�SOm@�p��$~�����T�sG��܋�
Ж�nlٌ�������2*UO/u��Zu���oLb�(�W�;��|�n^����vQ6���E�Gů`���
4���w�:^(Kѣ���r��u��Ok��K�̈́�l��Cd�'��I*�fΌ��h�/��q*Uv	��̎+�+�C��? �!�N)�]��kM|��bI$��+����VT�f<X"�9�6w=���*�E�{�R�#o�����DኃF��Ћl)���(����iq����7wY��S"\F�3e���e"�j�����4,��׸�X��E�t�з=�TgC��cǯ��[睂�
����#I�lT�Ig�+�.r(��ڠ��vD� � Z��1�E3�S̐�*m��78
,��9��4����o�"��Fb��	���k=z��8%T��&r���[l�I����ܓ�:Г�J�j�K�Dʚe��Y;�T��}@�1��;sSo�Lٟ9H�u��z7�X���XB#H���OA�2��{���!Ӷ]�|�蠎��vߍ��$��{d��N���VOW�N6�\3j���L�E�po�(W��5�*4 �Sz)�8��e�t�`.�D�F�{"���D�Ǭhm��ClȑO�>����F��0+[X������$!c��������`��"�����1XG�ț�<�?�m�9�:a�T�(�)���ż��`4T��L�)�t���l�`�՘�-N���.��5��;&����,ۣ@�d5ZA��#wo]��g�B��]Mߟ�٥�Lfz�����!�8g�<���g����V#�%0��j�hfԥ��a�n�*^z��� �\
�tg*��ۅ�H�&!�h7�c&���gl��v_�%���[���Ohx�~o��X�OIr�}Y'��캶��L��3X��= j:\�*f?���WN��CR��%.����ru���a�C�G�Dv������ߤ������l1��9��0R���K-O��54��#	�w�TDЛRLon�YyK�OU.��]a}�O~�`�JC��w"�{�$qHS�΁�E��`�X�e_
E��T�XJ����Pt"Uອ�xȍ�G��?RΑ�=�߉B߫43������+�(<}D48�<����nI�X� ��/�0����3�61����6*�\�^x�ڌO��`��q����_�[��ƒm h9bwD���C���v���b�:�s���w�����P��z=�îs6��a�
M���5"x�p��]_���4��z�@�cd���-���x���E��.���c=!�.[�čn�-iUÈ �`G� ]g��X�ChíH��St�L��6l�������Ep��)Y�GFR澛�E��詇x��^��>e�z3�1-����!!���c��/$��e��&�Xo�3V�%��SB^+c�Yg���E��C�dI4�~���'�����]��h���&alW2'
���D±�e���Ŏ��ꖖ�-�����.)XѦ��L�P�g��"�0�{[�m����74�����+���u�Wm�{d3�D%о�����`��js�y���.�6bW����t�M��t��� ѳ��ӽ�##�����A���r�
�{�"M�=�q��E��b�E�0�܍���˕���]�#u��04`O�eN��ˀK���@�u�c���A�8�C�����sά[�r{P�=�~�����8\8n�R:%��D��ҝ+�M�qg]�;�#) ��՞����T���	�[.�W=b��9U�W�3r�X������������I7�#�h��=Ў�ᔃT�!W'�y��kQ��2�eꞃ4��O�L$������Y0��z���W���>�g�C�kU��kŁ;��1�z�+��>#��5�����s�>t��Т�+��?��f/��F��`��0����,!Apj[$��l �*
o%8?Yt�gy�m�ED�4)^؀� nyi�1���D��Wu�ȗ�I�ӂ8����-^٣):��t�y�6��a�q�OT����~��ۃ�2�W�{u	��&'B���h.<���=5�?Ņ�%���27�F�b\ 	�g�a�������6�ׄ&hW�c��mf��G���#g��6��t�_"9��0�n�w�y4;-B[����Թx\{M�渨8��A���7
d��R��Ŋ r�vv��zOV(/����CU�.���_GV��[E@�L]Q�M/�	���W�L�!YV~Z�	�4N�o2>$(�ID[%转�}`��]z@4����B���,�ͫ�E#��80}�\?bQ=,+8�a.,$��Z�\!�{�V�]�=��f�g��.7��4�3H��`׵oS�Sٽ�v(���R�8���E=�t�s�]|���6�.ܱ�\@�ᆎw+�PCSx|�x��؃��<'�}3��۽�G4�+��Dl�_1J���+�}�h]8j�Z�	�{�|�WH���: 2�`x�b�F"K⤒�D��,�z���W>�YJ�ݣOy�I�՗0��R�N�S��T�.{�JC�M�5r������؀,gPH�p��jq�G�m���Mv#1�����)�k�9��٠~��32�b9]E\G�<W�j�]]���)�A�]���8Kd\s'{��%��˟Xd�2f��Ϳ��OD�d��`��z]�)�cG�5C/����L�)o�)͒��J��G[�<?9�|�B�ƶ=�����^V����&7s7i�{�r؁���v���{n��O��p�<����RCѹ��D���ɗ��T�~�&&{԰HY��b@����ڭ�-�5m�#w�D���f3߭��\��NŬ��Uܽ�3ua��Q����Be��%M�E������gR���ގ�ٿ����	��xX����Eו�H�K�DR��gP��:�G���ᄥ�'i97>��P�V�YH��8�]��Z�����G �
�9�j����|����� #�(��6g�����{��=f�1�m��U�U�=8w vL>��� �_K�8��=�6����;�����p:�]�d�3"C�����A�0O|�^�_U?�@����~|o��E�H��1u��;U�3�7Q�R� e+C�0@��B-�,0�f������4���.�jXR�r
o�.D��Q	���)�|v�>/٘�}�&":�V��d2Y!;��Z">k�UL�OL)'?�W�ـ�r������ZW�K���!��Y���`�ar��֕(輜�3�l�NF�ڒ�Xj�I������uu���4U@@����xf�"����]� ,ǚ��U���T����\H��i(JL@�j���[�](-�X�Yn24�>��[H2���rcb���24.�k6���$�27�@Ÿ�犒�!���-���)��6mj��i��'!�k
�m��!�>.�3��\�3��P��,�S�&���hS&�_�;�����+:0E�2O���Ð�z�B��PDOz:�"$3�ZnV?�{{{��H1��?�@�����u��FDi.咞M�ױ����N��n��J��#�����/������24k���ICxn��i���5ݎ��,�
Yx�>xH�t0��"Ǿ�Cgt�2sc���Z
p:G{%������"���Z�vB�Fc����Hߐ��;W�9�}�?nW���l��*ָ��������#Y�(�b���b���s�7k(}�h"�0��c�+���q�v<�Ȍ�L\Z ޷߮F>��J�P���hc�eڂ��L�tr�Y'�@5��Z����&G��?[7.�I��ty��7g�������i��c�c�
gݧ>CuW\΋?����d�-�N��n������ �ho0�|g����KTm�>��!����踕Fh�����p\�8R6h�7��6i�֏������@��y^^[��S��۷U���a��	���1���ک+��~;��%�\m��<f��A���)��L�N��Ы���Vŧఽģ]�g[qT�g��<����ˏ�ia$�?���k�TH ��Pd��o��g/�l6�<ny�T�9�H�����:�g�J6�/l�V:0A�C���\0�\���2���%�E�9�B��Ǎ�k�����g���~��nM��G���m��ğY��� ���
�͗{֪m�&�۱n��6����D�χ���,U��E���l��T��NG���1���Ŗ�	k�(Rj����`��y�u�S�ˢ��sѠ�+N��f�o!�<g�n�2cDdO�j�OWɷ� 壿�I¾��"��#�=\9zSjҗQSo��z��������U�4�4��l>�S`��_b�b�������ϸ�(F���Mj���Ξ(����`F�-׸?�b������g#�qco���.�J�r�������*|#C[ލ����r���x�=�����S�2^ 9M��uuA�e�-h��+aJp�[��`Z�7-�W�I"s�mjHG�������oM5�=�Uz��7�m��^�7`�a6��s}T:��2U��<O|N��H��=��/�G0��[
��r�I���xݲ8�?�Q`3n	�����R��)[ƑRچmS�赮���(c��Xgu%�* ~�V�ڻ��ꀛF��!�C���Z���:��w�P|���,�/P��n�AR���>H-7�%@�V^���5s�bĬ�X�3mO
�s�W��/�J`�Io,�$~B֜�6�=@�ҲLᆘ��S&H�^����.'s:�b�
�ⷛ���#���U�n�q��f9ɑ���Ӆ��b&�?�](�ڻ���6p�6qz\*��Um�ܲ��-a�.��S����:�x�;���=�p��P�2@�w͊n���T�b�	�VwQ�V# ���7���}8��j����h�����D���_U���=x�+.�a&=S/�=�m��2�F��܍mA,�J��(�Ѣv���o�i�&A��2�N,{��u,*@ҡ!���rnJ���_v+҆����&Fɨ"�~�5�Zg��/��r�Dg>��몁��`.@�cA�5��誎���]���#�8�U�Fڬ�����	��[\�6����H��v�c��6޿%3�U���̺D1�`���:�s�Jf[秫Ό��F,��}�Ŭ�ml$QO-�ٌG/Y��k������$ ���S�Ŋ*ѰȲ�0È<�B@�e(K��W]�O�]:=gB�!���o�"�V�G�� W�5��S��s�����zU�M��.�cp{�~F�$l�3���!�7���m��^j m��7f�V�>�gr�a�*�����:U�:V\h�Mαߣ����������f�>���\dY���:r�o�C�݁��o�I��G�3�L��ӊp���@������W�����c.v����+�hm�q�əoR*3��E]�wq8cS��V�>�aҚ���,\��|\NnY��_�99�N�(� �]�!��^z�1Q��@hæ�x_�m(MU-v�2�\Dh(��9x����m��L8�{��t�ס���5l,�p@Ҋ��2�4//�&~�Z6 ~�����B�JkQB��$-�	��G\ƾ������eG��V$��9����o7���|�*�eD�������h���gx�B���ci�*,xq�D$p\X|�Wy{��Y)���u��o[{����+���S�k��?9A�9
12޼c�z�(Rk�2��T+i]Q���y?`|&� ����mc���_��������L����4�,?�
\��w��o�	�/	4��Y��p�J����"�.^���X9���C�T�����0]�!�4=&�qo7+�n����w�'lı���υ(V��M�i3X�0T�?c�(��a������!�� �N�Snm��`9Mh�u@�l�!�&�-/�����U}Mv�a�th+2 ��A��#�u?�/��O�prklx�*ci6ACY]>�H�����̜ ���.d��ސX�G9 �f3I֛�n���i���!,�	h��)���$_͙��P���Yr?�� h:�S���DMG���W
b���������� ^��i�~��LRŲ�����j	"5�^�I::���_��#M��x��i}�JM{��E*+m�'��
�JL�ohS��6i�ty���?�VO�!��2[��2�V	d!�cZ��n(^
BwU��<0,�-V��-�����)�1̇�	�y?2Bb�b����8C���ݵ��80"�5<��2Mr�R,;���k���i�>�%���h����|�w� �sG�@�ۊN��L��jk_�ag}M>��A��H���DH$L��-B�Խ����Դ�5Y���yd��V>�5���)o^[Q��%n �������e`��W�D����*�֘`8�ڙ,�f�c�&2Y/u �u!���PȶP��R'��d��uE��!���[� �m�GV��McI�?e;�:i�c;׳+Ⅾ35�(�44���>���M~�2k��=/�ƴ�5��K"
���H<��2�9G����*ޒ>�w���U�B}
��>sÛz��\`���v���;[L�6��FG-�����W�l���e�=�zv�qh�	fV!�8�`=�қ��Z��Z\�e�((��6b&�@�:������n�aat�/�����T�x���μ��3��9��S��E��+���Ф��m^�C�{Ƕ�:)h���3[~��>e�vM�F�v.gT���&k}��˧5��6�V���� �3�(���-������in�=��^!��G$�2�h�-�o9	)��Q��j���w:�lC@���������v���X�6C ٬�����#V�JOg�����(�ف�(ͤ�#��G���E��g�5��\�6��R��J�CY���b܌3=�-�k 失\�a��[��L�C�N�A'!=�����V��w�M�3�?�B��ژ��ˋ���P4���8��b���'"n����r�z)O\�����^K�	���{ݲx#�S���(�F*؇<�^�/�6�F}U9�p-���1�<�r�S���_�$GM�VA�ю��}iN�o����e�Q�3fT�D�IN��%���� �D���y�dD��'��WADp��>E��u�X!�蚗r��x��5P��H�}�"�:wX�C.7�u/�8�I-+;KO�W��Q3��ŇiT,�0;S3�h�����՞��A�����c��j |�Y�[��@��R���X��)�f¨�~G ���gq��bd��u7����x���a<O����I*�����)�_cҎ�XR
[t黓�K������XEt�H	��/ҍ/1����V���hͶ+T����A��33���ǳ�M��w<^��<��x�0��g�}m}-�W��_��j�?.��?�]��e[�d�t(ek�^G�19͞���B�s�]�S8r4y�%6���Ւ�\e�ͩ$@;�Ƙ������K2�Y�Mh0ʨNڸb������P�R\)�^����P0N�T*2?��T���1��fM��ӏ?o.�j�1�Ύ��u�&S�-D���@1�`�&�P��+@Wڠ~5�$���V�x��Mw�\�Zl-n�'5.*��{�����y���ON��	.��f ��c���C$�OI�@�ٽ�-�s�kd�[�O�}5�y��6?:��ujyNasn��G��#]�崩N.����'�Y�7�v/u,�+p���
���Ղ��S���"�ƭ�����_%<6�hcxFrsg����u/I=�@�d�"l֍�z�#�uR��<Q;�;�}k�Qf���y������%���e�,�Bj�h{fm��R't����32�d�����i��z
-�L^�v���1.XXl�6lZ4?4��c��|�S���|#����j-:~��3a�\)���G=���D���OG/��4澡��C��5���sd��?�]NCj�h�,�K^ob|��W �)�?��S󮻒))r\<�zx����<3�� �[��6�x����	!��K�(�#��q��x�RV(��^���b�!$��*Ljw<`�:���-�7�~�tR7�!�3E�F"��ꬲ���'c�]<��X��0g�iU�T���*ï}_��u!�:�,����};�����V|��ю�4�k}��=q�}�	�ߟ��c�S�3�> 䥕|�C�b��z��9������ƲJа���%Q����Gq��ג�α�)c_��B��f���zl��-��|z�30�LS�h�<(̛߱�MT��
��(��A�>�����j�����k�{!(���9��Jв>���[��<@f���X��-�|z�-MNԎ7�{�����q��6x��`u���,�1!��v�ɨ���Tlfq��w�KZ��'�{�����l�P�$C���4�`�-	^o�wDbW�#��G金C������&�/1WE�#�ۓ�@!�mg��&a�>q�Ɇ���~jW�{(>npl�<��Lt�5�ι�嘃M�*Q��Dn��hXb�d]�eE�W�⍵��B�EM��e��N���9r��P�d> �M%�>M(,j4���O:�{��� �lW���O���?b�6Nt���j��_!Ćl?��q�����<-�D����K�|�W��E��-Z-�3���E�� :s�?�x��/�u��E�y>S����LG��q��l�;���y�!
��ְ�c�ԟ�-�K�yר�3�3�R�� �M ���s�uY�W�[�)X$��=L�V�G�����ki���_ޝ�-�B��[B9��G����r8Q��#�C���%6`
f�1��|P�Լ׃pK{�-
�5�h>D�DiP�@�/��h,e�Z�uSTkU���N�F�H�Ǣ{m
����C�U��
u8N�h�2���{
��IG��H���r�Iԣהּ���жf���H�����.�R+��G�0�5�Gl)J��^�C�ս̝��%��ѐ���X�Qh��_�Ӄ��Y���p�ba�sgk�<��%���kx�����{+���	*�ʑ
-���x��M�K����;6�1^�qV�4ۜ��<�]�Q�87��I���Sk��{��>���c�BbB���ҐRNF��&A&������V;&B[���\:�'Ֆ�(�6%��uL�[%�=^�zWYt1h:�9�Zf%'X�&�ذZ c�e�Ux�{��M�㣺��bA CHk*��gOU�qõ�#��Dy�"��I2�㋁o��Bq� JV.4�ܘ���G�T~d��e*��*�.��.u��Q� ���s�[���C�zW��w����-�_�Ċf���m�v� �t�v�f�P�g�<�i����N9j��P��,��E/�P�b����7_��m��ڶ��At#�Y������o���q��A\�]�j�0���I0�-3\f�X[	+&;.�U8���Y��iH����6�����rMG�/�B�^�����o7Tw��bE�o{ӄp�`�;_B ���{��f�+��Mw4ց
�D�>V�l1� �L����LF�"�z���|���R�F#})�x�U�*�%ޛ�K�^Oq�}�ȫI�坣g;�-s��o��``�%�H�74�䁳��|�_���W�ơ�p7�f�G�S_��h{_��MVMf�k+����p�LOzH�����?۵��w���<k�⸑W�1z~/���߳)YL���g����TBY�έ�F�*b����i{"�nzb���f0b��8�4�2�n��A5^�]��A���X�i�����O���?�t��G�K��;���f0�0Ӆ�P�	d�`/=����s��m�՟���v�%�%�1����-R�P�Z�����������\}yI�P.{��Cցg�Ք��J�oj�Go+Y<B��HC�+�� $��2� �����o��pvU��Gf}�h�g���Sչ��&�V*��':,B<���G����\�ף���N���Urt�3���$�t֔hՅT�
껾�+V��P3�C>x˫0���Ϗ�aU#��%���%Qr�6���P�6��YK��Cz�������שC�׷�����a�*��A4S�E��p�a������Ny[i�0(�o�li@'I ��Їѫ�݃{x껄�Q|�vЇ����,|3�f%�>,0�f�)v��L��[�`ԛ�C�w�T�B	��>P�q3*��FAXel�2ŏ93p�$Ǥ��:���z0��b�2Q݋�p�b����A+Y�z2�l��1��0gi�u_w��	���:2Yڝ��&���I����D܊�����BB����qx�qbU�Z�`�I����(���y�sn��W�������7��a��?�'�̘N7��	�K�$�-{[H6s���/@���vO����=U�\'�=�<����;�����p0���R߻��t���4r:&v/����`�>�Z-r�B�R� �����@�]x�ka��K���U��A\���ʛ�TAx�v���:�=qA
:u��>Y���u�i���|$�'��e4���,��Pb�p��S���9�6�V�5��(/�l&i���숟�yӶ������p����F�C�O�{����ǦbI����?���,�)MⰮ���/@+]7 m�~�b?�mQ
�	�+S~��(�ޠĶA'k��$�T�j/��sϲF��P���Kr|`[H�WSٸ%�2��D��C��;Qʗ��r/�����2����őS�L�V��EI'�pI5��u���o��W�6#���L�5&��>1�����F��Tz�@U��)_�[�4�P�߬ޖ��E�0�)�r�����g�dBD���|�jg2!`p�e�t��2/'��
V�pݡ���W̍v�d��!?�����q�$���^��(�g�Al+��c�Tk���Q3GT�
9�dP�(�5�D�&h��W�:��ϑ�?�(����"ڢq��%N�Za2`�����p�nQ����J7��4�j���t�q~#!�)l-K�hi�D��,p�vF���j�u�dS���`.��/='$�%�� +l�^��^t��3[���)z%��,�a���ʸ��p��J£u
#�U,X`��64Z5˒���8�h;�)�)��������x� nD��d�ps�Kw6��i�������-����f�S����=���sDI���ς0/�3��$�
# �U-�h6��BŇ�R R%:��#w�k}�ǱgJ�&M6��<��Nen^��f'psn�@*��V��s����Iv�Rx�_�oZ���#�J[�.����5#i�O_m=���X2�$�����m�Gѷ����]�9��| �Z#_+�U6���+d�� �;r#���M���1���ѣ�!4z�W��afӼ6M��g.�Fq|Dã6��h:����ڷ,u�-����32u���s{\=�Q��˼+Xy�V�k谔�ݥW2���?�c��^2V��ckhAP����-��s���V�. E"|2f��#5����{����!�f�B5��7�`9��
�U�~�zJ��fо�m\���Z�� Y9�iG�e�˔b���Kw����`��5{t��n��b�.�Ub���KuԹ���|͇O�᳚��a��ߛ���춤��"?ِ��}����^�eViTw�H
�DB� T߼v��t��B�d�[���4f3�`cX��b���6��]���|�M r/�4��4�,�IEi)2�N6X�\]��k���9�8IĲ����	xBH��-ѡ@/QR����O�V����Rgێ�Vh��f�,O�>Q׹��W�6 �T��0���Դ���xIL įiÿ+��<�%���KQ�2�8W����V\��xu7�E%��/)]_��h��,ps/��m��_��4���mt5�p�����?�Q ,�~8�����N���0`��$�SRd�I����+�ኯ�):1w���)�WO$���fj� ���2����-�i���C��/`���L�Gk�E�]w�a��>���"�vO�����X�Lg�������w:�>vD*�9���/JD���
VQqOPeuV��q��dH��F@�bX I�"R�4��!�O�լ	�<jR���p}%�~�q�C|֊vv/�ё�e������R��pc��Q�-1�$���6��L�����v�Q�����H�E�"CXt������lt1�q�݄?�}����K�r(
����2�?��2�ZgW5���\s�X;�#���1�����b��I���6�t��X��º�9�U��9��m"��n�Z &�Hܲ����M� \W��'��{�paY����t�@48�+�?�:�x��y�A�Oo�(���;��j���v�>��:�h~S1Ó��;���=/y���=j��u�g6
#��O�=��*������K�z���*���X�#]vw@6��l����q����z�)mJ��N�R�_��ǝ���"O�4�D����d������+(�n5���?���x��,��ɘ7U�ׂj) B�LX�~�\��$"M�K*vr%d���/��,��XS�Y��Q�h+��{Թ�b�c��Tmz刕�t�3nO���Z��H��⪰F!)���E�:�{�G(�����%bq��{VB�N�6R��\���r�q�NZG��ԸV1G�#�1�~����_�����2�tz�&�q����,�Rr��E�P���F����x��y�n��>��آ��]�RWX�>^_�ʀQ0@�j#&Y�HZI�oղ�y5f�d?�n���?@0�2E2&ʥP_�T�Baxvwj[�p�I{U�dкTyw	j���Cd�&��zf�~9�������si�ɐ�	�,��RmN.��� ���m�Z]�GK,0�2�q)�y(����B#[y��ސ��懧���QdK��)X��KjN��Ӽ���U� I\U�\ˎ��(i�
�*SY����4�5}�1�/�}���ϋ�ɨM�@�2�B�Q�$�$�j�R�e"&b�Z��A��Ј*E�G��3�ė����r�{�;$i��@2g�г������������ϴ����{���)�f#}h��p���:-�@�`HͶQ�������-���>b�E�:�W���Rqr�;��M��B� �ulx`$G�~��|Y&��֡IN�I�$���.54����P�U���4���y���=��3�%�m{۶��:fj��9����2C�ۛMg��2X��]U3�U�.n\͍:�#�_�є3G���!D��:q�D����Z���I�M2	�\���d�:-��� Ƽ�7$�s�mcMSyp˒=)@�p��F���U��-,�t�<�ß_�0�iq����>�Vߦ2�DˤN1Q1	������˭�4�?D`�.�7�� �x&v�4=�uI�+5և!�r!��u=exT�S��k�s�Y5��D�(���J���-v"�*�� �8(���:(Ɨn��ᔪ�38���w<�q9���uު�.��]�*�R4q;��nqv�]��{U�����$19O	�.���r"A̰�M-\�PV���S2��PK*�W���v�"����֐J�ȹ�68�?�g�h-���be��W J1Z$9�ٻ��#�yd�@M�Dl��9���_��]f4?����M���F�_����?<�Q��̷��g$uLSIhO�D����ܶ"�F�|yF��#M��ML��J�l0���П����m���+�fwm�a��)�Q��Du�T'Ky�kW�8P���~�k&�&���vf�v�d�`�p�6���v��&75� �l����+Q����RL�L���X���d,n
�-�;��N �3�A�Jes�Yךɑ�Wn
�n�/H(��`������@@=�g �U���?rg��Ww(.9�tR�3e���*0:��t��<��n��C��v��,o�6�^�-K�$=}���C&�6Q�F�����ק5R�f�ޒO�YZl!"��g������$ҼK�����kB��X�G>`�K�#C�[٤������ g�A��]�T�-�8Q��u)�p����b��5NKeg>���`����F[��T\�s��+S����m3k�6d%�^�������	?@�>� JPT�_F���{��Ғ��C�,)\"]��4�f������O�Q��Х�R!�I��ʊ�F���4ݥL%΃��ń��҈YV�a5�T�=e~��w\=�������
�-9y�Y�g/�d\�<M�A:$�(jD�yU.�$?�ѥ'yx�h�+Mק��WB��rܖ��;���r�Z���Q-I��*W=O~!(P�Cbx���΋2jd�g�,��U�<uЦ�5
e���)Y?�č�7��>%Th(ׁ4s���"�h�懘	�B��ܹ8K�4� ��M?��!p�Ѹi@�V���P�#�m7豴f��>�r4r�\�ۯD�!Fa"L���P0;�����6���p����ڑ�@�S@Mඔe����b���A����A���ݾ���6���3f
�kC����S��uQ�׈dعqR�5XK���<�B�����cƢI{�� �6�=J���B��G݆�Z�e+��z#<}��N���|��##|wtB�<9��.�'�������KWx�I�D]\��x6oB���}8o���x�Bg�U-�=F�cEo�����I�H���.�//8hn��0�Ù�RM��-�l�rI@QN<�&�/L�޽ӊ�����z�	�
�O�ѮL��Q���J�~#RfG�P9�h�A�&�qJFq]����b�X��攥P�~p��U$-j)4��3��9�i�ʕ��'Z3�&����L�g�Y�̎c3�#	�X	 ��^ug���ӄo3��g���;�����7Xq��ښ���_՚g�C�5���F>�R�C��G=j+î�3B|�n���
>�q �,M� �9a������H��!IZ�1��6e=�y1wC}�̥���@�j>�)��ƿ��$U�����P���?j��)�OR�>�߁>,,�YJ��f������g��-��26�Go�����Q�g�/�·�q;w�į�a��F$��|h���)?6  �vֶjs��-Ŧ�
mT�:-t[ܷH>؄c >/�׭���@9�y�۔j��g�J�ʌՂ\���T7��z\6��ԟ�z�Д]ꉀ��Ř�c�\Z�"��_I�l!Tȧ�NiY:��}�h�\���^�Ih��'�s�~z]��_�¤��e=�)�(�x���E �SFz�9�V�HD��n�֓6~iCi�օӌJ�Ԥ
7���]~�eA^"�����p�8p��-��%?Q�L���`�\��42�Jo=�1V�+�Ɉ̏��b������r�۰{4�dJ��no�3�]��(
[3���ǢoU��8ǫ�4I:=�Ϧ|�S��@�u�"����LL�����Ă��$��_FHX�s��Di�=���,���Ә��i�o��%/�BT��O	c�ь�Z'UU�	t��Sk���q�m,t�zH���%��i���P��<��C���9��~�hN��Z���D����dQ���+'\��s���Nj�h7�~å�O��#@�����7��"鐕� 1�ئ�JAޙD�C��	��GѺ�P�&��긔���ԏ�S8�x�`sL�Lr�Q}��d]���<�%wP�3:�CĒ3F�z"��s��z�R�nüm�::P�s���K��q���=;W�۔�,��ڠ#C���!L4�l!-��!�v+-@3#�!�.i꾪�C󱩡�Fn�}��;��^��P*u����?�TE�K�a�b7vT�]�(�p>In����ķp�&���,����P0�)��p0��������u���R	ä%d�7��OZ�}\�IU�?2� ��>j�xYzm��fT�u�I���W�Ź�񀹬��Saf?�oq�K�S��R����l�]�H�&��\�[`��p�������[�Jݰ�0��(x8��D:�>iH�y�^uJ!���G�J�\a��vf��eʊ��z��i��C�
�Qo��Bɜ�v<H��Kq�X�����du����᮰jB�Z��Ku�/���@/�X��Y���L$r���In��FgV��O����@cΠ�'���	Î�d6`�����^B�?��\�{F��#�مr������&E�&�	&lU�֮�?�Z"��Uq���4��5i�O0�U�]W��NmQ��ĥ,m�5c�̼�߆�"��Oޒ�}3��4�o�v	�
1.�'ڙ�T�\8�~Y���� ?�\���_�Ʌ)Z����&��?���@��e<�U\o4/�D���ל�6���t�a��SW�Q+�J�R���a�xb�d]ʒ�B<��M��k�G��v��G��rMl��faWw��3gf㸠�����I���j\�&5�������é
#"=`/�ov�YqU��j���1 '@"�+^�s���|�6)ZZ 0����(��GV	�ImR�<�%ݰ�gK@�Trr���S�떬u��z��QF�؈�tO�3Ǐld�n��Aʯ&ri a%��H�&T��IHA׃`N���f��\8��?8��-(-z��2�J6n��cMlFwd֋ke�I��{1��}-Y��<w�X��L������6[���4PZ�6�.QF`��K#k�z(�(�h����"^��)�8�Q�wDV��8�@����Ӱ������-�hey�k@������f��	����L���GHWp�0��c���Y���׍(m!v��p�l��E�~lf���1�G�	��
64�nw!��#���`������t���,�3̚I��r��Q(B���R�$��KA�FB�c!m��p�Cw�AC�|�#[�\O�+r�]K��	�ë׀��p�A:�j0�0�=-��ج�k7�KFo��O��`+	�&k^��2I
�^��jv��o�E
F���[�F���=}�+a�5-�X��@����̎q���>���D�w�2����B�A-%��cl+F{��]���~,�p+��h��{C�Ҷ�b()ubNՃrq�H�_�L�z4�]ǀa/�����S利�.�'ϟ8�J6:�ᖆϴ��8IL��e�<�l�(Rn�u�Th�B�DV���W2�N�k]*���Kvy��jI��Ր�}nA���r7�)",�k�
�6�A@º���h�Z[N{��@dM>����s6�(�~@lML�C"j��<��/�u�͒�f��Wd����RDC��Ĕ7��Son�ېMl��F �M)�f����������qGē
��<�k�z�M�і���
�Y��3���_K9�����Pܳ^��Dm��op�ʠ%!�H�o���WJ	���B���|��J�>,H0�-%�tjEW�\���x�Bn��Hk�����k���ňXŇ��}J���%~���FK��J7џ!�#o�[��:���L�'[�@�c����s��ૃ�~�ĩ`�̫��l�C�Z��:�'~�o������[lEv܍TyO�ͼ������.�x���Zs��S��D�F%���)� >�,�h�z���k��S�� C7`\R�#��o�`�2�h���c�S
҆2�1)"�s#f!�PC6�m�+��?T�u�O���B��c4�Q����MB�A�\�s/�b��Y��"Y9�����͒��j�=XD��J���H|C-
�Cqʅ�#)d���ޅt�[����_3
���{|���޼2�)��y�� 
�bӬJ@v���U��|��
��a��b=ߓ����`��ۤs�SN�������Z�	����zs?��F���8���ɕS��a��ô�m*��N�@����c2��6���%�����~co���J��]X�Y`Lԩ�M�h��B��;�d>U2L�e�Q�f����w��J
��`̺�[ �^�d$��:�t��́xwG˃ʫ_�
��^�S�Iʮ�-�5�8�l�-�GA��Ł�� �O�~��e�1�?Rp?p{�2�y㽱�Λ�LB�Y(͌�i�S$�!/ٶ��e���Z�Rq�A��	�Kt�b6GBP�S�.��v?����mjB_���bz���+u���]���J����S�+� %�E=P��u�4�zM�*
.C��ŶN6���d�-2r��H�}�nG�!�{�GJ�@�����ih���39�1/ "s}�(#CI�6����(X�
@7M�f�2nb�B5'HI��e�\#7�.��g�O��ʯ����P���Uҁ*�Y�w�����&�	�=��h����8i��#�����L ��_t 9F�J��g���a�\��wW����I�ҺR��
�]�cYMn�OV�&M�eYn�8
�齜g�
�%}D��q��v��.�M�.�fUp�z�@�&�e�t���L��sĖ�kĪ���٨�b��+�8�Xý�KQ�-�U�ck�K��l��} �>v���a��H0�mX�v"�� a��H'v��@E�gFGY,0|�
�̘
R���a>@��Hۃ`1|��}�����ۛD���X�q� ���!1"��@Mk�m����l�PnE�pE��9 a"��=�n*�	c��P?7���Qr�~�QE��x���Ƽ<Lm#��R	�3�x�>H���ջ�#���Q�5��
�R���k(�>��
���pf����� �����q&E]];��c���P=���K��~ч�� ��|����WS��t����(�'ņ|ܱh�Œ#֖�לx
E\�6>>��9�Gsn�"�t3jc�?F+��bՌ9��e{,q6A�z���3K:@{m(����8i�u��!m
#��!���I%F�ӄ�wY)Y�L0g>)���Ǽ�iwu�ǻ�P@��n��U>9D���9lܱ_+*k�Kc�6�}W��J!R֊*4������B�����z�g�I�]c;�;�H9yAӔ#��2��_c��*J��ф6��,���c6+}?���Ĳ�
��d:n[!ϙ�H���W��͙��qǁ�fF�L+������ż�00�-e��R`�����:�c������u���5�L���Acɺua�������[��$hS=
�h7%VyYG���X��"�"pZіf��n�=�[�Bڊ��GY�=������U{{v^q:�����!�9Wh	���¹e9Ἴ����"�t�r�<��U��N�I�usǑ�H:�]ј�Uk2]v?�{C�����Ȍ��H=C���ۨ��tK�~�v�(�����H%)��6��V�vyDC!zt^oZ-1�;�x���AOo��," ���*�_	<�,c[�7���_�q�t�v�Ș�����I���Q��F ��kP��&V�N�9Hd�6>�Ν@ �vs��syNA�u���֫�H�.R{��4U����b���+Q�j�;sG�?5T^����m�;���WQ�U5�3��y7�%�KG8WؐS�%�"_s�9�r�!Ϣѓ�u����ZXo#6��[�`_oe�l���|СX,k�����ޛ��D#s�	aq}�"D�I�^��A�I�-.w���Y����n�� bL�f��P���`;'�"-?�� XvVĠɽ�<�P�(,�4���ޣ#VW8��k«��H�Aє<̤�=`Q �����9;�֤�>Զ�џ�6?�o7�^��U��5sV���Ǘ��N;�;դ3d�v��7{���<R3K���My�@�Y����-���[����5핽d:>��O�6-?��uoRE���y,~��8�c�7�ҟa+tQ�Y��y��WF�CEZ�����b�4
�{v��|��pjlP^���B���3�ex�/��.��jT3S� 6<��=鑠�G��/{�G@���`�xF�6-dJ͕�e%����jT��Sk��R����������fW�")��+�q��Q?Op���tg_��.@o6x�"�sxW%q�i]<z;||M�j㝎�A���YY-�׵R�����KB"�q� �Y������+������X�}�D��3_�{}=���Ŕvִ>|`=B�9��vE�k�n�g�Q'D&`���E�\�S��Ёu(�M2��j1���W`<K�3$�tT����T��8^��$׹�a�Q���ȫ���w=@aP��o!�ge�@m����7�þ�h]N�k���_y�T$s
J�j�g�mJ�#d�?P�wɿz�V�ͭ�-��H�Fl��l�D4kkdtu���k�S��nx6��T��pq+��?����+?� j	��wD�u�gR��u��7=G�נ��s�6+�}�c3&&��_Q���j,�O&�H��O�NR��{7Go'���ļM8\X�+�x���s,`�zo�F��e���p�ƨ8�0��3o3ī�C=Ĭ�Vˢ��Q��7�>S�b�B9G�O������ZÇrp�@��tۦO"f^��J���?.nDm�d.��Q�s���q�%���&Cn�Zf������|+32�x��oe4�p�i\໇钙�!�S�Q���)+&:�fyO��p�D»s��-�&�T{@��f=�3BR�<��2#W��J[z�T=z��Boc�ԡ��.�%�g9�3�̟L�K��O�5ď����C�|D�G2�D���DO
^�$�d6C��8��,��:��Uha��R��H�/U2e
�c\+Z7Ō�X��`�g,h�Tu�H��$Rnq�+cZ?~`���ۧ$��ŜZ'�}'����v~��x�\��%��w�nA������. �s����-l ��/���f<C�>(@����$v�@�(�5\T�;5������׹��`N�7I6� �	�E���I�]UE�J��:`���� �I�2���~�^�C�U��Oa���Lҥ��4�u��8���]qV��`}���1\h�UTLM�w�o5���D�5����KM��.��� ��s<��e��=y��5E���t��'����V7_ʩT�/�v�PZ+Th�ݷ�a�.�r^4�H��O7[�>Q,����KGM����lK
q��&]���)��s����������,`�R�)�|a$�G����-�ohte����c�O1�қ�RZB�R��9�?���������S���Z@�Y�+�&ɹ�q���#?������~=�p���y�߽KI�B�k`��������\B�gn�q��^�����?s�ӊ{�˷��H*��C�h� �;����{�,l_��,�F�����H0���U�q}�s-Z+�:yL�W��t���9��Qq&vNT��m_��3j|e����çN�f#Y�%�Rɫ�lW=��}ISh��W�<�W2R���!��s���;� g��LG.�ؒ��ڴ����gY(�u�I��WE���XH��L{�P�ߕH#�:��[ܪ����JTJy�|�8�T�c����'�^���$M���V@`�������ޖvzF����;4�I�;*V� �p����[�?���c�=֨n�}��]wC�o�d�乪k���,��k����r�VK(n�0���-��<��z�{�2�H?���	co"�ґ�M�6��C���d榻�G//�k�yI�M�){�,��{��z]��M#�<2��fk^��D���m�GV�hE��I�1���=����)#��l�� ��:�2��fP�ʧ��] ��A��l0�/�4�%�8�N,����b[�j�}�mL�QΙ�����_����T�i�zKw���nU�#�In��H�ҫ�Fd��ݗ�& �	��;*"����_�����eL]�Q.��U�$��Ȇp'(���CqHh�b'{ij�}�}�:B����u��_�$�Dd*MME[�N�|�Iq楆��b7x�~1�z�V� ;�_���ذ5t�ie3��S�/,9��/j�kI����v_�뾪���)C��xԵk���$:���%A�w���Ӫ�D���Up� e����}�ɉ��#g������5Lg���aiQ�	��yfma�B�'�m��ç���'�������W?���~P�j�WK�{ueo��w.����9!���"����b�<�Iϱ�r		�����b�eZ������Y��L�T�[����rHV�T�[��t�֓'�.]]GR���6�5�%xiԫ��n��Y��%I��� �oB�òH�N/a�6���V|=SG�6x���)�����uǩ$G��{Xi�0�_�k�����*O��_�:�r1��B/�,{p�v��F\u����%߫=.Fv.ɡ<d"�dv"'#��(�_�U6���h�G�
D.�Zu�Z���=R���ҭ�
+��1Wu7�)Hܨ)4���f���g��7# s��s��z���&Lt[�T�R�&������`RD��,�Ɉ�u.tu��= C��
+�y���'�����s�V��\�,Ҷ@� �c�kw�e����t���Q��q�r��f�}8'�9q@Q���3ݬ��֕+���	�)�����v\�(?^r�}���,v�vw��]�3�p](k�ϳ~���2V��������a`�h�^���4�pǷl��<������]�}aς1`:�u0>�w��hp*R��%z��G�'���:W�Z�|�C����IC������Cx�Uќ��tS	�l( �Ж2Y���6��JL]�����;&�%�NS�I�3+%r�'�m��j��ZͷL��s5���yڎCD�r<���}���Nx�<`��0�n.J7��Ev8*/�]|^F-�U���Í�&x֮шQ\4�}�mԂ�U��Ԋ�Ǚ�J#��GkC�\�rLgb���c��w�R_<x��̖��Ǝ(����c��36��X��>�
�9���}|�^��Dy�����{�2���,K�6lK����>�M_65yҥ-Y�l݅-����,���&ٿY��\�J��&�������ݔo��a��q��bͿ]�+;�AE���!���M[�s�f�`����|ZX(��b��s�ma�T�Pq*�V,�b�'�o�9��j�8��%Y.p;���;_�W��ކ��{�Ak�?ϕ"N�J�ΤI���%����U�T2z�Lo����'j����뱡33�R<S�2C'#�\ǆ�7������č ��cs�#�ng��B��%��ǵ��G��7�������Y���{&	7����x��p�R1�!ժ#0t��e��1y]��^�H�dE���߷�%Z�T]��R�nlD��[.�]�?bh�폱���jdRT��Ba�U��6��&��	]������F�{Qw�
�ma�aD)���-:��@-���C�0�Z�0�|�b���6a���g�i��U0�b�����}��1Fg�}����2G��In��򡚬Q���,"4��MN(�S��G�?K�b�C�W2� m�p���k�O&�Ϯ���=��	/u����D��t�zCL�ӔjgT����;�*=�f}�E�$�-|!B����W�p7���_�]݉���De�ߐGq{+�}{�D��u�K}���$����C�8�t��	|���I��{��"0+e���p)�+��O���d��܈�������$$6���?��x�#�}�b:��q��\���V��j�4�Yy!
)b@�ī�{`)���w�VA~�����о!���
�z�������<\޲��0�kC�I��R�EVߝ�c�� �ʀ=A��2�b+�J���v�P&_,�	K��;���©�N��t7h�m�VG�A#�2����.j�a�n�iA��'֠t�^Z��_�_�:8�����Pyk�i��q.9o	���ԑ��f;d[�$�w����U/*o���9}f�Y��>��R�
����$-�~�#��ė���s�(��92������j��o�.+�/6�A��Ok�JÛC�HA���tk��ٓ���t����S��L\�6n������쐖6(��
Cj�[RM-�E�W��r��Dc��/���\ĥ�*�����a�>��<��`"{��}j���*�۟k�(K4���-'�jf4��C4@�PI����Ųb-���j�`@O�Ȃ�����з12�H�%�9F:Kˊ�q��9|y��lv�B:(ĴM��
Y!�������[�Z���e�8�5��&���B�N%�ﱋK�TF��ߪrm(���m'�������%��Q:=��]��gJ�M���}e��)��W��8�߃��m�B)AT¸��?{�:� 
L)�v\�A�q�ZK��}}�@��{B�_��#
T��?j�ǎ�f�!��S���^���4��I
���A:A��^��:��'����̏������{W��+И	��h�܍�B�Yl�sT�"�r�l���5���%ue��v�����":�4iN⑨ �Dl�N%���w*�t��~	? }�[.��K��F���/$�wݘ+��&�B$�{;P���.K򾣺��*&S�s{���6Hd��!��e(��Y_�!��+��'8_��h���;�N
=*\��k�\]h/5S�I�(�/�Nskww ��M��R�@3�룟/,2C��M�0�g�J�1�j�\i��J}�N�K=}�t�ħF��r﵅R��� B��"ȟc�'�ە����(�
�I�BR\����)U�Zd���Br�#ޭs�g.�
y2Z�sC�����@���c|�tj���@�mE��N�A�Y����_�8A�����/�B��a)��8�ܥh�+�al�eh��(�kIq��}��UR�"�쮰�����v��D~��
G�Yڲ��
�ex��Y�řw��?�~�X����g7�;�u��I-_�U��8�Es���^�����戃RL�n�ͨY� K�qV�8(�ԅ'��|�;�ڛ���5�mcF��M<�2s��0��IQI!PЪFd��'V��Md�ty�V+���¤��i?��F� )f,�`��l_�$�Ջ���tc`���;`x��%?�䍇v�E�'����zV0����u��%v"e]RlN��7δ�� �d;Tl
�c�s�D�i4�
���A#5;�ۙkVK~�$mq�zVN��O�xy��BRPI��՝
X )°���%�ׅU�Y�#�9|�p�V�G/��ޙ��B�t _��(VR�����(k�# R^�/7�^q��\>񵓔�dG��V��+��д\��*����$N�O6/]d&�Pk�4�������2�e��R��c�0D�� l����jVv���,~`��%O�z�q~��m�ڷ 왛2��ȽS%W0�S�6nJ	Dxbk�|��{3+e�M�����7�e'm�:�-���ce5eu%`X�����L�m�~��=�pj�񇊆 *8�����S�������=U5j�_˵�+k�/�ԫ[4Τ���5w�� ���Vb��ҁ`ק�*�m
CՂ��N�j�#[��qO���H#!�/Df�)��Ů���u�g�T␨6z�zy���@.q�5���Ւ��B��v��)p��M��F��5�� <l���\2��`����b����h��8�>����8=�>cD!^7�5nˢ2�g�iS�N��
R��~��8txK����`:11]��
��S 4��m=@N�d�d�<�*$�17U�:��6s��l*䢤��f��`��Csuha:t��b�1^���2IK���k/��]-��Lͧ�h�Q�ث�_��~:{��#4����w2[q643�Q�~og��@��)Ek�
?a��G�3��`=9�C�*�������#��������*M�{���� �����B ���@!";�����/�k&��?2�S�*�E��*�u��`Cu_|��z�kb��łs��p	�������Y>=_q����dڠ�i�Z�������V9�pQ��be�fS�@����=�;!�>��k�-�\��i ֔B}G��1V:�x��!�g�j�	j���ef�����4\����u�(j���+=y�.�o�;�{���^"/'y�Fd�bL��U�>gQ�p5';�j�ӟ���.����"v'i��d �(V#�����N~����l���oS2ݲƜҲ��S*�ڴ��ĜruVb�¥�8�@�@R� �n�?tJ~�eyE��W��?.�����&s�W����.����سT ���#,�ͬ��Z0�gpd9�%���� p{��i���2�J+[�� )��}v��.\����2�O��a��ҵ\��4\�ƌ��g������m�/�߸h�ʃ>wSI�$�Ք��_�]�v��������\T�(��3���o|��1{�*�}۸T] �}�JG6tܝ������k�?HC�+|��}��
J���h�EP&�!*�-��zu���{aH��ź�D�ѶVk�I��]fʟY�C8,�[;!�ܶL0C�P���x[�A���1��L�U|����V!z=��M��!O��떑2(��^�d__�I��������\���k��|�ѥ\�9���@Xh3���m�#�뗴F��#�@�W5V����
!T���~�4Sb��x7苖Nu����ܼeb-'�����]�2v;�(�R�1u#N5���ikeʩ{1��0\2�į���"�˜����.Ȕ�� ����i�o�a�"�U]��f���bߙV�b&�o�x��ڡ��2o�R����os�K���@]��4J�:!��JJY҅x%iW�X���f���)\�1��7��j���۲e$�SpkU�`�� ԑ�2,{�}�G�j�=�/��
t��hC1�**j0������������ث�>�_���I�XcO�Kf��U��q#l&
qӕ6ـ�\�np�����/�B����h*A�{,D��=X��f���^��.���!��O�������z��}=�n[O���ش5[�k���A���Ox�.l�^�F��\���R8C�+Z��2u��R�t��P{�c����xvN:�
�m��C*ry�@DF7-,��&������LO};��>�_�����zW����")lFP�<
��1���W�l@�{�k$�o4!ię���0ߞD�k�� Z���T�E4��ENUU�o�x�u~��a�5�Df�6nbAi�W��i�J.e��F;[���2z��	/����&��]Z� ��䰇>�~�A6t��dҨ�,��So�mN�K0��v�����ݧ�Y�#�<h�u�k	��J��Z�!�5�M\i�M�"n��P	��=�Lj�%Ǆ��Kdù�}y��~��$M*<ڱ.шl��4�pO|#c��)��1�<�@8��Gz��2��e8�s�c�E�vҔ��?�{*��zˋa�9y=Z9�k[��`�C��\d�7ڊyThB��0M�ꏄI��u�3��M�f#���i��ae��w��s8�U7�$�5e��&�g��e�z�S������]��)fjQ�@W���h��K�����4��8J�dS���/C��zxL-�x�%﹮�73�Ӏ��h�@�$�ĥ�/m�3J�e��x|��|��O�⻔`y�LL�٩B�4
������� ~;=�fJ'f�&!>�r@�iZ���v�&�E:���-�L�V��^�H�1-A��U�-3+t��b��z�a:<c�*�̰��|A2���~�<_�+�Pa�ȽiS��o�j_L����݈��nر.��zE\�^ v��?�j�ǽ��]
��M8�d�*�G����_�C�un��&a��� R�)
�$X���.'�a��N�ޟ��%�֤��;����f��Ǝ��7tb�z�D�إg!:%��.��v�a)�6�y�R@&`���4[�!T�4����r+���|7�$��-͢�i�{�~]��z{�&���8��(�׊�#!�I��u�Le�)'<��D���oN�E\�{�rZ����`�-v�����!Z m6���;�ʕ�w��տ���Ͻ�Jxl�J8�bw7�_�%gFV1#C�_�����:��tnFIJt���\W��,�-��W�6&��oEDԻk��9���^UD`������;���81�솙��-��ģy!��g�e"��]l�:B�<=X�n��y$����l�F�����'���Yg�h{�T�j�nH�~���o�.dyÒ}��j֮���c�ȦNU�@ە��-�p ��O_4&�C��0	�z�jHpՀF�Ɇ
���!D���&I���=u��Fʼ}f~�Dc�����V:v"{���U�&*�{��wl��� �2oMs���
��:4��;FulB��NL赕4c'z�
��O�{���|22p����*���U0��o8*O��q ���d�wDWy�s-��:m�n�H<iN�v7oJ)��ż����vR�J)�����[���v0��[�Z�n����u�ʢ�K���*�
��ڲ� ��c�ڢ�"T�֪۽���w�QHA`G�.|�c��1}�RLU�շ蠄0R��W�t_���+(� ��^��. V���C5�a�"^o���KJ>A��)�Y�י�x�������1�,�/��fFu�T�]���SO��Ľ!�H�ǏӪr�k*��vc�QCɞ�b�+d�'P�ag����t�����s�1p]�����4�f�*���g�z�/M`��/�֓ .�=�T\�������-�8S'�R�ᘧYz�n���qV�K�f�(aGBfY��;yhm{̪>Sd��b}}_h:�C�0b�*{��>�2���ט�E���
Wcg���trƋO�}6{${�7m����Y=ߧ�e�����c,���뺫Y���F_ƛ��n�Z�ͧp�S��x"MF��bVF������y�b��H;uu R,r����Ԕ(�
���	=�"�{�3����A����c�z~�[� �������wp�r�_
���<��M�+�����@:<x��`�ӵ1���(�Ӆ����t��lG<����A��4��6K_�X����1T5��P�	f�� t���*���%�E,s�VV��8s<E��4�3��E,�e����m��s+=�[�����C_0�?���檉�;���]���Y2��D?�-;c��q�~%Ɠ�O�+�,���DN>�y��:$� �71���F/�@e7xKx��q%ߊCX	�f۠:�:�.����6 եU���A}Z��N*���Ѽ+�A��o;SMz  ��$�G��yȴ#�����xdqH�U��k�C�@lZ˓�b����U�f���݋�M�]QSA��`tb82R.��++��(C��
!\�j齨T����IYzL��0��/M����R��7���V���5=k㹆��`�,�yB���#������~ZQV�2���Ah�)�a
�-�����o�6�>~�y���-ȃ�D's��2_�1T�@���ү?��޵f�(��!~2�E
���Pr�&��"�^¥�&o���y��|�*
\fG\z�v�}����AW�=��=�N�D?���2
��b} du玨Y�=�"T��r�?b��8S�̸T��{�+���:�Rn*������œ`ϥ^;�z:e���@��!�ohU��?g���/��yr��pO��h��E������-pB�n���Y
E�Z1A<:P���5��Q��"?�`A`�aL�t�D�)�Y��*���x7�J�W�j�b�U�B�)���	�њ���9��;뢐���?�lL;3�خ8
)-�&j��XU,�tCZ��I	�$6�C�暛gM]�#��]n��&jW�c�?9���W]��Z�7�&8��k�d�k@�Fs�B�@
�p�`o����GUa3avNw�ζ��>1 ��z�o�b�t'��3B;�wJ�����K,Jk7�(2��o�a���u�V�-����z��zVۛ"�����>҈�S��r�__�9}�@<�j�iB��G)A������x�%dT�D���>�8s1[$!��L����ŚR�����B'�º����snj�bt<$-�;Y�zb܋����:�����������j;B�F�ǌf��V�L��t�@iHG-:�Z�=A�GX!/���H�ə|��1��hg��~Gi�C�\ۂ�@��wBC�{��X=,����I�I&����u%�M%@�"�(�$ׇ7���sW�o��'b^}͊��������e��5�W{�U�w	M��Օ����{�Ur��d1;.�1_:<]�噀$����m��.���u"�ř���V�oQ�M����<����@�G�|�Yr�V����L	3��ze�]ᣘ�L�)� �5��"�uU���E��g��\W�Z~c
��8��T)}o��^a��5�z@�Ofأ�e�˶[]��|�]�h�$����e�g�?:����6�w�|0������i�ׄA}���N(��>��P���]VJ�F�'û�
���0T���g��k���S�a���}�p��*�>=t��C��R�t0Y'.wD�,��o_s������&����Fϖ��Xk���[Yq&,�������k�p\h�0� A��kw^�Cb���-�[.���]�u�E�xU��?��&�L����ntK�V�K�_�4��H5��~�N��7 ���ܙ�F�A�:a/Ł�i��]��� vcə�HÓwY�G��;#�K8��Kz0TU�6��Q����Fp�<z��"���<?��(v��A�M�?���G-W%�er� �w2q��z�qs3��Qi��sER�["ض��T�_*�[���q��<��ֆ��-���؄nX }��x�u�[���~NņC;z�iJvL�����Ž� ���{m��m0��M0�v�9�VnZ]��q�4���ϱ����~M�p1WWGvV�R�	�2y����}Mf<h�3�O"6;ɘ�\ �����=�����Y`�4ʔ�ܧ������\�,t����U�)U� ������D�(��k�澊����_�O��].mFg�� J��T�<�j�>���`eJ�z�j�.�P��35�A��Y�pv�x{�Zv(� ���2���2��l\H���_�F=�N V
�~;e�v�N���Zx_�@��\�>V�0X�;�"	���G��R� +%�KG���4��s,Ig	��_�
/��[�w����S"R	������[X�Mt�����|�:��k��*�}0| ��aA��	%��1�@�,������ܿ/4<j��H��>%�?�Lp��y�;Z��A`�G�4[&��y�S��I1�*}{���p�Hu���w��!:1ѫ����� ��p��	�u�r�P�I �-�ʙW�(F�^�|��U�����`M�GK�uv��_��g���9�;n?rⸯ&�p�P� �V����3� �Mw"�m���I��#`����L�C�#}�K5|���w��9/�Y��E�wOA��4	'ɗ��!{����:	�;�g! ��j�"�{�`i�	���z�q�+_��<����ݸ"�o ����Q��	B�q��4�*�SF�JKj蜨�vd���S����V��I{��&�Z�!��x^T��-ցN$3�˸���N�F� ���S�\&�[G�r����T��&S�ظ2�/s��j@�^��c��clD,%ף��7_�	��-o�R
h��A<Dr��0���>�Ԣ���m/|^_���p�_╷��{��	d����蕨_��H���� �؍?�,h���E�@[���;R����/�v�!��Cz��.I.k�FA&���3q��@/�Ӡ�lZ�Y��zI�L���K��ݶC���+�пř��4�� �[���4���,e[� �(� ��=�E�t�.��^*�����nR	a|O�Q�"6�a�6
��{��aQFb/�N��\J�j�W���5U�dX�%�!�V��[��S����SM�?w���e\�˚�=@��-pḬe�t.^F��V]v4H����J#^i�Q�T�a�j�Y��l�3>����?8��q�Q)����L<C���y�cP�C����?�����t+�`2�I�^����F�Xs����6bK���1�j�˨�#��?~mX3W���L�З<�P��}�.M��U��� ŕB$�F��Ώ]���]��p1^x[�2�c�
Q6��� ����0�{ �6D"k���(��V.��Ӥr�ߋ'�(S���x����ς+KUmB�e��%Z5����L�@����y������[�%�<��d.P S*bŐ��(+���b��R�R�&��C�yK-���7�v�����,�1P�h����+��G�Fi?���t�U�xې}8�p,��`�
��H^�Ndp��g�Cv��Y�{4�����di����<��[�#�G�:s���I&LHƿ:�<���yh�#�a�eY���]�	/��'-��qG�ze��rĿa�b����6A����VN(^�J3(�����{���Cy��L�<���։��n�)>��=:r؈Wn�=���y��?���1��E�-'���X0`��t����yd|{���ofwU������|�-��+zRmw�\��U'�ܿ��@\�|���:I$��C(��:�ŢA�<����nT��E%�Vr�nj�3 ���Q�؋�3たs�_�6���O�U�R���|�l�ο�]G���@�#s�vo����+B>*������
���j�=�t��V�)��� գ�W��AN��K�#����Z1ɺ����n's��E�L^8P8�%[JYV����=�^�������t7�P�e7��>�wS���&F+�I�B㨑�nK�c�J���{������8��G�.�`�S��gEU�z0��ה�u$Ng��Jͮ&�~.q:����Ӓ�`�Ss����dw��-	<�OW�4��&ur�Ǖv��5�j��t�Ē8!���*�i� �?�kWI��j0�W6� q�ěY?�� �<hh�/��;b���� �*?��$A�����t�� %趷Z��n�hxzjw��+���[)��@��4ߴ��{�����1<'�~Na��((�&H&�"Ky6Lo��5�sy��0b�E4��S���)�<����[	^ߝk-�j��	���ن�n�Ƥe��C�+��NV��ۉ1��*�u�v����Ť��u�i1���'ޠ�'ѭ�╀���n�\���"��⽻IB=4+m>燣Zyb�/�Iq�+?2yK��u�1z�F�胺Vk͑bh�n���^:q2q?� ��eB�t��E���+(��he�)�<K�Us5[��,= ';F��o������ȏ��E6�,nt�O�&�Y���'�8���'a�:AX+�
սU	��n�Y�cek����	t=�i�c4�+Eח9���`d�Ҳ��O�j���Yi�R�,2B��f׳p�}�t(7�R�ƀ;mw�T�1ɍD��ԄF[4n��7��hV��6+>�Y�+��(u��IbV�v�ɧ.�?�]j��-H{`����}f�01��y3E������pT���Ji�u�]M�zl�����9��L:y)^�/S)6�W�G�{���$�%�?��Q?����Ӣ]W�2��`�[���7Z�q�)O+���Cu2�X貕�� (�7����A�Q3�l��j�vi�_�S{GhW��( y���d��P�[}3�D����氕t���Ӹ ��si4HHg3��X)�l�zɥ05�å��;�d���SamV*�?B1>E��_Gr�z�hM�N���/���7L�����C���>�O-����,ӄ��%�%��Y�Sy��,���uO��d$��=oř����މFّgt����N�
�w��_X2̵�*��Գ�M���H�b�����{�)��qd�t\��]/��r�����Zc���E=�3G_�����Ь��W�����FKx��iJf~��[���7���Ij�7�O����?���1��+/2+���%B0�4~�9DJJ�s������ח��U����$�3d��a͒iE� emL5Q�/�f$�{�_�Y���?��Tk���	�4� ���;�F�2B�(8e#:C�+��?�ak�ʩ{�/�LOFo��!^�x�]�,��X���J3˪X5hD�7���LP;���^�h*�{���[_jmqE8;�P���_���ZwF[
%���yy��.���9U�hZ"ɷ�}q��"���ؿ��­f����X�[���-)O#m�e��O�<��},�i@Jj������ l?oy��o��h���z���9����!nm� g"L�!���N%��y�a �F��I�E���ґ|$��Zҙ$];�����,,�i����:_�d�$��Dτ�]FY�^�٢6�kB�i*pa-� -A�ܥ�7�d��P�T<v�p�'���$T��
w-f�}3;«��o|Ec�h(XXDC(s�\�}� *Ez����% M���I�o���\?3��V���R�
��~H�Y�ڡgٷ�Yu�d�8,H�����'�j����G�ǲ��g����%Ƽ ����-��5T�-�x\��#t�� �3y����h&s���?	�E�F�<w�|Ӱ��z�~ܤvJ}����6zEU�_:���>?S�
-!�9Y܏��^w�u�M������a�Ί�8,�0Vћu�>���-�aLU�cp�����u��	�=�
�b��'�B�孿��È|t�'���H��`�ѓ+����uԂ�5�gI�E��݃}�!�StΫqŵ'�G�(��E��˚� J�U�k�q�|��C��+����c`�u�Y&QFd0e" ��q󚈀�~I*�^����������m����>��3x�-,,5h���ˠf�2N�j��Ȗ��]J���G��M��V��Rk�-,j��)�"���/�"��F>D\]B��F�e�G\����0#)�����$|��H)��%4�jBM+�M����{���V����vE�F�ol^u0���s���V�O���5t����nb�]ߑg*�Ǚr9�\+��ϗQdд���HA��AR��2���~��R;�AY�pp�	��T������=�v�ۍ��߳�0�/�;��G3y�c�͈���v���BO�ZC�Geve�y��ˋKT��x���������w�(Y����
p�����m�a��Hπ!տ���y��gt]mc�M�-�xk�"��/�~��|V�7���<E�G����f��Dtk��8>Y3���A~�� '�"��}h��j�Z��o1S5���x*� �����������{0�]h���S��P`hK"R�YM�
+����Ү��Es{U�k�
��X���ZZ<k�j�yUVm��q�Sy��0N� �+�`�m��¦A'����W�;�C�@��F;^7��Ή�w3.���B�q�	:zTSt��<hC��*��ɶ`%>��XeW^z�j�wӀ�%X��/ ¬��(T� �;�L��)�` �222�����������.�]��0e�be�e\Fʪ9��ⴟPq$�c=�����(|w5�{�L�G����:�!��s��I�d&��#�-��.p��MAGo}�>�׽:�ƌ�o	�ݾ���#c�!⺯^=�md�W���
eN�ѧ@��Qx�	1(���)��9�+�hF,��/id�����xqq[�� S0OC^���J��<B���5.�`��\��~���3asQVO�=%
/j�*K�x2X�{z�8����-�D����U�	p��9�f��_<�^+�4 �k~�C"�������T�c�("s������Ɋ���4�t���X�ik�a-�'q���S�q��oԹ��"�,B�!nW�Y��x=V��@�\I�2qF!�w@���=(C�!	-��+⹠#!��}�KG�p�����p��CzXV�`��0��V�Vh��-Mh��~?��p���9|��)S���ˍ�շ���1���c�$��t��v�u�$H�yNe��/�h��֘�*���8)o��� �8b�d��d�ر��w�h�q��]]��d<S��Uj��M6�YqS��#] 9���HʇH���Q���}�y�Y_��&�[��c�f4?��&��s�wBϪK��DY�;���bn�[	w�Ӽ�-���a	� -�������0���J���B[�Uj��I�k���eا�w�;iA��27|$�Fr��A�a���U�0�ݣT�$�Y\�����J� �AR}&QD��I\�|É�d~�qɞ��p Z�p�>k?<:�0���HY`���W���a����>�D�)��w��P��ZY@_�X�i���}Ҥ�Bj,��
��{�?���]��F�#xa���G�	T�%��J���E98�7$fl]=*������fm�t.��`53ϡ������w3��'d�[w!"G}l���Ed���7�6[��L����"��Z�9�����3��!9���e���Q�]���h��
*��ϐЋ�mQ����ϻ���.�.#m��li�=�fb
���'&s�~�.!��xz�N�O�מ"0��.��;��X;�S�p4�V��Ϋ�H�����7ϸm%��
�j୯/�P���b�8TeKJ�<�緶B�����y�����u����,b�SBRO���P��X���ҹ����"`�/�;6�L�!y�wJ���g�e�P<�@�,ij��a�d�	ê;�ZYF��W4�8��:rU�b�1A&`�_d��t�D+ߏ�Ϸ��;��ё�!Sy����_jvp����'k�`�>~=�f���Q��Y��X�8�)(3��}��q�G�H��t�	w�-E&V�Z<a6z��}�>�a�<mS/�>Ƃ�̛֗�����U���g�z|�ꀤ;�����7�z#n��1�[�&��u,�iP��%���:��[X0�޴�Z۬֠�$ǯ����c�T0a)��L�= �0��t[ȩ����u�M�<� �+rXR�x�\���C��ƨ:�˛G���N3��1��g��Į����*d0)cc̤{8�J�� �Pp���B��B��lf�^���`����NA,� ���U�v�*o��;[D��ş%�V�X�cX̴��QIi=�ѫ�BaY���c�Wo�S��Dg�"���:Z6����w�i%$��.j�kE#����wP9�S(ْ��:y����s�:`#.�;�4��O��Swd3Y��U���婝Ώff��r� ��݁�/����M*7/��`��:���n-!�aG�#*d��,0�BY�`_�={�o`E_�MN���ž"x̨��A�@K|x4N.ëG1�f�TLq�,ڨ��7ǉ�O}�Vt�C���s�����}d�+��1b�y���I�s��*zZb�N�ӫ�ʾcc�)���|�j���=�*&�D��<��4)d_��I-t�h���?KIP�_و@O����t|9�AT#��pH���7W���\���ض��TC~����nZ��oI�J�[(�sw�$L)sr�^{���ڦ��4�*��ma���΄]"��L>����Z�M� ����P�(�
�B�#ͭ��h&��ZP5s�V�6�K���#��L���r�q�-�☞b/��f�I,Ŧn���y%b.a6l`'z/n ������:���<b������y�AzU [�u=��</!�Bƚ4����{�e>
2Yγ�YO�q�[֣fڏn���Cw7ː�Cn2Ź���s��)^Q���IP��'8P��C�+�GƦ���=��.�cƗnZ��G���� �I��sR!�W�ֱ��y)e�*j�y�JX�֯���k  �Y�Sp�8$u�}k�OB[�-J�/ D|�D*�:@$S(� �I��w���;����u�m��-Bn !��ƚ�0���M�0z����Pai��׫�9����G\fl�LVλHd�/�Z�r앧KE������&w o��OS
ȵr+�v���pB��ĉS9��E�|W�B��u���g��B������&�ר	�օH������Sc�T��qC��e�_�����W�,N<��G�!8���1<��$bh�_��AY�2�\�f���W��B|���V�g������zM���5oU�,�r΂����ļ�$@X�w<��*��c�M�IuN�_��8�C��t�w-\���|*�n�ݯ��:~�`�mB1�*��Tխ����:{�o����v着u毎*����P!{�:��f�E��baW@>�vT�sJױ�$r5�s����j�����#`����`�o�)ԁ����%=US{K��	���h��#��y�%ΠN4�*���"A���mo��]����D��TY�R?���&$F�[�@\mA���n���� '�zq� v���q�m;�"ǈ��u���C�4�& �(�5l�MV��\��&�ۼΰ��0��v���ų>��8�vI羽@�üX|_~��!4�G��x���&�ះNeJ���k�`�%��&Lq�%�jy��tԹ?��@��0��f���[�R��s"IOx���ΉdyZ�M�w�I�UC�g�~*�d��N4��&ٟ�N�i���B�,?mA�Z���y�G�`sB�zK8k��4�@_�ZHY�`;ظ3d�Gt�Cg�Auy���f�@z5�כ��ho�ۃ%l��d�/ϒ�ft*���){r��k'k�P���mI,��E���7�@�?��o��q:q���m	����H�GMbXA�@���'��PZ�ȸ~�^I8B,8T9_�6e��Wh��maV"��Q8� �`0�(9!m�YE�u}�ܐ�Ŗ�3-U��ٽ��l���j��n�8�IN�SD��
�:/�z�7e�2h�������Y�+߸���*�^������?�ײH��곏��\��f
�vU�c���}��������}z��{�2����|���K�k��L,̱�Nr�����,�����eJZ�&R����^b��ZM� $%!�&A��	|U��FN�B��{��t��r�o��>Lx�f��Պ�s� �#,Lx<��_ӳf��;*�02�Gpu��(�.��~l����JRL�]�t���x\S;#yr�Ķ�Q�ۏ+����X��^�u��)F��,Y)$N8��R�.=�PהI��j��Z�*�s3M� ��f�ۋ8���o��K��}&ck8�|�>*��S�ٿp�d�h	���~��N�����E���Py&ID%}xWr��@ s��K���:@��'JT,x�������K`�PP��6�u���]5��bT
�������&m�.�� �2�^w�P�?M��)M#_õݴ^9%x^���5��c�<���j���o{n����q"��4s&�Y~���Qi�������`$���Nޏ�$���M���A�%����؃[VpZJ�>���1Z����?t�A��|Q�i��=vz��@�����OZN��_zCl�aR�5ز�sa�u�� Z"[��I��Jǰ=>����9�ʬ#����Y̯��(/l$KXJ|k�b�ш6��t�¶B:��d�myL��0�-K_S��x��D����>!� ��� ����\8zSVb�ܣ�gzq!�G���8s����^�l%`D��yV"�*c�T=��E�9�О�m̥QN�O�?��*@��j{&*���;N�8j]��E�=1�6D|W �
=�Wz�\@"�t&���g����,�8�s�?_zY�<��*-����>�P�2��1�F/]�@�x=u��/�L�m���=����V��b��Y����X�5w���\
��8 ����򻪧���b�	_-b*-癱�Wk�*RP�A��6�Y�x�2��~��!�6'�=��-��f'-�ya��^��c�[�oٻ�����
tpМ��w5��c�Y���2KT+���i3s�}��{��a�86��n�����J���X�ڴi�*�Q�ΐzS&�'�����G7^T6%8�m��Z[���� rV5ϣs8_;���_�f
<�øgc{�~����� P��h\A������T^r�6a�*�D4FR@+�g�Z�1��e�WZ�%�o�۴d,�OxB_r��/:;u1J�%�����ħ�O��@^0ú֦��z:x3��u&��/T a'�������K�	���?Up���#�rL��0W|��
Ǯ*S����
�C�X4��o潉�ɛQ����ծхŝ�t����7�4cpi�'���pr�A3�]���Ѧ��r�hY���^L�0��C�a{��P�Pn��F<VMhBT)��`����G+�)�6l���]L/�_�3��5�w��DYa+Ҥ���/_J;��-�;��Ʀ��=9�ZX��T� �yn܃�N�m)��-���(̪�1Q	j6״�%��7d��ܘ&$U���Ի���'!���*�#E���S���9��P��
Z��g~���w����\�����.�Φ�j����;�Z(n}t+w]Y�/�#�X�j�$k�0v.y�՚5&�@��h���Y���I=�����Bw2UM�U�"��8<{V�1LqvU�)L �,�.����ܥ=y�`)��Û��3��CV�=���[�_P�
���i:� ��6 �H��t�7M�:~���0Ci�noD�͢���r��d��;=,z0#0����T���	�S��O�3\ܳ_5Ov��`�Z-5� �L�n^��"�/�/v/;~��A���҂�2_�cWg&04�c�`���頜W9u5,OU�.X�gS�����D!��. �&�~CsPx��	�i�F=&���=l~�G%7Bl9���S��ë�|����VS��h�*x{�"�T�Ĕ����W�*�r^O���w����(������J���v���Ԟ�Z� 7[m
&� ���ˠ�1�-\�o@�3/�ٱ&��|���/vvѨ�����x���=�����`��Ć�[�7�� 27Λ���zI�~�T�mg�A�Zk[�Ϝn��"/4(�����~�B�j�{�r?�'��w�I�-а����Is[0F��D�t1�D�o�z苙TqZ,Q�`az�|�q�r	��`,$U�T�Zu�l#��;$��a��=�F���"�_n�1��T�a��<m��(����gZ���&Z�d\s'�Z�D�_�����<��9q�TSD'Ձ�&��_ v�\{$8[I8q�qo�w���NCU��ua�0��x�ؒ=�(MKM�,W'�wqd�9�� �F�em1���>��הm��Sa��p֑��!�z���~q�L^ɷ(u
-�����d����6L[�g@/�F�{#)�ڮ�&��U��!��.1�>�#|%/'��>cҬ-�&}
��f�ĦS�h����$pޏK��L���Sѵ�"Hx1��p~�K�Y�J�^/A:��[��,�n	!�G�09pK�0(r��E�@�e��d#M����R�n����s�_(Q�X喅߁�
Wd�G.��)�Q����r.�� �t�3��1<�QT�s�y�4�6[i� P����|�L+Z8����^fX�K�����Q�Z̻4��@
�ţ:%nЕ� �y2wv5�z�BЅ}Dھ!yAK���Eu���;�
�6�|�a�R��=���z����SVyn��n�`���CA�́�����F�~8'����,s���0`$D�X���x�1��D?�R���<S������\�rl�T#�+=˳{_����	����(�ތB���ۺ`q�-��,����d��R��ܿ�9Q�]���}h��c�m�ӝ������� ��d���pHc?a^�fJ ��t>[���7W�q�+.~���ua}s~4qEW��U\j�?�2��<)3��O9Rm��6������O"���4�ig�\N�b��e�T�b����q�f�A�<��%�Qζ��D�[3�� ��#AǕn�̬��h��q;�FeB1$�9����K�
dD���xy��s	��+�	4p
��!Ե³I��s����Nz�H
1����=�|�� q�_��������"����K�F� g�_b��~1���:7���̥ g��~,G�1y�������ఱ�6I!Ej�۽�T*pJ�^�r�����чX�~w�ck���p�Y��k!��l�Y������J1�>Dի
 ��8���;׃Gz�Oh#=�������C-�k��=|�|/=���.�T�DZWZ]�@�����\؊�ڨ�?c�Al9%>���ӆ:%�3������j
Op�]k�G\�]'c�]��T���͑�B�w�S5דtH��1�Fy(�(��JC���v)�L�mv���`������i7N߱�����!�L��)ia����٘��Br}:�v�(�r��� �U����8 ����1o� +�}��O��N�,�&�fJf�,��z׼6	=(&��Gx3|�#��޲����i�h��jON�t��B���G�$��S�iȯ @zV��p�=�*΍;R��9��'�b��~�J�a��r�fMS�6�$IxG�琰شڍ��k �7	����[hLn
��x�ʦ��W�/��2�G��s!�����;l�T4�� �9!?�=����ĥW/���o�~	8�vh90ר��Eq
7�$���O�M��Ǉ���������-�L"}ZN�Dۼڏ��oD�ey�����i��O>O�w���dp�� 8�\�O�;��k<Rd��XCn0��	$��X���,&W��c;��B<DTç7X̚�h��CW/;m\G�Rd�s�Chv�a�^Ȼ�O���z��$d�&y[�Vcf�N��_���&t }\uO3at(�N��A��9�`�`l�%�ggj�Y����D�ٻ��*7>�"��Z���7�Rh8E������j �&��B��d��'s�^uAQ�\�y��e���FDl9"u�K ��q��Ig)��WhE�k�R��[�8��u�Wfz�^�R,f�	��u�����M����c��}�,T��%�oA�ꘪ\���b4�f��,	F��w�:!�{�Q��p��C���������qj�֔x�2�l��JN�ԳA��K4z�_���A��VZ���Q���ɳ�5m��rw;}�6�-�DQ���&����������DO��5T��B�;�A�3	�A��]n�k�'����0̰����[_~ԸD����򁢇�kS�1i0zH�`;��#`]�v�"\�D�s��s'��x�����(�!��/�U� ���j�N!�O�wTY|0�?�z%�,k�e;�X�v��2���N�o�����ts4p�y�{�D���#�}F��MIy��QϒgZ�[Pz�L\�!GM��p�S�����LV;��/����(�����Z��dtut��`�������Y�h�{�<�]��>*d�;�B�|��T9}��Pf����s��h5Y�g���7ji�:%�W7�kY�o��]�7l��b퐊gƕ�P��3˙}�X+�|��yd�]���O��Wf%�4\�(����� ���NRds�"tƝ��h`�1"`-�t�~�A�*ȆJ��z��*K5��A�w�R�K��	���������ѩ�5Ei�N�^��E qZJ�U��<D�����:ǩ��xr��3ky�DŬ���@ڞ���n�z{|����]�!u��HZ�;�.�x��Ɏ���Ҷ����둇n8n�(��Vb/6�)��%Y}\N88�����dB;z�{*�h�g��Ai�iPz�,�OM� �����vM��u4}��M��Y�84����τ�	��-�n|�>,�R:�
rAt!�ߤ}��Q�垱3.�KV�AZ�j$X�A��LΑU@ԧ{V��:�-?P��$�^z��C����	y���.��".���S��dέ�rH�a���b���|��	��Ơ����f�S��σ b��n�|�9�ڍ8h���R��s��B�R ��'��lA#��_����\.6��2 �j��@+׾u�m�K(�'��eV"bg�	�}���e!۰�>���T�w3���q��'��%���ŕ�W.&+z���oI�
�I����'��J?(�A3Ga��Ac�XJ���;>
��z�^/#>�J3
���*��Qtd>�Ճ��)���{w#��sj����� Dq�_�..+XJ�Z��!��:s�Z�h���8�)�Pt	��g�a����5ݜ�FD1��<qQ�]Ό���IQQ�p:�B�3;����q��.�m��J��/�L���^�ṕ
�w�o�#�s�إX��� ��1(�	�A��ҫ\z�&��xBZ��<sr&l1Ē�>gŦ���ϗ~�.}{K��>@p��ׯ�Poȿ�<�E��[�6�"gă��&cj ��,��>�NF�Զ��@
���W�.�ڇI��}i��c@ �`cE32�"���[7I�H(0��ɍ?���)��*?R�tRj�v6�eC�%��H[x�_#݌�{�PH���St�8�#�~��y��]�`	i�)c�DZ�c5.�b�=�P���6`�2��֣Fc��#���n��MΏ���/(W�u*�l;��G�w̜�/ϵ���"1i�5Ffc���]���	7�� Z�ő
q����H[��ׅ�E��w&v�����R��(*ʜ�����a��˹~�Y~?f]
�O���溂�hiǴ�nRœ7]|ߥ���\d�����G� 1 v>��@('I�i��,бgX�ƴ�SAp��c�D���3t��&�l]5��>7�,M��󗶂�ԗeQ9_b:I�In::�^E5�U_W#%wJ�8��p�Dq!̤ʿ����et\"���o�4� #�?�e���u�����z˽��byq�|�|�b�qG�'�ҳ���'ެN4�&�xw�������QK>�F����Ziֿ��L6=�n�V�v�%h
�>��\�,~������;�'pP\��&a����1�_�k ߐQ��.�~W|kw��_�_,�~�Md�j.��GR]�z�JS�	�.O�k��1>W���㟝V��������<��B��-(G`B�_�`'�V���|y���� ��:�*Q�d8�V��J���,�4u�"�.�u_�>i�S�Zy�&SR8��� bP	=�y6"�)(�A�}A֣�����fm��{Ŕ�R�o}<��$>o�M��������BDw��^[�x����E	�#9}���!�1� ����Q��y���nw���o�N�WHvd�s�Ҫs�(-����6����L�(]��I[��d��-����#H{��j5��$���!3~�㴍L:��M��UT(p�W(�\(j�X6��D����aR��m���%�/��{��x5��%�UO�Q^⼏�e��Ф�g���9E�MO���HE���f���iz����-�h���X����%�G��Q����S�g�)�_.�=�oò�NgU��uː�#S�K�W��Zz]�S�Lv��R���"�qg�}�kLӕ��[�
��d1H�C�f����fg�
@������2����.��}��rȏ��'�W�t4�+�2�0����g`�����<��/,���e�i	$m���B5�扩�RB��&[�ѣ�Y �5O42��2��9,����{��7��wzLf;&˟�JGre��ހl)�=�����%�������EeU8*mr����-Te�&$-͖����/ʛ��M�%��0�[���բ��3a�rj/Qߎ��x$��c;���gk=V�%t��A��hQ�L��W�����'���BO��՞�I�T�I��j����^d;K�j�f��˵�֩UR
a��פ�����\M�Ns�O:j&$�?Xvh9���ao��}�9�[p7Nኒl쉯u1��G���F�����u;2�Y�L�`�TW����iC��혴�<]��'!Y��)�1�@γp��GH�|O����n�1�+�����ס{�b.>�&���Y�ϵ�q��X�Za]r}T���?��&(�c���j�o�݇�㒴��5�ӯ�s��=G��P�t�uV�"Pu��P��u����Wu�}�Kh��vjcob���c������c]j	��8i�}�zC�-��R����6���1�s=�t3s��t�C/�\�%E�R����g�����������	�|�]�����'~S�r4�&mό��Se�S�,\�����l�<���f�kb�Be~�$J?
����}	l|GF){[P)�'y��$V F��o�^�A&�`vy*��3��*$h��m_�QwL�5K��Uv���^$��ߏч�Y]��b��_]���_dM�%':Z�Y����%�8s���VT��b��"5��}T'*��'�(�T	
^��C:���Xc=\M��7�IP��y�t��&�9 �Q�����[:�*җV
�U0L�P�0��'��0����R(��M��g��Nś�w\L�dy��/��&��a�[� U|)y5|-B-0�柛����ټHB{�����Q��H)��p���K/}��p���zV,�H�VB5���ɶ�3���+&�@�g=�u#�VNb���Ű�՘���Q�X�H -��n�zX�bS0+cIj�+,?FH��@��2���=h-;���3�0X�\U��=�C7�t�f틒�U�;hX��w]g_��tʀ�l��p���A}�i���)V��:N8cG�z`#f*�%��p�?�Kd�R��p)�W.��T@����o>	:7������9�i�D�����s����1�.�I]1,�c���8&�m���W��;�c��q�{��,������g5�b�`�(R�����6o��{Ni�>�u��������Ls�Qu��_���sĲ:���jB���`�uC\W��K�ݜ�kx�u�N��)K����p����9�s�R#�_���I�R�7⒱#_�}�Ҿ LFf���2�g�t����%8��jѵ�oHIMD�R��a�&W��5몋j�;L�X� c �^#.�����g��NDa��bܖ
%��V�눛�����B��ܚ3h�Ϗ�-�o���[i�2=�/��q(��N
��a�B���]���*��Vj��s�Y��n}>Hv�8&'� ��YBʀE�F����C9�U��8J���ʮQ�2"���n?�9X��h§q�VL���n\��
-��Kث6���J�w�ТE�+�Y�
g[�c)�\x�B�K�S�nٺÝҵ��]}��KBr��V��E�LpA�j_�u��$D\���;�� L]@�����]�u+��������[�N��$�]�ye�h`���A��������E���d'i���5��tWrԼx\�J���C?����k��{��ˍ�W9�pHs��j�3ʟ��D�C�ً���;�n�����V��+�A�O S��o"|vv�%m���[�VT�i�۱}�~-߉��}�"Խ�^4���u�����u�:dpO��j�;�D؅�p��3��[ц�df=adUhⷄ�	�0�d�]��b�7����Uܭ����w����FSYp�T�Z�Ta	�?���݉����G�J��P��'׉�Cڀۋ��	45�7�=En��P!m�5�D�C벳��P�ڞ�a���r��#�մ�i�`^�`�7��d͟�����r9�GK8<����
>��e�������Q֗�?�W]��2�5����!~�{�^JMȉ�P�ϋ����s=�8H�ZB����J~������ ����ׂX�i��]f�˔��!�'�Ȣ���=���=�9:K21�m��M�G��y>(S�؁�%"q*�E�>����W؍��E�8�� mc���<�e���ZjO�8���o�b�V�����	D�1G��!�&�r7z���f����X��uF�!vuH���?7�v-Iy�W��>��N�A ܭd�6�=���������Ϟȿ6[z����a$�P����ٌi���>�~�ݍ{C"�a����Õ$�)�U�a���� 7Ak���)���(���O8��\O-����[z��ڤ����^ke@,0�78�B=�j�;Z�rI�.ҏa����Y�H� 윛8��s�\��#�}؅�ʬY҂�E �H�B�i|���Qj�r��`��h��߀��1�fv޴]��d��L[�>P��"��/;R����$�f�����V�э1����u4�+��~��;<i|�?%���y|�)c�s���Š_\r5� �7�N�z��{M�޻�BW�'0+L�\ �D�6_�d��x~m������坒�U�XY���<R�Gq怱��)s���
��~�	�$:�S'��a�$��ٵC�����<�0jN�Ь~���#�d��M����5��:�e���N��vyn�x��;�KG;�q�k)I{�S��D�N7 T,��0�pΕ��F��ص;�iOR�b��8b������o@_l�� vxi��V��� [� �jS�G�5�^��X�,P�T[�e�b���w���W��>�Y�o�/h�:e���ՓD����Q�N�� N&�e�&���В�Ƿg�2�'ѫt4�C�����[��xZ����V��;��]וgc�\e�-Tr���I��{K�n[��:߯�~<����n=��PK:��'ծ��`�l����>do��Zy5������]��F��i%$ߦ�k_���H�]�?�by ��ˏ�0$��S�>���D9�Մ�r+&9�ڰY5���Q��a�)��;M��X�-!��GE��Tp����|�Υ�������@�'Z�3���������BJ:[��\k���]E��༬9Y���M���3.�����;gB��S�t�bު�ܷ x@T�6H��-77��b�_����M&~<��n"�mGEB�TI��!���7w�3�@Q�Ių������߂���%y�i�J�hJĔ��_O�3�z;�x)���Vl~p��%�����=�	N���/ÀX��]s��s���t��S��Z99VSGSr��ɲ�]��^��+� ��0� 5��Q��~o��.ߔ`��-G�pm�!k}P1}e�ҹ��\ά�p�J�����3�J�z��s�ш��WrZ�P裄������@�u��yb#�5��g���ە��s'2OY�I�I�wjA��<^�� �t9�#�H)!�����Ȉ.t$�$ ��W3�Ӏkx`�By��]�]*iK}v���ο��|G��\YZQF~����vfL���o��8f�;O��k�X�DU^.w��?08n��NZhV�{�F	��,�
�8!Z�q��W��1jKtv6�K�/�Q��+/e�	��<��,�ʦھ�X�,b̬��`Z]��ᴽ�� �������Y5�8� �S���16���r�-�ڼ8�.���U�'k<y�ug���T���S�N6�D^��d�<r�:�%ї�5G)f�ɇӚ���$�v:����=n<ոV5���g�	!m)�d�c�՚%���e�@�%Qѹ'��/�Q�%wv��p��eA�� 2�����8e��kҷ�{�\�tKȎ���cN
V_Jy����6���k`	����d-����iyK��_����Ӛ��"�~a�C���]�}g�8b�A��)��"f�]&Mpa�;��N6��7�|`e�g�Ҝ��r �`{l)(�X�I��X�������+���m��7^g���������c(�CE.e�����_����͖��ZvxJ����=y׊W�dV9�p�&���+���y����(ٕ���v�B�����e��"# ���}Yl�5g��� ��>ۈ�#�/�^l�y��1��("��x̻!���Q�t�Sa * �k��"A���rdzPvwSR(t0/(��Y���d�>�Ϯj觘d���,%��C��>	~(�Q���_%������t�`S��c�< 㚆̖s�fc8)c�uS�2����{l0�¸:�����G�W#X���F��K��D�]}�.m�,sZ��Q)��N�@��f6�C%��Afa�/{2E�h��e�f;�q&�u;.�dЦME1M�p!M���t�\5ÖA�����[��K�+5�
��^��4�$Ȝo����4Ὃ���
i���r���eF�%��r�����8��B��q�(��/�,J�bx��,΋�T���š���c�a��������w��'I�]�]��K�Q��`�#/G���7b�P��#���"�lZ0�N�/\X@GtOIiP�1�z��,��4D�#����d�xj�[����������X����6}A��K@�*���=�g4t�i{������D$���ͩuzdц�ȀBk}/Ӄw����D_�n Aڙ��!_� ^ʬ�.Z�<l�"�3��D�<ga0�lZ4j�j>^!Y�Ȁ,������7R�I	j��x��Ҡ���� g���Y9'�~O0�9�a�@9x��$"��޴��.
�NI�Db5N�?�"n��~
n/����f���&Q/�p~[[���2��$5�=�.��*4L+���Qx0���4�.�f6Q�>�x���Ź�9��6�~@ʅ�q�J1;jZMJ=V(����{L�_e�p/ �r��b�51Mئ���+&&]�-o���a������>�ͱJ�4�����-�f��{;��?E�Y�2 4��7A���iH��>dH��Aj�"��r=�Y��%o��$�RQEc����dR��!�#A�ʵ�=���ƻ��A�1���1��J*�sУG�=�}�P�8{6�g�Y�E�t5����!�oX)��iZ�C��)ƶ��YG�0��E�M���QJUn�¦�[J�/d�_x�A��	l�y�v�P�sH'�A}~AB+Æ�3�Z_5@ҷݥ1s=��KU��g���G�,KG\\Ln��ꔁVD��'�������'s��{pi��FC����P�Gp,i��Sy��}`��S H��
[Mad��� �H��d����A(V���f_�#+�7��V7�"(
�8N2��,Bs\���`=��:~���#n������=
!��@=��X���̗�ߘ9�Tj��c �i^�`�l��D6W�������{R%*p��z�.|b�D<���,I��o�qOxȯ�C$T���݉xֵ�T\��� ���J ��f���Rg!�� u u/�1���ڳ�Q�a_��+�vs:�z L��r����7Qh�%IJG����?��
;#��R�
%G�o]�'q!e2�36@�4,���<#8�I%4]����,Ĩ�#9]Ym�}��/,�0�˻Z�p�ӹu[�˔D/��-���	���z���/_�D�{z�o�
 -�;P���j]ɕ��V7I-l��?��H8����q���ZG�l�F�r܀�z�3%V�V+�:K����'�������,vG�~��%I�V��?S��9I.6��RY!
{�g�t�_����ȁ}�3�Al��Ӣ'�%p��b�'ܚ*���Eqd��!�^�V�i�AHc��i��5$Bv���)��@���rQ�G\�.�{��3F��T���,::�PCu'���wu�h�,(Œ����;[RV�#��BA���u�ϠƅQB���㞰@XT��tn<6K{3c>\C��|짂���v�SŹ=~Hl���)�R}�gy�A�#6#���*�孭�x��vG�%��^n�:�I�������$*M~{R��T`��yW����ʵq�v���D���<��c���w��yv���H��J�R��7%�x;U~�R<�3�5���ഀߺ�cX{�^5l�%t{��!��� �ݤF$=w$F�=�l�~i_#�]���%�!����Z)����9�U���z��o���G�b������?��J�)_po����ANJ����0U֟*��q7�msP��4�R��h�Hݼ�L���� ��A�K�l^էn_�	�'�[��=a�P�VP����c�w?��a�@-���wl�ZN�# 0�l����l���"l�C�%�2����#9\<M �]�K��wy6�p*�N���1�Ņ���9�8�;B?.]�_e{L!�XoD[;�|9�u�]�9���dB��nj��
˰�qN=刬M��ۣ�����qؖ�jɩ���
��	w��e�&j5)�'�t)�`�a^�>zf���WĆ�g�����,6��s۵"��uy5ǹE`vm�J�k�`x��L���W2�0�&OOT�#`� `E%�l̟��ʟ�F��xf��u;zҚ�3/��Z�n!YKG���������d��2�@��O�4�b�0~�����.蔕�|���}���sSt8;���z8f.���޲���Թ�=͏��/7e2��ڭ���X�c��i�*�h��h�^�#�����_'�&��L���A�en���kKC�]z���j�l[LMw<�7[�8�Cr3+��x=�A4#�w�> ȑ}u\��p��u�e�C�=z� C׆ӭ��)Bm,�a��Y�ʾ��������������9	A���r�Ւ�0F�tfW��
#�6�\���	W<�z�2��\Eb_7��%~�}�/������#ָ��ݤL��T`��Ų�ښ͋:����n%����Y�y�E��re���z�iZ#[�K�ʇ�e@Gl���nU��4Q�j�'ώ�+�!���A�Aoa�����1^��hY�i4�:��v�%�r?��6�M���L�?�.g�7�q?�?<������K{�A�ND���@��Qt�Q�Cxq�\?[Y�C#
T�oo�!�ɴ�n�x�I���.���Y3KG�|8:��� �P����gB�	3�d�_�sa��x� ��UcTvh��J���x�o����X
QJ"��^+�M[��G`����L×�/��*����f�J%(�?�.Z{�0,>���2:$��H������'Fx?i,�:q�>��v�"�lk�7i�)ߤm�J-�t|q
x���*"
����C���s(cʷTM���p����L%3n#�oΆ�����ߣ%�O��@�f���eYE8LCIB������^�br����	v���?>��>9I���<r���fٍ�ŨȚި��:{.�+V#؜Մ )$3��w���܆ Dw�"��ܕo����-�k��p� -~
��
d��+�B�͂/��	ݙ�(�/����P�Ϥ���ݍ�}{#�V�����wIVl��_�l��"ǖ!pgf\�h�O�m�"���Y8��%����\��[N��Țg�� oɯn' �Z,u�:�*��{	
�k<Q�Y��:Y�W�2��_�:�B̗�g����Q2h��X�(W�{�6�a�/毹i���K~|�9R|�y�U��L�t�W��Y�vt��SØ���|K��)��~�H��鋒e
�a�b���$ "},��]=?�G�,�H��4{E�sU{5�v:׀�n��w"��iUtZ|�֨v���h���)�T;�G���\��#�2��4�B�MF{ ��f��6���oP62�Ff����mQ��\e�h�(����\�Xu��i�`�cnt�Z>��'�!�G d����7jٔeZ�z��&)	ɐ�)��*7~�kS��<��i��^:xo��<�'���8?L�krY��AR��M�~m1?�{S�TE�I�F�@���@�v6#�K(^���$wxQ�Y�����w�b��oBy)��`����
��.�;�Z�����
�Fm��|Ըt����"Y�mB���v�$l��2ZG~�%Z�w���7�Ǧ]������e�׹��P�wp�h�z�P�_n����lQ��nI��)��?/G̚�9Z��|�ċ��vۚ8�l�z@�X���6!衝c7�"�&��uπ3��~����M��	)m�M�M���XG꧚��SDu�nZ ������6=�����N_�:7\=�:�D�e@'g��HC�O� �gw���ZRL�K�Ls�nT$1r�tZ3�rW�U��L�f�h=��tC�}�M��[Vƒ�n	�@f��,'𪈁K��eD��� �L,�Z��d��="�a��&�R0ע�J������q�ꮃ���da�4�A��5E��� Ɂڄ���B݈�G�uvA��#��kgsUۡy���+�n!�t+/��S��q�<�`�i����(��{�E�yt��Ӈ`�"/��G'�1*Ⓢ��	䕱��z�`{��B��Y���
:28.`2�����*�T��v�l	�B�� `�����@3G�pD�+�2�����z:�ч��T�u���.�/�w�͖�#j��E��.)3<v����*ȟ?�k��aoF$��u�R�a�&mD�#~lRP�e$]�:=x�RIY�بX�����BI9�C�t�C]x���ɴV�w���Q��
~A,x��beM��{@��ےDuʔ�ð��Z2*�f,�a�|��6����a�����K�	����y���_*G�^|���̻��tB�NI5������6xѺi'��%����N�v7�"5*���lmj�?#4Y�L����!V|��tl�=��k�|�z�*&��z��k10ЋՁ����^�]�W0n
L�M�EF��W̥���u׊��2y2x�;�lBd��[������K�r^�n�_���δ��:)����W�I	̀Zˇ�����I^������ҫb3ݣ�.Oqk��i,:x�s��Z�;.�����;���SL�N݆T�)�h����R6p,9���FǋKc��+��*+	͊��ʟ��- A�հ�;N��j�7�cr�+[p��i$A�H"o�t���1���79�3����'����G�:y�6��@�-�͑tz�����n��>o]��d�����,G)�K2O��w�������ZX�������J2��G�Y[�>:[�L����}>���b��d��f�����^����Tڒy���c>�C����h �o⓮Y���/���ñ�J�(�%�:�A�wP+s៹�`�V�>Q�4ʮ�U�b�+��N�"V1 ����B!U9=�!h'vݎt��<�P�s�Y;GT����U�撚q���(�2;���Q�㽻]��W���&�4|"�[v5�{4�	��fԟ���U���m\�%5�`�F6���;�S���,��_��ކ��S����s�T0���l)ܺ�ڧM�*��B�X45�v�D&��>]㩓���+s�`q�K��")q��}�j�B��#�꼂�wຸl�����J{í�_�惓Y��ۗN�z
�CA��l�l2/#��A�w��H��8��'���C@#mE>f ,
���YL#jM�Pp��FU�����h����{�XE��I ��9�u�]��w�w�l�m�b�ѨM�� ������nv����{x}��$�m~?w�D�jR� ʆ�#�Rɡ�c:�G�i�ꃿ������8Kz"9�қ��M
\J>}g�Y)�E)6�Wq���;��sc5.'�8�#�=�Ĳ����(ו �p\)����� `.. �����Y�����Aw 	MRe�c��'Y���f���a`<��Y.���
4�ȟy��b�d�}V�7�JRJ���!|;s���"1�zh��#ׯ�](��"��;$uʼ���a���a�9����I�\����`�߬<	8Ne�/)�|n�]��%C�m{��(E���5�ò��)a\�e3'�k�fO��$�q��݄�D����$P�����=�6�yl����TZח�Æ��.L�,!�������%ݿ�z��.��&��6��F���XKo9�"T��>`�7t%=�@r�1��Zg"8
�í�u���T�yGB���~8�ԗ�{�X¶��o�î�e�7�W:�M-��F�I�W�$��)��0S���	���Wy0�ʶ���Ug���0Y��C���^��1=и��9��G�vs��ߖxS�0�/#i�G�	�q{�(�.�gD�)�5��lg��e��[U$to�� �{Ѱ�p�Q�(ӽ%a%[�+���E:�g��c�>=�9 #�5��F7/
�R��Ǳ�q�]S��{)�  �h�'�;4�sv4�ˑ���EF�y.�@;�E�jX�C"YL�Z���13*6^4xt%�֍�ȍ�C`o�V��{rZ��k�+?�N2�A��ooY��!	�#���_�7��p�:""�ʣ����� �d�^ �d?ф���Hxˮ���8������#��;�I-W�#`�,�`�.��'R�w �vj�ejS�ڠ�3u`�Z�'[
�>�i��2���H[llz	qC�0T-��������M�v#��/�����Q��a�׏I��ʭg�_�D0�	���Iq"sy� R� o������~x�Uf��F�Ƶ+�)p��f�@������*�ќ�a4�0v�& �f�@���y ��D�a����ſ$����[���I��A�����%��l�O��p^i���Iw~�Z=�7\x@�ZC)~D�(sڔPg_��`���!i������{����m�p-¯��d�(+�ih��ϐ]0�$uf���HU��xR��H49��p1	�M�i�����z�l9B}g��u6�怴B�����T]��B�c��>�p��_Dن,�Mo�����ѣL+����my�ȹ}�a�W�o�|>�i�����%�AMo0Ԛ�=�]0����̅MV̟H^}z8��,e��H"�;�og([I��(�U��2}ʥ���Ns?��o�d�RN�u����"�R!��%&å&�Q�����^����n	'��D��Z���d-�dɫ��9*\P�N�H��]^��%�nL�yV�R���.O�!��y3�&��U{/��T��3�r2��e�G�T{c�8��}n���,���bK�.�48���H�3B�UC
������l��&(gx&��?���e�S5|�y�>��j��e�M
�@4��P���Heur*�و����1�,"­���8w�����cA�6gxu{���84��,����(z+y�uia��&�	ƽ�����v��'�����ea���;$jK�.�w�E<��d޹-@��	�i����+@�|��l~���<���4��`�Q����:�yiI�L�E��}�Fۧ;�	^��S��6�J���6՞S�������;���n��H�يƐ����&K�G�*����:j��v��YEGҋ��73sR�f�آ�ZkH�̞��`��%��!c=LHը�Vh�޿�L#͚��?�޻���!�H�i� �X9�$�����!���y�-�=bGI�Œ��vR�!w�쪩��E)O��{Z�3��p�Y�_C:��b@�[�ּ�A�,��j�E3�=��a#�3�sL��3��Y��:������@�w�/`��?����.�Ti�46$y�q��TR�G�;��lг�4n>��Z������@D�B��"\�[պ�((G����DEVz4��@P���PE���	�{]�C�|��X�Z��E@0��D��g�Jg�[�Re��p>2�y�!^��]
�΀�:^,�S}����W�wB��fʸ�Ex��r���5�$w��j����_o��ߙ��w���>����Y�d�{"���N*8�p�Wh��s���ظ�o  w%q�`��ɋp[܀h]�pVݦĆ���C
Ac��c�?,�R�1|�d�&t�� �����s��,�\�_��Pq�|K����p�&��)H����
8��m����V����^�ލS�o˄�yLgW����8!��ިԳ��e؎p�@c�i���uA�J����s}m����/����z��j���/Ԝ.%��[x{/�k��&�:D!T`,ݼu�q��å;�f]lH���j|~�X�`�,�&��+��J�V��4��DKx.�y*z ���3��nZ/�"
Mh�i��S�R��#�z�,Q�B6E��)�����H�4b�8 ���ej�0�g��i��u�� 3L'^��h�ڣ$�ypm���y������΂ i\������t9���Cb%��m�m�IQe+��z�:k{0[�u�wД�ែpi#.��]��P[O����d�Y
/�(��y]�
K���y�¡�03�9;�.M��좳4;��m���iw놁xC$7���K�E��yZ�I8��w�k��w��~(m{�T&�C�h(������G�a1ʑƴڎ O��g����RNס�)v�탦h�ˈE9d��ԫ=J�Bҡ����iγ�Ĥd�qٷ�k/fC����tH?T �<]�u��m�;�R�s�b?�g���1ױ�	�{wv{��s�vr	l�C'B�'2,����E�K�͍�엞WP}��ؑ���z��S�|�r����Eݲ�z�]���^o;�R�pN�,Ԉ�������go�$*v���9C��軅���d+�	!�xn���Jϴ9��tz#\d�#�"�r��(ćs,u��+��-̰�+ !v�Q������(�}�Q�ί�1�>iJ2e�OH$�j�?(�Y��
��b�-��}��o���E�b��%Pm7�f���B)B}>zg������l��q�e��A�`cu�џLXn��j�+�/��MЋ�]y�y���My��1�
�;���|?��0N]<�Wu�k=�by��\��){X��)��P�``�a���z�wa� A���A�'A�p"Ƴsý��V$���Y��b9��������]ۭ :wm��s��I]0�@,} "͸�H��N?%�h�����;T��%��ݜ��sI>���r��d��sM����<��<�^��l(\{)�/��?b������@_d���:nn�$T���l���}c=hQt3mњ_�D7�}"rQ��1��p��Zy�o$X�ZY 0In7-ƥ��^���%zaD �-���5�
�\��~7��{s���c��Ki�5<L4�A��,��`�@�&1�!�Y�`�Tk"�N�
�Ny
�Q�\�֬�JB-v��a�xр=+�v��ox-쑁���){���������n�1t��]���g�Q�³j�39lq?��X�,,Uwƻ'�%�蕁]t�B�|S�x���*流�[_�s�Ag���&2_�u�i[� �p6��(�y�2H#�jw|H:�t�٥"v���Q��X���$��I�4!ӭaQ�|X@e�?�.��oJ�I��{�%���7<M|`�q?�7���T��R��G���c�T(Ǵ +S�q���"
��N��ٿW�x(�e�h�&�a�d�
U��3��7��k���Zg�2�akl�EU��P��m�de1t�G_�b���Y��o�/�_[����5�*�\�����b�M4��m]�M�{�bA|���-77�c`��\�Q�Vu�~�I���Df���3��z���q �-,���Q�]�&�tqc�Q񤚈�?g �8�e��d��S��+5�I�\���t�
%C����[jL�6� .Ő�M����U��C6�}X-��&D3��&�Y�/���� ػ�<0��,o����0�����V�H�]��-<d����E�J��Z��
�:;�9)],�7؆03L�h�/սX9P��S�������;9��y�7N�����V�{Ȟ(���Hd�Cۜ@�E�yŊ~���*u[�k�aR��k[+2|э�R�C+#'��es�K���9�N8��g�VW]��ٻ�CF����aj�C�	^V(x�|Zu��S��T�1�:�$]�$	e�P
�D^�2-���}�M�|T&Wm;�V>5Ӷ���(�@��7����蝮��X�Y�{�nb)��{�ǉ*lD��7���\2�&�dATt0��́{��F����Ub��3h�t`���JC�5�� �㴊3���>��[	����H���?H��Ұ.^��^W��[�㍵�O��V�<�o�12N���[�|?�Vr����?;���'x����eWP��EbA�@�r�L�МaR^8������\s<���ɠYa���H����#�3?��w��Ӝˌ�j���j�9�h����_A�V�}�g�{o�ϥ��>e3F��#�jR,���q�֋n��l�A�,�����S�����RS���,���ٮ�:�x�(�~;����\��y�o��v��f��b�����������@��j��(��F!�� ��=C@��Qx�~�A��TR�*и}� }�I8R�gc�pL������.﹨OBϷl��A��
�{�.R��/�_mI�=�nC%6R��;QԀ�`BZ�l������߭�#������Dh��9Q.�h}�	��+��Jc�p�mN����{��\�t��+kj;X�ۈa�:�����E�D�����
�����u,)�Md��^{����I&םj����K{�lб��,���E������^�������bo��R�,	���h�e�����~�;ِ%����F�!�p��U��0L(�=a�m�;&T�T+��z����������L�]���K��^#�o�¸�}�-���x0X�L�m��Lҹ���rՕn�C$a��G����'մ-�b��3������~D�/��7U$8�^(/��b X���a�B�	�RƭVZ����U����x�Ss�b4jv��0N����.6�#t�+8�*�+�P'����%J�d�\sW��`6L*�{#�z�~���2ۭ���[���H�n�ּ���h=#в��x�17͞��C���C�:���>�ɬ�3JƠ��T-�8�*&��+܍D�3�2b+�-C���v�Ah9�Z�U��{F���r���i� ̒�d��e,�ږ>A�n4@J�Lx�:C��
�<�$ŉf�ױ�0`�n2?tA'!(C�dc�R8:�T�I���x0`��%��F�d7\
	�!@��s�X��Ț��ؾ<'�r�Z�~�}T����)�vP;���c.�5�ضv��bݪ�^�z6}\��KTt��8�R̵�Po�N-^�b��F�~,�u�������*�s���(T�Z(k�b�͝�xe�5��wUE�[@�N��@�I�L{.\��ݴ��1�D�	n^�Ma{k����Ùw�M���l��,
,�+�fBM��k{�����D2q�!75#Fp3�+(^�6���0D��L�fs�<�¶t_����r���
!5��&�r�څh�%�c�5�gһ7���g�]�\=K�@r~G&�(��p��0�YI���a\�.�K�=nt���D�z5{99�|
�~*�"�SV��SD���Zې�*lSP��@�y_�+�cY��|��`����1G���*t|\�p��7�M7��%eo��	��s�~�7O��E�wJ[C@��Έ�-����nv|�;
,�N�5_��X�'��3o� ��\ �[AZ#c�!h�:e��cp���1{ ����\h8vǌ��$D�i���
9���:�뢥�T��eE|�$$D�<�}��_�i?�)�ө��C�Ȱ@�U���A2<��\U�w�0��&k�ռa�K��y�L�f0 �������l~�yЁ\�h�)�jKM6O����Q¾�qi��I�l[�Wc������+~C��/�i�����rb�;����ˍ�����0�u��Uwj���yG��c$�;�����@LZ#6���� א�,�������~n��\Q׻p�ⱨ CԸҡ�*(d�������[�-!�*(ˬs��;u��êW ��	�f tS�a&��vF�P��:���\%���6�h�lА�*�"\m�ݾ0>l��<kJ`w͠��N���6`b������U²���:�ݾ�-�^*ưwP
D	Cad`���j�-��V�l���־��+����Z=%�@}��M�vF�*�~�] R+@�����7wN�F��)*Ȧ��r�@Wj��*|�H���`�h8�g�v�%#ݖ'�U��K�.���C��|�Ŝ���`m�}W:1sP�f)+F���-� ����[��`������	5���j��"ӴB�؀��)(h�z��΀.����F����t�v{z���)�JP`pF5� �R��mn⧷Zú���07����p�DA!�jA�4���-ԑ�b�i�փ�2�:/1d�h�ӟ2�����~/��ĄV0���'8��^ �w���&�`����>�G�z�ٴ�y��Y��~^JW��֌.EU,Y8d�w�q��%ے�i=���\�	�����$0�r.*B�O����,��)#"n�P�m{�=k��3/r���������4�/��i�ёP7�vstsD�`��4��������1��H�}�q��B^,�
���M=`��hŲ��w{>M*}�y�n8>.��h.����2�d)�Kz�p�~���y�����h.T�8T�B.�����5��&��:����<fV�!-.�E
# ���	�����9��^���m鎀Ĩz��
>xt�M+c�4�J�m_�tz����,�������]��]LA��
�4B���\�cE���ȕ�2�d)��y2��)}��g����qQ�#@�}N�|�*���w�m3�4I�Rz�p6���^e��f#*�'��ZM�1J	�?���m\~Rxb�+�9Dqd�$h���7]���&.Z�c�����ۀ�A5<���ҊH:��_��_���0��F�.����N�b����7_�9�J�s�>P�|i���ֽݑ����m�H{Ѓ���S&I,�"�&�9�W��f`/N�Ɋȑ�%�8�N^�n_\� �I"rß�i�|�����V�=�H@n�;�H!��H�=%�񉹾+�NB�Nnއ�L�(i�u������*�x,�@6>}�a��;J�ۉ�WQ K�m�q�q�
��D}LUQIS2Jh�Z���]xk��=��}���h����+��S���]+%�������O���<�-��k�Wף�$�!IDs-Z�c���&����@�-Ţ	F밺�F����0�9]�Gp�V���"���a>B��Y
�?�aio�د�
t�+��6B�㔐g���B��3nh���:���޴0��SPG
_�N�X`��l4@2k��%�f`o�}�Ìvn����œ�����n�.��H��K�~� �����.��!F�+�%��bW�4I�O**?n����h�Y$E>����:6\�<�.��H�q�����"�:���2�-��"���L���+J��o'�U֓�W�_�3�O����_]�0R�!n|� Eєx�����Y�g�V�eZ�a�H�Mh��Ԁ��n��5�&����X�̊��O�«���2=����c=��MÉ�TS�E�}km� Mo6Uo[�ëe|Dc�oG �c�[d��v��#��06@�(����Ȇq��bR�=>�3�aV�^}b���Ѽ�Ј��&]cU�r��.�^N�P�*E0�Uyq�܁X%K��Y$�����ߘ.���N�T��u��3vTz�a�uc�[7��"�t�:��6�����{��ɊAM�-^^\�{�ᙀ�A����^M�����g���m�c�U-�G�rQ~��FI�x����0"���iY�nHy�[�H8ڞUE��k��|��/P�c����A~c˭��e�w��K�Xt���$��<70�/����'l.s�YW+�;�a9J�����ҥ�%��v.��3(A̓P�����|��k�8�sm8���#]�W�4N�Ԍ�g����)�k[-��9��1�k�&��f���Ᶎb»�Jվ�J�T�br�D$�����!����)��E�}��tਐ�>����zo�e5���>�z%��\ ���G:aí
@�2mR��f���'��Gƅ��v�Q"�kK�k�ɔ'rT( $V[���3. Y�C��q�u}igx�|\�yE�N�N�z�,��($�kX>',��K@�(��.�<F%db&Oug���ìx�=�aH9�;d��ag_�o��U,� ���Q��������gbX�1���� 0
����+�I�"P۶��a�2?Ĝ�� /���)*�=�;�C,��
�$I���q�=J�*~�F+(�n�N�hFb�0�&���\N�U�"�1�c��fjX��;��J�Tf��͋;U���>��#ˤ2�w=������F�7Bʵ�]��t)]\�T�Ӳ�w�Q�N4�o��8)����m�Мw6@"�0���n�z���@Qq+ڲ�~��@��5��K�)��z;���B�9��0�������|�V�!�˳J�_`�>5���7��ʣWMs�8�#	B+�јЪJ4��̧���⌛�4���ݒE�fƷ��ize$a��s��E��t�q8��2"- ��XMm���F��U�3�[��t(:j�^�9��7:�˻$STJ�*����^�1J�ϛu�Ɩwt����W�r	gVw��p�����`��#x��u��QqR�:nC�{K�)��y�����W�t�=��i��ىу�l-���vB�a(�TL/��s���؁���OuC�!�J��h�Y>��^Ӵބ6�MO>��ܚ0ƅ�<0��T��[=h��uwi(�q��C}t˫�~tA�������&� |yjއ�e���%����q�^�����
��=V\#Z/!����I�n�<�}ZMZ4������8�|�vADr�|QG�s�Ic�"����it=���$p^ ��}K�v̱f����~�M��^����g�sdz���}Kǉᒬn�"Ji���������1�.-����G��=�|T��Ok��&Vd�j����ӿd����m@�ڶj��YK����ta���n	s>y�-��x`���>��@K��ڍ�l��\d���}��ؐ�dc��J�aMg��H�7��i�ĩ��:��5mp�"�V'7�B0%�K�h9K��'���%y�_��j��i�W�#�*SGxm��2}/�����uӰ�V�/�
��&�t%���h^O�=��&���l��0���M䚄���蘼/1�STO?�P=�
�$1!m:��bn^!0E-��D�ѥ���4�RDgH���B�?T6x�3�-.�H�SHٌ�]�n' l;��)	7�4Jri��>����_�)r��9-Rcx�΂��k��	[Eu�U�\I�@� �P�����d�'M�r��l��H�m�����i�I'
N��G�Gr�έ6��R��{��Z?/9z���U
�A�_����$K+al�"�5�W.ۑC^�A�t��H@��U�I�V09p56f�P!/���qEa��~z{�/:iҞ�&�g>!#.r�����(
S30�L��O�l�T��(�ϟ�<�3���,��(q_g����������ʮM ႯFYSa�G*��zF����Z��I
"˼,C�E�[	��@,&��t&���\�h��>�a|N><d�]Cp��Fz�$c�"N�7�]���V� N�c�u�����Pd��J"�:O����D�\Q�)O�Ee���V}Fۂ&�r�Q�XZ�5K����|���~ڒ���MP��M�Sө�Yt�� I�w�,%�#O*?wv�ɕ1# ,�9`�'�l�^[�@�/g��p�M>F�-�� ��Ԁ��׳�Y��~�W�� �\�����7���@�H��V��q���H�@�W�zl
��n�7bV������Hww���<D��~d�>�aނ\Y�b�w��/<�78薕����Ь�F0��lM=f�X�w��ju�5�V�R�aa��!�@=�2E\���<Y����.������{���U��k@��|v��3h�:r���Z����3�n�f`��gc\Q}p�<����Y�9ESE^���?�:~����g�����|'��veV&t��fy�U���0s�(@���-8�{��L��AiE��Qj2�٩����Ɋ�!#��(!e����-��q)x�L�r�L�M�<���V�Ȱj���y�T(��E�!}z���jc�P*�K��]���me��7��V��D��٬]���=�2x�:��@}�W��%A��Wp���ZͿ��ϔWe�mTq5RI�Uʊ9U�����H�dk�@zA^>��ʎl�=)�CV�Y�:P�띾��R��i"�R��9~�R�����vb7x��ʲ��YM�#$���	��͗U�����J�\o� .-(���̔�{�՜�;�ce�c3�9ʄ9#�`������r��U�NDվH=��.�K����N�Z̳�U캪��\�4ƗS���ʓ����æHM����!	ׯ�b<��L5G6��/��asz�+d��h����a��I.�N��-�T�C
�����Q��%X��HpM���9�n}>�՘�U��Ӽ���V}/��#.ؤ����+�l�ǻ�������A��/�7��!�w��W��K���OGb�̥R���)e�����ٵ&��~����EtZ~�n:�ݧR�0�7DmN�søK���I��,ٔ6�[�8��-@jxYSf�%�^	u�/�a }wrL���+w���T�<�'V��~y�� ]�V)���w�ct
��	��F�?��O�!��\Ob���gE�_uw�6���F� �'Ѽ��~��iB�0%�u�o(2���z�lU#9K�{�Z��C��}��(y}�P�A�$�!���S&�oI�1�@�ڍ��2>�+{���R��!���,�,�u�!$��nP����-��ԟ�&�@:�+_���~1�y&�b�H̘,��}�\zr�c������k�z?.QN{-��.�s�@��I�ء偫�o֍�C����q,�WAZ;��i#�l%�d�N,���ݲ��!����
Ζ�S�)^��֒r�7��g�CU��k�/��t�=Q��������.ަ>ȼl��v�N �k˷����[˚�uhh]�1]��ോ�6�q�=7�^By���;��w�˫��N��5Q�"�D�'v!ߗ~Q4�1�A�[U��$j,���]9�j[�d4!�e� �p%z��M*[����Ed�o�o��/�%�[B>A=���L�:3��L�� ����p]�X��?|Ozݍ���gO�ٮ��u��o�߹���W��>������t动3	i�ʹ��DĪ��S�}�/�dY���@q":�Cc����Կ�������)��Ȱ�6Ů��F��C'�@jƯH�u�)|��xc--`���=�C�ݎ��ͽ�蘳��iVu���PZn8ٻt�0�e�j����o&�P��b`�N��9hRE�m�`���Sy/��A*T�{O����\�ǭ��`�ԗ�]��夽�,v�IRr���Ո$��Sh�<�O!���h֘3y�@���ԪO\U�KO�]�>%��I�N*����Y��d�At�2��R�K-�D>��J��M���>�Q�z�]X�y�	.���@=�|I"�:�<��<,�ⱸW�796vj2>0�&3i(Jf~U��;DNV�N��<=*~��U"��]�`L��� -$-���eY��1/��T��dB��~�nL
�k>��ZRm�P�ʛ��U�C�l��-S�c�D��������J�M��"��v��MX-�b~��4��*����[��E͐_A�-�x����%�u�˓%�6D��!�����*�@��� ;$y�?!d'��-
��
:v����ٙ��KK]w������G�y��#)�n���S:.�+Oȳ��_+n���B亠ʟqw��	��%��ҺZM��:<�UY�
� a���C�T<��a���#���h��T��⛭�bX�Yc�M	g�� ����tb�1|�؃d�@^[�yQ�>�]����Ô��LϨ��Q��	�*��7�8Y/ h�U����Q׽�G�'p���+�ɻD��
�!�ۋߐj�-k�U�����ׯ��A�N�D<�~͉?��L�e��@����F�b��I=fI��<�׸�Lj�;�d	~q8��,�`�U?(�_,�;�w�iR��3@y��8���N��|���OQk�����Qt�y*�o��p8��~���"�~�q��5��M��oC�o���� 4zR@.��/n#�	3�����#֧��}%�v3`߁�9ϡ����y�(�ו�d�z����i���O���Ԧ�7o�/��7PM��g��=��v���
a��c �/a=E�r%�V֓����i� c`ޅ#��1�pʚ4��D��������%~<+��z�PQ�(��֩_���I�&��wχh�����V�Sr�����-=��K<z{�]�57������3G���I�~a�^*�$f�rE�Y;�f�z�eE8��<.E��A�������1��C�`(Y�=�	���og��o�&O�[�凹*')��~cNdf��v1�zR&v���ӥM�:�¦� ���u��åE�/"�:�'�$s�1��AM��	O��Ĥ9�_�ɚ��Bc+;�i����g:,��q�����Ԋj���ѻ=�K-B���8R��})�[�le˴ͥ�� ׆p�Ӧ�0o�{�Q]ug�-]���a\��/2d�`T1D���z\t&j�skƠ����裔i@��r/�A�\4���f�?�^���eW�҄� mHװ���$2R�r�LX����uZ����Z���O��5}E0k�
�=�5~+*���<f�3wXn��O����`V��۞����IV�=;��[t���j�C%�8�6�X��lq�6B8��|:	�5��ҋ��Y�,i��Yg���o �r�]��O���E��-�������;�����5�S�ѥ�o=j��-�k� ���T��8�O�f͇�#��01�e�h�s�X��#���Y��w�M�O�K�nR���
��9\5�9Ϊ?�c������@����r֧ �ֳ[���$����
�[]`�#QY���n�C��#�o8�X�u�8�2�Z���T��|�[j�m���t7�Sݾ{���e��Y�N.�Hɔ����5�Ym��:NV/���@�z����8]�>���5�r/�bz��vH|���Ѡ1�J��c�T���k���O��Ǐ���nK' ���̺��-z�\g�!�QBv�Pv�_֩�zDw�ES�A��B��D�Wg����*i��r�d�@��U����Z�́��J�o��wW�����?9_y�T���[9�uJψNG�-�^��lb�D~�����ϭ��M]7��l��?Эp#vS�:�l�����4ZFWIYa�QW��~@Y��
?!��R���Z@U�w�c��}���Q�3�2��XC��F:� �Xi�4�@9F���H�r�4�[�2G�I A�"�1����V���R�й��|��J�µ`5MK%�O��ԕ�uqXGz�xV�`e�rh+��u�}wm��]�gϦ����	���D�B~<(m_o�����̀�1pJ̵�BxMg-�%,RW�D�hm[���˫ss�+��t����S��}?���s�*y��2�Fۈ�6�`����
Q�:�\�38E� W���a0�O���<0.���Ó#��ܫha)���@EW��.yO+9�\��CC{���nN���4�Vqp_��Ϋ��\����R@�����3ߌw9��~����|Eƻ�qo%gԞ���D56����̂���PHݙ=�C��
�k�������A_[TϨ�����P�*g�1G`q(��MՙI)�ҟ�3��M������|��k�>�NJ-��Ÿ��	�DB$ѓ�!;5��+
��;5Is�
ams��?�
y���w֖$�Ҳy��M��^��ׅr��a��ڲ�����Jx��4+¼���+9��<^�Z�r�>3�QrÃԵ6|}��Ѣ-��9��9�-M��L�}��|<̜�6�L$�AH$*��u������p�"y�SD���E�����e��[�2��|FS���V��c��g��V;��{nF<>�����?��9�%�j���՜~�B���&Ɋ�[�����@�E��KM���l�>ճ�?蜅�@�;VQaz�V��%��Re%�w�n">�̒�|��w���TF&��5��ó:�/��%����s��\\�k�A��fq)�Q��m�	ע79L�.�
�pgKV�����(��E��+5&"0�x�$�ҷ�P*+MFG�Κ���c��"޻ב����0�Y�J���|�"� 9�0�f�@�֫�]��9��w$J
n��W%,�L�H��{h�L����`��=����d���qZ�YAJq�3�ǻ��C��3�;��cNQQ�� �|:������	�W��p_�ΦǬx�(įU���֑�(�C�E1�?�1��.vj��!�P�;q&+H(����B��oe@� z�R�(����a�X����_A��l�&�p�n���s�F�%UF�C�h/m�A��^�UZ?��W��|�lv�����O������AM��SY�0���
mM$f�{� J/y���Cw�)����wHle.ٹ��?l�	����V,C\
���� �z�qԵ��!Qp��z,�r�Alz{�8d��8g!�������M��2���׎pq�w����H�ju�9�Ȇ���ݴ]�|�	��<Un���K��sG)�-}7�#?2MְYO"�����Cԥ�(pO�U=�:%W�]�t�VO�	��O�Z�Z��L2ˤ=<*�17�X+�4�]y���YP����J�K1Up�f;��m�v�U�$�*r��ahDB]��G��o��Qv��KvD������K�_�������I>(��4�KG
E��lMkϙD�/��blSX��w�>���y7�9���ϳ&[T�/�AIҺ.�)���Ӹ,_�����#��-�W3��8y���r��?�I�,WL@mϭ�9�d��fA����R�ˆG�/�nh��ʖ�¢f�2Kr�'�onP�������O��I�8S�SF�q�`y�Ms�◦rnBobO.�P��M�?���3�l���&fYn ���O��,�w�q7"@�1J�\d��*��	�d|�L4C���/�"Tǀ��Zf�Ս�Gu]���1���`c�_��Ul�*����ձ�:b�J�lY׌/[.����U+ԩ�yq\�A�K��S�Lǃ�Wb"����5�̾.t�C��dfq�r���|q,��]�����>-!�tS��s��� Ā�1���1�2���=�Ü�.�-K�H�<���B���= �1��k
� H
`z�c�O9��%�͎.P݄���)ʮ�Bpe����A�Nv\t�������b�]ϧT	��p.�~8���R�jJ�A���t�j�W��u�g�?�y�;����"��Ț��l�n�����di�LG�j��c��� �7h�S_�z�0��}@h�1ҡ����mː9��j|VmB�>D���Q�L������q][h����M\"V,�`��g9�g���=3g��E����;oZ����z�KC���6L^X��%QH���ڶ��댖vd}�G"USȪP)�#�NIܛd'�L���r�bW�c}�"��R.%+�9X��k���[L����߆Ɋ�sx-`	)��Řj�����q��N��1�G���Q9P鍠�#Ʌ�EI"�?`��"Ui�X�p�ʀX��ͽ)��d
���p>!&0��K.�$7�يz��CQ���5bw�h������g#Nn'�C`~�>6�L�{�L-,T�Ѹ�T�+r����8v�
�B�qtUtd�����ғ�n��}����@�� ��3pqNK�T�ǡ���-c�>>�C?]`~8�Sp3V�����Y)�֭Y��8�������{�t]�	�H�KA}�Y<P	����N(�L�Sy�}q6����hfRfB�^���U���h�R**��x �7�3^9�_�9MN�9�kue��&$M���ǵ8�mT�,a��&��ةA�Ag�W��v^�5�Y�����@����Y3}�����$28�a��	X�1v�o9��F�y
)���m�/?6+Yc5�2^��
̘�A��zVe�����RZ�L����L��!=0�ߖ4�+��ھ�J7�Z�*�����>���Td���z���>��o��H�Q��lL� n�ņb���?m�],d��e�5��mW/�n|#f$�u���y��J��5Tʪ�Ω�lO�-2o��< ����/V`4tU��γ��_ 
�t�A��Fe���������Y�p��8U�wS���+`{���`�q���[kT1"�^�i��������횩  K̕n����9ΡX�}��r��	�3�Ř/�5��7q�����ۧ�V�
o��d^\��
�SѰ[��0p��M�����
��<i�yF�c�rw=?>���HqY��O9v�̽��Ɨߣ~�24�NkA��^վ2V����G����P�#y1�A#�^��%����z�k)���W��o{f��7ȍG� {���������h�n�	KB � �C��S��W��#�;���� �<~�0��&��)<\�h��Fi�Ebc�Yk�;���YK�����yz�����9���tO>P�2t]'��rn�x}6 �,��	��]��?�˒�P/r{�v���)S\� V���_m�����@��N;jhB{;��<�j��շU&�^v���v���uV�Ӡ�rd�� Lj�^b�G�oʇ��F��i��|��{Q�t����8xq�jc��}qO�-����@5�B_���&����N�?�T��eM|��{�X�X�w�Vq>J}%Ӑ"��C����j� ��R�AkN�☊�֭�Ee␝���{)3�ݽ����K�+ �nS�Xhe/�嘃�����������yE�o��-?�����Q�ސb{� S�i���W�D #�l	2�KV��D~��'�x \-Q�{T����U�����͝�V�T:�|�-��Fy���/����qh��T:��#�ƪ��6���r}p�J����d�@�,�GH*'�I)$&��a���
l��#�ObM$Y,��� z��ߤ�E~���-�sTs�\���n=ɬ��{I�7�6/�3�06�n���J���|Q�'����W�RFj\�?�Gd�l�'�X�%��ݸ��ݑ7e��� ����ւ�kr�[֜)�X3g����?A�\��V�]ʴ
�w�@�I���b���a���Qj��\(43��3���*�l3���y�4���� ���i��]�q�Lw��X���՜�&Y~������� 񔀺�/�M����4\�Z�N���؝�wes��j��<:���h���B��v���O�uk�
�ɯ5�YO����$���j�T�
�wٴ"��`j:�����{�=5�M�N�7ȶ��[q�p�Eb�c�!�0$�~[G����J-O��KA;�B3-9�b�b�x�KO��|��A�z��,J[?D#�ყ�,rH��?/���p��re������4�8V(���.wĳ�.���S/+��	a��
�Z�%�5첎��;�� ��j�<n���z	圆�y�G�S�(�A��eT2{�&4�-|�,w�D�#
ӝ���_MD��:�sa9�M��	2�9��q��-|�ƽ��=�P9`��~R������3����j������D��ecE��A2����u�Uh��4*��Z.v�J�B��`pg��r�"�X��Z��b��T �p!"�\���|?E����ƕ�Y�J�myv�H�bC�@���I�V���D��ʭm�@7zo_IB�'T�����`"����gt�[:�:���@G���b����W�cLNz�mfd�=���0���z��,����[�Y��76P�7&fKf����]lb�<��Fc�uou0���ir䊥�rޔZu��68�v�� � �7v�-�E��bQ�0r��u��duK|�;Z�*k����ll�KG��ٳ��b�4���D^'�5�C5rYCz���l�]wx;)�Ϫ[d�c����Z!Ӣ6EX�W��Ff�EG���,���X���U��ʼ���8��=�����6[�#RN6g���ps�5B��Yńv�݆M����}ɑ��2-?�m:m�U^N��S�3X��7�8�����n�7;��6���]x���-ҢƦ���E�2_Z���M=�) ����F��N��?Ҟ��4�*sV'%m2����)7U�e
�Ɏ�0̄��`;���9:�_��z�^��*�d!E�!<�	�J@�w!��Ծ�4�]]��Y��]'1�{L��*b�
�>A��/đ���� <4�ܰS¬�����g��?�8�?ñ��S��������]#�ƋY��2�����lj`b؟�橽8�ƫ�?z�]�R1z��D�`d�9͵O3���;�~J%��YH賖-	�����U?$}@
r9-Q`I^;;[���̮���x	���2����Դi��W&}*�J����U��FW�4J�O� ,R�
1�.�;T\����v�u�h:=��X��\����V��nG7�>C;"hki��<U�ۮ����q�H����S�JxǦAYc���jd��Q9O�,��yȳ����-��9�O}��y�O�h���bMP�jm���& �@sc��dk����	�6"�̢�ѓ25W-��*K�7N�*�,`��b״xR�=��=j��D%3!�����C�H����.E���5x�;�T��^��u9��ԙ�W;(��h6�����3�T|�,���b�݁���t��V�%�6�/�J4YA�׍��؋�A��h�u�p�'���L�p�9�!ƥE`	���+J!1	���p[�1�q�Q��������@��Z��{�v} ��漁#^܄��Ҫf�0��i!�r�m���5\�A�ջ�&�J��Pg��TD����#��'-���R+�d%EN�p�yYH�c�A�8	ИA��)�R�Z�mo�ş(���_�L���<N�co�� \�D"�I��VYZ�v`Y�-���B���L�\z�:�w���$����t���c��fP/،��FM&J[q٭pm�"�Q�E���v�^=Ҟ��,����M)'��>�p��ݫa�����n���+G�Js �z�zL�"�
q���]���n5�g
�7}�u�A��z=s�?{ص�$�B���U.��=���^ޤ7�y�����c�΃��(�I9@��hϯܾ��C�$�2q��w�G�`��Ƈ��l����m�rS�	d�Uˈ�;�D���6�4r�~���z�_$�p��jum���?�mcX��/��$�1�� �>�si܃������9�\�'�@=xLqأ��OM#��L	�Se>�y�%�҄��=���5��c��y�?���:���w� ɧ�a�єƵ^P.؊0mh��Z �#��������-Yq���W;]$�k���"��h�;
�{��f�9j=�#/�o �r��Y'��`h�8V�N�	���,��z��1O�E�����+(���L��e��[r	����U���`%Y3��oU�A�� .���p���ŕ̂�l���i5��lZ��]{��y!PX$N{m�R{d�Fگ�����]G�rP=.j�zp��Չ�O�MO,"61e�l�l[�Q����[ݧN��TFx��U��h�YW���Mg#��F3R��Q�z4cl�b\զQ�����b��|��(�iL���%8.�npD=h�@��S��'�[�߹A<��J�2#ڤv���l*�9����F�\���
=����5*�eA��s�iJӏ�7B]���+����k4�����	�i��~X�8Ҧ��k�dVV��L�j{�� 6�_GC"b�K=HyX��y0�	�l�&���	�O�'`6+��P��#�������]�N��iˊ.��
�X?�N(c�e_�%�*�|�����Lk���a�IT�I��J��� 3�/��׷��l5��l���k�0n9KN`ϔ�戰�L���5�P�e,W�m+W��cR����J�v®��:���J�Q���nb���ztm׸����iJ�0"W`H�:|S�i�n�s���2e�$�Ն\��nt��8Q��_C�	 A1��;+�e��Ą2��Rd�92��l��yP���{`�f@V�ɯ��|<��<���̀�n
�{��[�f��W�o�3�L8�nR��5�|�s��f�(q���,=i��KOו�`R�X�pŬ�&]s�@��z������ٟX��(O����G�:��aR$�WʲAK�륿=�=��JZ4nS�g�-O"�}	S�͌(�,Y��+�Z/�5���/�w������J�Y�Y?�v낭P�2�o�(B��ߎ�Ӹ$L{��a.�����s����0��6dRUN�k��:5)|�H�^9 6��6�1R+�f}�6P�a}~ʸ$ڦ��<���3�奈O74*�~i��PC���L7͜��b<+��H��]W�R{ڡ[[I��kF<$��X��1��f�QTawoA3n+ק������#�7���'0h/"�b�*�Y��V�IC��n��������W.�|3�����M��䧹��I�?MV�d
t��>}/p������;�ǁ�,�<67n�H��Y
��W9�%I'DM��M:Q�]Y7,�`����# Ju� �ʢ9�W,#2/(���E�%�o��S�����z$�Lّ6d�t)%e"�wt/�F�`�u([�pO�1��'�tZ�!�r\�/:�ǓO��kx��)�")EO�t5��&@mw�Ǥ�A�yHr�	��;����?��D�g4�<7ϋV�@8�1�&��{����u�1E����~u�7���F�3�=j�m�YpDn�-�v�!��)����G����,������ɻ��0_��Q,ɤn�y)�XG�'��n��lG�G��'dS��u�rH`k�ȬR�PD����>�6;�f��}�C���F�nS�Bn���N���}���W�9A�;��N��FB�5
&���bd����s!5P������㖎cHV���-@R�6[�{,Ғ "�p�,��]901�Y\�&�%!�V����M���@8�Bd�_���@����m����j�������'�[N�j[�m�5���)��f�3}�3�n��C��MN��O�ka���w�J����g������+}�C���t� ����+�ZP��3.��0*E�����ǵ��Ę�3a��_ ��JCo5ѯ��
�n��t�����E�����Ugߕ��?�-����m��2��7��H�:����Su�ms�8�1�H��ٮ��7N�=`�W���7�@��^!��yʈq�<}&ɭu����#W���}��?��3$e[�\�FQ(-xAx��|q��[��c ,���@
��z(O�2�8�{b��r;�[�5N�2'h r��� I�̉�j�����#6���}�~�f���c��XhB4IWh_�u�Ǟ��֍N����i����X�)[�T�����,o2��y�WB5����߲�ш@�3i�f���Kp4�sK�廷�ůV���sd�T�������I�Ƞl���z�H�4����5�8��L��FF�1���%��6b��8�G�����M�h~T�(��C�zjc
�����\��D���X�N`W�پ'�U�a�����ny�s���;J@L�u��Y����Uʁ������">�uK�_��?��@��I��R�U2� q��U=�#��ϛa;r�X�r�3�	h\�"2l�W��N���l�B>'Kt�&�ɧ��N2$��|��ܫD�b��n�����I�h�(d)T��t���G�Tsϖ0��\�x�(��Hp�� �<:o_��ejp�X��'p��D��խ�%����G�~�,7h$q�"� :�1P����CĒ�Rd��*+�y�,���d�?�%���
��jaФ����̩����(���}j���6uU1%E���T/"������I�ж/�PMGK�U�Au�Q7��6��Ѡ
����{�V����*��@���޵?}��P�]�K͹�حIh�PL��]b� �)+S_�9Dӟz�j��_����������خ���c7Dʱ/�#��	甇K���D}c/�e�>�ÿ�A�4"� A��nÃ��z}I��1��\�`@�6'?��-�48���KA@���n�R4F���2v0b]!�<"�)�G��x��a��%b? ,l(����[\K�ƟyV����C��z�*��d_���:�����M�#���`��xX�ь�f[�O��}��Ft64X�f�X1'��Lu�kYyy����kYݔt�w��뷣��y]�H�|�$ݔ�S1�E��;�ZV��1S=H�a�gF�W�_�eM��hJa
4�
��7�I-*P�=�A�ܵ���q��A"qy�㐙0n3Bi^0*H�	��5����|v��Qv*U���l�V+8�p#�.j�|�)�>K#g!Ǳg;a^�i���W�gAUVI��u&ߍ�U�+���2���U�#7_�,wH�WE826�#r��#-5#'���E��9i�^���9�`%��ӂ/����n�_�����ټ2޽lDe�7&y��C�|@��I$>>�q~Ur�X�t��Qb���ܤ2F�uD�i�Zz@OpRJ��|�	�~I���Lx��G_:�E�M#��Sw��%Κu܌��5�рrwX���li����Tt�kM�pH�wĒ:_�c4�*�I�
�B�c�Z��R��8�y��1�n!?�X���˜�⁾�X�c~�F����w�t?���ʨ�-�;fy���Β�6U*�8OgzE|/O/�!�;�����yܟU���f]�/�q^'�=�yC;�� "g3�-�4RCo^�n���d�3 ����O5��o_8�3��$������\E�A�j�m��ѶL�Ȥ3���@��x���h��/իH6���J��hm6�p(��g@�� Y}qq����y�ԏ�Sk�/<�d\����O鄆r����e���9�&;ڷw�|�$�������9��f�=�b�F��>����ۂh�;��'��ɞ��ڄf{8�V�p����ŗLT)t5$W��8����x�7�(��~��3�to�dU��1�n�d#�EF������o�W11�͟�AA&ӿ��Y�m�_>r�atR��ؖ#s��+�Hڱmk�P�E;��A�k��SY�`���q�۷3���p�t�A��`��z����u��t�����p�����P�Y��`�'�.�����k�3x���75�Vd���+h�"��K��Xnn�'Q�\Cځ�!��W"�`Zt�dP��yqJ�����0����1��
rC��A��t!�?*l�=��g�	\M'��<��~���a����y�6�뾇Ή��duW\�Ҁ���N��Nׯ�˧��'� &�m�t_�T��},\ܛ(�kG�e�t�\���b���F���U3x;�W�|����9q���d���a�w���z�U&U�Ƨ/f"��1��i����?]fp�pK�*�ߘ;Qxm>},D��(TdaS��z�7B*�hF�}.%�/��J{!$�7j�?k+%�7��HR?���j��fO��qb�@U q	��C'�-C
���+zF,��W(5�W��m�
s��[�M��?�s�a(�3k�h""�w~��R�r1h@����7�Ч*�lcG�3ܜ�i�E���J��$��J���G�}x���'FQх���o���va�T����s�J�C@�rK�(��M9�aZH%A
�����B'Y�f��;��?�9i�������8�c'U�!��Ǚ�}�4�%�������1G37��;��&	g��<��A�xv��1�y �,����[w�������FĖ&��Z�X��b��Y���#O�K+�PX�X8�0'w�^�Hy\"��@�Nc����.�J��0�Z��&o���zq�耀�� ���y>x6Ű� ��5b%�ĭ����u�]�C��]���_{�W@��w]|̼"�ú���g	~��>Q����}��
x����t?�?J;�+�ļ)� �l�9��Fⱝ�إ�*��]��h�ߐ�,�Vo��ߦ�X�P��m}���}c����5u����	6q����O�(W��D6��/��h[vɽ$|�(�5�>�ú���r����.�������8c?물�a�y����\����6�\�D]���IC���nt ����Iċ��?kҹ^EC�L��u����b]�:,d���<�˭YW����2�]���T���Z��}iy�t���vi��Ҥp�(8*��c�X��%��@󔧍��D�)�G"7�'!QFb�,�:E��w1���t��]�I~�H�j��������ւ��+{�zj-9�)�w�_��v$�.Q��\Ke&qt0LY���J��P���i�FZ�W�o�aI֝���3��}�#𱣲':�ƻt���ac?�]�r��ʃH:&\fȱ�5�<�8_FF����ǱK��*0�����r�+"������@ر7Ɍm��{z��R�5�DKbPT�ޟǘ��`���,�=Z$���!d�����h��8��CtZSl+�[�"��.��C�p
T5���s������+ \Ʋ���h���v����v���@��syk����k�Z��h���I�j�>��[W�b����Ia�C�Ơ�x7��;���X�@��x���� 5nJW�=�9ӎ����w�xOd}���k0�\�gz����$/X�u׸�u!�/P�H��c$�����<��U��RAS��'d���o�S&�6�eJO�F��pf@mભѷ�!omup�/5h�33{4����Nװ��a&ÞIA���}�EM�-!"�^��<C�,�Zik�eҺVc�����:�	i��䵹��>=��������0Ia����GABǀ����b��|+<P�Y͞l�!E�D`�����/���CT����P��}^��4��K;S��GM$�E�v�k�t4j�w�RJ�!%3@r�/�Y`����zle>k��� ���i��@�ϝ8`]~k�cXY�m��G芢%|��m��j��[x꜁(���O�8�؍^F�Y�����! ��3y��B�a�* ?�a_��Mj����$��$r��aR������V5�l�I3�%6������.��ة�f�%�+�)����č�q�ǯ;g
�(���T	s�<O[;����@R�vdB�Ѩ���![�F��D�	!󈯪��F_wD��F�ja͚��v��i�p~E��?�r�%,��CL��W>R˼���{@e�#�g�Lx!�G��K��svI�{\^��ٷĒ��X�X�B.��H����F���N��P����Z)sG�"�.,����[�[R�ib���^��W�V�h N�/)�Xq����� ��Ks\)s�/3H��I��� ߳����s'8L��2� �:��(�]?��1�ǖ�-:� ��T ���<�k�cm�&�X�h��h��?��]U���Q�*=�Eb��}U��魗B�.`n�����C?��bx��6�| !�� W{�w�������1r�6��a��F�4�6��~���������m����G��&�S�ڑb��Y�?B�U\��کAx�w���5E9~��<�b!=�|z����e�ֆ��Ռ.�;���@/:m�1�g�s��9@Y��ۓ�k��@�C��P����ꔣ0������e���� |\���=�@T7��zv�\�o5����%O9z�*�S�yB$���C���ތ0T,m��j7}D_\ؽ�"���]-x�����9$�M�U�J�{dB���r��#"͒CfB߭�}V!�٫Ԝ!|JPZ�k��J�B�~3��-Y"�*k�Զ�z
�����[��I����L�/QW��hW�H3���Mx�͉F��@��~��s�٭)ȶ�ۡ}��:G��-C�Q������#�gIR�Ǻt�)\�Wm�ё��-�m���̙�tr'��bO�;�����c7U�A���e;������c�32:!����,[�8�����tc!	�S)"nz�oO��;:������LVj�[k���`����VB�������J��c�����٭�aJ�1խ��΁22N ���z��rcp��|0 ��?u6�5�>WB�!���VT���n�ΰz���3�t�����-�2��L�ҙ��獸�a�/qD�g��N��^�\.-b�������<��I�T��Ǿ}T�Ss�5��^���87�j�2���Y#N�<�%��-(;�;7����cW� o�@��S��U�mp���LV7��p���$o�r���q�P�	����K��?�@��*��@���ť2�*:w�h&�ԫ���l·�A�"�p�F���Gp,/��S����Vn<ph{eO�oF~���(^�F43��:�r9�lCcf��4A�toJ�5��t��z�Z��6���&e��/�}�p�<��[s	��̘�x�×���k8z�����
�\Q)��s�E6� �_�Sv�9���mvq��d,�
z��Ջf���Yh�Ǎ4�r���^jqh\�!�bm?Y�S�B*��5���2�&>�<5@���!�_U������R�!�:,�@I��<�g�]���_[#��<0L�E��U�Wg�t��)X�|�a8��	��ԯ椑S����l�Prp����vV]EP�P�u���?�eA6����l�ΐ���n�Vc�b��'?�x@*C;��Y��a�>\m�[��NO��Gm���xgS)�'-��W� �E*@���/�m�e����ۨ��u�P�����g�;9-`J�Q�\�!��vo�}Fz��X�^3��h�喿��)*���#m]��'D�e%��O�*$l�t������FLb���3�r�D&$(q�-|u�Z@<�o�>��5c��$���Q��E4�+\��,ɻ#�h���f)S<I+��γ9�FP�5��B�}-��pX�W��8�����f�^�6@U����t���<��n���F$H����@�-���j�2%��Z��5�{���h)c;?�v�)��杹_����}�u�I�1>��fkm�D�Z�A�=��H1���u?�<�jF��sL(X]���`W#<��A�s�*0�J��q���`��듃[LL����������*�0>�h��0!y)� IQ�j&jȋ�m�JˇHڃ�n=>6�U\�A3��L�D��������
����w�ɑ�ů���2��t�*���}As�;iZ�Tς�:�g$���秆��s3T�Ƈ�&gt��mDF7x�!��8/���Pv��V�0}mFtl�%+��TI��p�'��w��`��.?�)HU�&�OM��s���_�������6-z�l�PFO���\2�y~�<6�uPC�
:楀X�y����1i���,�U.���h�r�+���ˌX�w�3|��"WA��Y@gg%�RO�x��hUVVe�XJoTn�J%����R~��J\�/C�X��w�JB�hu���)A
I����k�m�/��Ɗ>sC��vS����y��D��i5T���J��z����"��KS��bu��&�꥘�F݊����z�E1��8VͶ���O��p9�o���2�������&���B��+`~nHK+�G�S��'���S<���2���k72|�@1��&̈_ ��f�U�A�Y����W�5�6R�S�q��K-\���D��[��\��Z@�t	����Ҁ+����t�S��8� ����( /�#��˞_v����
��!��i4�����I�����B�I����V9���J7!��@�:�*ޤ�<=]���f>$���ݝ�*`�1����Ji;V�h���a^�ҫ%M0=��3���"j_i��55���!A� �IU�S�p��Q����	�-���b���}�S������)�>����&�!�S�U�⨢I�Q��i��yj�S�B��C��T'���@�n�������\�!r+���G��U�������|��i��&�Hb���^'T���&��N�k�,:;�w�'_�}Eq/t�_i�p���:�̹7Z����p����D��̵Ύv
�%+�{��p���������$i#0?w�:�j�M�r}��oP�(�R��~��gv-Sƞ �8V�^h哱Q��b����0�$� ���.`���
��]·�* ��$E��ql�VZ#hڏ��G������$T��J��� ]�rC�%�L`��T�kA�&B�>�&ƧMC"C� "��u�~���x���!�����H�饟��4��Q$lr��+��e�Я���t!���:�F<L��Qbu�ێ�Y�xG���3H�f:fҴ̹�\��ᬷ%4s�`" ��ʣ:w��Ė梽��h
j4 �rE�2�֝��2ϑ�3�̾��JH�G(y��}�ݙ��Q�?*� ni���}6o�e$�6�ך]�- �c��ȋ�.ѱ��d��W�E:dx���@k����`�`��8	)���0��n�
c�) ����&i92��q�؎���G�{)��ŉq���pC�c��4��H�ن��&�+���:O���E��^�R��y��������D����҃�C:5R� "�����3�'�e@�g6�*�/M��X/j���y��u3
�N��Ĥn����K�6b�0����>��$�j�0��8�A��_����u���r/ie��_rT,�@���s�A�*f%�����6��)j�E_lkݫ	tX@�Ж���6Z�q�����[��^�I�O����&�h=@���o���z���=�g(eg���ld�I�^��!���Yߛ�E�W��t�	�,�-Q6�b�u�g���m��2�ʙ����*�.�]�Y25�A�W'satz�\5������	��*4�?��d4??�+��h�fM�]F��nF�3S΁�6˨��P�МaK�]��v����/I3Jq��n��j�20�R��������S���p<T���5+B�|���R�U�и����(y*Jl�h��K��!I���o	I�+�Ba5�����>�Uo��c@�Q�$/� uv��Ũ�V��s�H��ˢ|���׸>��=K4���V�)S��=a5�%A8�&��q��������q�'�:�1o&c���.�tIx�%0f�S�j=�b���q���4}3&�#��84ek�7.�w�<zi�n����T��Be��5��#^Z���ߣ����T�b���A)�ר�!S���mT�'�3��r�r��t���r��_+��R~\.�||d3�*a����Ti� �@a�#�/����ïҴ����;��3觠�&��gs� ��{|4e�=)�-�<���o����f,���)�%�!���ſcS���d-�d�q���s��#;���1)hS����ɖ=ku��aq4�.�,�S�| ��	W��O�&&�h\��I�O�Ǌ�m�׍U�	��
�=�I:��afd%gVѿ%����~�:�Z���6a���!0_OA�ydK�82*��c"�^_~$3Z=0����]0��,�g�����WG�S�K�A���G+���kC��B0M�$�P��n����Kz+�7I2�*%�~C
����J�$�h�}�a�6�0/�<PP�ԀRh&��Q޶(���_�]���V��-�+�`F!��!�#D�1���l5��.iV�1je$�ʇr��� �Q:�L���Y���y��I�>����=�ʚf�lr;�uJ���yNzu/�lQF+k�K�2G5q�ȓ��>Z�Y
�^�ѽ����P�RG��R�a-����7�fJ��S��G�D�r�h���3�c�Ɗ$���rt�Da-�"Y���H|�T��9ݼAC���չ��l����)�H2j�x�ȍS�x���T�:�n�����r>���#oȑF�#k�{��i\��l���L�x�Hy����}�j�2�/-�x��z�8�zc�H�$��̟��dvV�Q�ݟ�8� pHl�%K�}����qa%T�iAs�u���4[�`^�5]k��P�-����ND�����-��Y�M�	�Z���欒R�ZER�vܬ �a�H��r����e���������]���:Bj��n͆�^J�#1�}��Ԙ�>������5�m�9�Ԉu����G����'�$�ɟj��1sj��ZY���1_T�b�|��5� �R�z��?��'�B��<TU�i�^�T��sw۽��n���S���	ۇ[�,5�7^�ZRL,�k_��Cq㉎��:宿�@�Kh���R��&q!�Wz�W���y &9����u�
~��z1��L�e�6��'���P!��$��N�p���E�{[�z���C?_�g��C`q3�=��#�zy�ܦJB�3��O������[�AQ���;f��vv:�M��#!}H2j��"��.虘P���3a��mk�XS~�_�\4ʰ����CR�?!�(��`Jq�8�r���3�L&�W�G����Y� D;���&ԜC����=�A����.]I	���ӽ������0������mB�j8vD#�}j�&�J�-��{;�!�#��P�\S���&9�O  7�<m��e�6�j�B_�9��i�Gi�hF&�'��V8��!��
��_^7�9��J&��_�%�� -��,J��a�s%���sm�"�-)=�5��LbN��6�d����z�3��-8ۑ�K��wxS��r���'�=�a#I+w���R,�uD�ز���s�j�7u��f�ơ�\�5��QM���/���=���������{'�������3���#^�3.;w������G��'x+󞺯+M�s|*�^��:�����l��EUS�d@D�Ұ￠W�zC�$��ά��(|Q���\Cϥ@٘C+�����aT�6Ce~�����}˴+GȭWW�i�n���p7�N�\�ӝ���,�!q0N	2���
�C̃��v�g[L
�CA`�`T����oX,�%ܨB%�E�(o�n<����ν�T��`7�B��@QT��:cn�A6&�����f�����֒��LW�	�<sd�ȎDw\U�P���VɑC�DV�4��nk���	@�@��	���D���e}����%)UQ�ލ�<�?|�-�1Q�Q�������_���&xSʇL�S}�U���`[G�񆍡'1&�4�M!J���ˆ([�NdC�xm���n�����e�d}`xx��`,���k����ߒ�B.�ٺ���J�G�zvh�|�ʯd�Y��Md���$��f~���}c�<�Qw_�����#Fԭ=aG@��Ƶ*Ź���n]���x[
� х7����E��e'lI���v���~,zA���CG4�('��[�!�v ��}W3�Bqۧ(D���6��A�a��b�5X���C��+:*Zf��(��c;Io�6���Jq#n&���3��~DYӭ�~}3�'�G��gJ�f��AŶص��M���bN�2���{��%Z�b��E��DY��}ugn��$)�t���N�vV	8�~* ��ɮ�:�������f+�<x���F��e���4�k=Qzsgod��q߇u���Uh�.�5z!�H��9�d��1��gz�تђAJI�x���/�^F�$-�u@K3������
P	$K��-�h����������|�Ҋ�0)��\��g�XGC��Q�)&��<��g0�芜7�.3o�#���L�T��Y���W=8d��H]��[����4Q�n�*�2�nך�����℧.Wᶯ�o(��w�)zƑ�y#�y&�CS�1����uA�����x~E�"�U��b���������)2�Eh�%��kV��U2U���\��$[�g��;��S�9����s�\[�k�*�e�m��w=��x4���>���.�����fTgѶI)f7�x�ؠڞ�4�y�k��1���$�D,G$�z�F��-WD>8��������]Y�2U��d�o_�h�i�k����ϞFt��d�7RI���%�d�h\ׂf���9G[�՗��
���D�rk������b��� ��A������Oœ�}��<�������8�E7}���cʩ���Yl�Q�N:F�)���xy�*I��P����淶�I�s�EsB��ƚ|��F`=,������5Kr�:�wO�P]6@�D�{%�
|�H�J_R;y��;�C5�Z���C.<� �2�2���lt���R(����{-ox��E�x*�(�bK������~ Cգ���1@�z��L!������ZF����Qo�h�e��c�bt¼�Q&�YSiy�~#�D8&q��$>ɝ�Cϧ�m�x�����A�Ȭ�C)MB��jeԭ�</���mIs�#;�{���c�|�iyz%�O*4cV�>cc辁������#'$�-�Rjޓ�^���o@_�@�r�"����b�<�#E���=������e��);"��N��5\Ѕ i�5�SC#F��YſQ9R���i�0��M��z>�A@)��f�MlT�k�BrrXB0�+�|!�y��!��r�<�$�b��__�@t�5��}�ܜ��@�I���\�Hx�V�Wp����L/����������9�h���9'Έ�]�I�x�bzh�F�B{qͥM��7g���@�����L�꣈r6�T`�Z� -�_�}w@��2�6s��W&�G:]�Ϋ��8r(�i�X�f�dZ�a����f'~�ɱ��V����ŶC�	k%b�K@��W�o�R�~��a����Ҧ�޸�țl�!r_�������Xϓ�>���kp���P�5�0���`d';��=nb���|:{�U���!Y�LӅ�٣c�8�c%R��[~x�2���1��/@�n�4�����"�S.!��/�
�O��I�y�[��}=����$�K�z���Onr<���<��p�i��X�� ?�X���׽I��}��@�П�{R��-���
��B+[��1���y�͜>���uW3_����f������='��ţ� �2��`YO����J�P4�����쇪d�C��M����n%��ŏ4�rs�[�3G/�-;/..����N8&q�R��m �#y ��0�0�n����R��M�6I�Sd�z<~��0RU���w��<��Ġ�u�u$}�3��+--��/��0�F�E�ϼ�O�g)b&�w�x�B���8w�s]��։��``,h��d�8cvj$����n���*�>��O�*E���喭Q�D�����たn��t�ھ����\X���,-�L�]5j��LзV�}�`_�_�q'�槕��b�G�3���cA�dm�)�\��F�2K�r"�R���m!�xA	�/�pHё?p�)e��®�����hTgmlI���}�c��`���k}^CU��h��hG�͐�y�T�w�;���׎�UB��[�4
��1 �,vj������-��(t5�!���Z��^%��~z�w�A�1�S+wS�������8�0-���O�x��6J�8��n],0�]������<0�9�d��+Ɖp������_����\�-���$R�O��O��v��P�2��J�W�S�W�ؼȺx(���uE!]���0d :ͻ��x� �@�6��a��҄�wZ(]ѻ����$	ȴw��	Q�*cC%yy��	�DkE����֖�ԋff���~D���-y|7�w�8p�Y,j,�O���˭�S!��k=�)�@�gㅭ3��y��łd��7�~�Ąj�Y$f�wo���Ī8EtB��6fk��µ(�a=�VQ�Z�cb?#� aaB��K&��nLX�J�D�^L�N��֒ؙ�� (�Z�^�|@�};6�$�~&���R�S���]k:�Y�ၭ|�H��=�(�^:r�%��e�(k)�6������d��<�5_uvqT��P:A�f�#��#� ��|*9`���W�z���8�8ݕ&�@0�&�&O�c�l��V�iA��ݤ
�Ё�aq]���}8��áI՘Ru�.~F��Cd|O�Q/藌� �_�\�`� �'&�8lȘ�'����5����g�3e��ǛL�5��1:[�=˴���ǜt�At���/�������mR;��γ�,�ov/P�{���sK!{��k�A>�딆�)� D��IC gs���OA��Γ�P3�1���w�:	,=��y`�G{"No�K�pDJ�PU�hIE=d��hU������tt?�/,=�:Ҏ�c�.���+Q�hG��1g��kw%
u�o:%���t���7?�K��lmؓ�����X?��c�Y��A�`m�Les��)gt�%k�z
P�^��|�U�,�k��<tdd�#�Y��E��nUA�@���=�������L��A�FsQ�ķ'�(Y����=�G^i��!4�F�v�T����L�a�O�+�;ԭXĘPU�w�{t��õ����ɕ�[SLiE�|7�)���R�O��N3�kkr��N�#�;#ԦͽD���M�س�����k�^I\u�K�P�΃+2uPG*��R��߳���A]��]�ꡢU�Fu��M�@��w���09V�Ѻd�D2Y��X4_�x'��N��n�%DT�����oۋHA��?t.�.�t˷��<�E4$;�p��.zCw-����X��׷��9(��������H�p��"]��%MȖ���gt��c�%���l���A]�sh�?�6�����%3�ac����
�zȉ�L&�Au!�P��VMF��k��n-�e\׏f^��L�Zk����-�G��N2�t\K�B	�4�34C����;�-���@� ��$��l��I%w�>��'#��Y��K�oۋ;.Q������@�e2~D2�������<��#b*����*��>'kw%�0V�:�4�*�`�m-�j? ���
�r�~-t$�5���p�I����e���-J`����׮�t��S�9��;�}�KgZ"��m�:H�=-T0֮@��;�ljC�=���H!zSXgJr!��p�U��
����k�5T"�8�_��A��\�E!'*��7u�c�$�RS�\��|;/�6�'�>�!R2׳��K���D�n6�pI	&~����7^���\k)�<�8�7�7z���v��(N8�$����	�(�D��`:ħ��;�Y{�@Z�>�%�3�U���P��o+5�3�������i�0��} Y�*�x��2ݢ�+ݳ^��=*V%=�#o(�SM�Ń�Wڸf;���צ6�T+�.��@G}6��J\D���-C�_&���r��!��EU����v�Q�q#�����X[��q�M]��W�{$���~�" ���7��:���'ܰ�\!�K,N�4�'8]C$���N␐��G?��0��^;��[��{G��ߑ��<��"_�V��� ��j|_g�]�x��|���-*3�N4G�}�U�����٣\�;\��N�f2�4�K�u+/��̭<NIj��%3�K�-*dզ���̢�W�T-�T�c���&�ev��+oϕ�CO��n��12i�Sdۻ�u��0�;�F|�v�q5�f�"�%�G}詟��ة~/_ %��m���'�X����[��t����S�\A~��`m��B8 �\Μ_�Ȗ㾎���©U+���������Q�a�<q�_1<d�L�k�����Oc*��'��4j��.`����?0@_	���-xЖ�j�U�SC�o�S�dz,<�Շ�In��R���c�{ڶ�:v�D��K�M�h��M��!(��;����v��H��ē���#.��g�}���k�BK���X.mҺ$(��������w;^㷴����}��U<� p4�<��������B4��Q>��g���1Q;#��X�Z"5�KdO��E� b�c9T��VE+&�j��}3��M]�|�m�X����b�7)h��W�v�N|�t����w,�|8A���G?|�c�_�b-,���)�S�C��Iw/2�r� %�� &�?����>�W�;x|����1�Rl���0�����wm LO1��6���K�g�h)�� ��&�r����f�Le�tp^#>����d#����v�vّ߄���z�:�x=!�Gaw��x��;������F�4:/}>P>�zZY,�d�-~WX	峚e��7��!8�x��x��
3�0,LVV�@��b�Q^q�;ɜ(BɆ����Dl��=ʞ&�y��,���x�1 D#�ܛ¥�tb]Lm�:��YO�o>8�B�8�,Vm�?<4Aƞ��Yh<�-���)X��G|r���,U�-4�H�u��u�=��j8�e��[���;	.� �w�dv���Ɋ^�ĔK5���3R���B?����/�/*�����~	a�|���aa�8�fgz�ߩ���K�t^Z =��7��(�S7f��0�TP[X���Ic�\v��7�(`�_������{$EQ���X��_<���.c �|�Z���&��Q���c��ۨ�� ���0ӍC�y"^b��ux��88�W&܂Udr�
����40-�y"A�=�~��յ�/lcxҙA�׸R�Z�o"S_�C)��Y��7H���4��GOͫ��8���a�cSG�nc�����%͊V���9J�[�����"���=�1%	q��K˙��	��h"q��x�#V���w�8�91 7��Ѷ���d�Dz�G�pY��d��H���.Șq)}#^������Ĵ�|��\��?�5�U�a�̣֠k5#E��}��JJ�f�$�o�P��0h�
��*��&��W�JIo�~0�c�9(D(߼3�*z9�=
��� �r�%��ru���%�M�bo��>&�ȃ<�S��~�a �X������;bpb��K�Yo�O�\�l��2*r�%��!&�¬sf/�m,�s���E�i�][�k��5rޡ�y	܃2Y��XB��_�! �'��qz�fn�$nhN$�G�M��Z��b\U�?�kpn�⠹HV��I���\1�Fie�g!�FסE����_9t&a�I�i������5����d���h�_H؉�/�jwfVH��[erǧ]<n�^�6��HQ7�j�'|@' �����b�-!x�C򃎤��]�.Z�,�[Y�)n�]��'*<d X��ՀV6n&?����)�������v�`���&�B�Hmi��[d7M�3�`_����߮.��Y}����At��e��t=`@P?s�coku
�l���Ql�k&�D|g�G#�M�i�A^u@r:�R-�G�aK��R_���y�Fyq�.�����A���l�T̾���s��;9�h�B��9���Gl���4|�kH��X*=�l�V~���4��^�oEe����=yٿh�f��[�#��zʖ��ߜ��ƴ����_�L�`ћn��K�o���Q)�ڭX�o]T�(��AK�'�k]�s��v12q��X�\0=���mw�Y`�X�3q����+�k��BR0�8���s
�1)U�c�mC�+ QQ!�g�G3S5�ސ W�V����B����A��zDU��<F\@�-�Z��5������W����v�LsZâ�Py�|��v��ɛ2tN�.���2����l�$��GU�1�#�`�4��]e	��E�A|u���:;%I^~hN+��u�����iB�x���->r������}��+V� lq�e���z��#��O��ë���mK�uc�S�ח3F`5��.h{���D��K�y����rygM6�Zև��7��4���䫀�*�)��%Q����y/�o�zh�ߠ�v����1����9)Dj�s�{<��`��x�2�e0���*����_®����>�j�P���#r�#�]c+�V"o]�͐���R��9ڮ�O���fg�A2廒b�9��"���(:�di�R�tp�M$�<HU���RԒ!RYrKݠ�G-k#F)<�ڄod.��圪6�ُ�gF���-�-#_�ō�#���VJ��UbߵQ���H�&���h���2��	W��2l���1�m�1{}'�����b�>��$��C��B6�A��k�8�.k�Yâ*DJ�$�wxv0��TŒ<���|u|.���/塾.��]�x�^�� S�
��ϫ=�(g"�_����r�>P{�)U��d=>�N��;���R�Kʊʊ|�8�����q��=�0,˦��߉��a%D�t���B��З!s0��.7F*�=Z��?��*��*��&��q�Աі�Eid�2`	����2$�2������6��Lr�'��\��% �N���M�Y��Z.Z݀UaP��I����~!���e�ґ�\�C�:�oM}���)ߗ��M34'
	Q:(�?x?|�B4���n/ ����Yb&�9\�c�G�X�d{�v���W�U�����rK��:�o�ۅ�c�B2@�e�ʬpZ�Sz��,���]��2G2V:�.W���"��y����?���u�s��/�`'� �j	����#u���
��h�=N��K�4��ס*�9��I
d+����mW �A��6T�I���z&c��qg��^��Ӧ1��h��`�����hU�)�yh�ӎ;)^	&��^O���zg�9�TV��Ƿ�Sgt>��c���+mI�?fb͸/�)\�[��	��Ը�/��>v9g���86� D.T�?(�*"pf����]l�5� kA[�^�<֍�렌+�po��趾+�:� k�?gQ��2��-�i��Npq�#a�c�1�$�7['��ާF��N�=cL$e�cy[H��~;����J���#�żCX�3*�Ն��Շ���e�\Ra�,:���{.Nĵ���u�f�s07���p�� �BWr���S��#��:�4���� [38SQ��B�v-6�Ͻ��U
I|3�C=��6S���c�@-Ѐ�Xmr���
����RO��JUW�|KxJw�LW�~ihΠ_���n�`��m���� 
0��Ɨb�4�"��ɫjGp*�2H��*�I˅.9fN��8T�X����%YH�`9�T+�����Tڷ���j�P��E���E�pq_�xs5�ε�t�OU8#����6��n`��	�O�֏��o�p��E�<8����|gVM�$Q��~u���e�TƲ�6k=��J��ԉ'2f&)�gGU����I{���b�yCg�D�ji���2�����Mג{�:��,�*�'�7�+do΂�n�̗in!|̢��-��kͨ�+��,�		��ɾ�ܐB��HbW�k�P�46����"_6;3��S(V[���p�d�3������1ɇ�b<��f2j�:ҙ�OF7��o��4��� 䶌�5Pc'��k���9�/���%ZU���a�}�%b	��Vʹ|��?Z��L�CWU�=`�Fr\�^�kƙo�=螈��"�J����+ȇcN"�3��XA��[����)���a�ZŦn�����@�O�P�/(+��h���'�,v��j������D �ѻ"�>S�q�x�
��#`���`�k�[�l6��'�u�"��W��j�zC/�=�=)C&����$���y2�z��5
lQ���P�z����l��KJ���
���b�og��T�R�����a��6D���}^y���q����4��5 ?��͹������Z��E�*�Y(�E��@�� �િT�3ަnYR�z-z6�i����)��W�Z�m{y��KH�UbNnc�IN�.��6�˩&t@095l�M�$��#s��i��x$w�TBy�Sɬť����k�q�)�ȅ	��s�T^CT�����d��:���%q�4K']m$W�2���;R��C9w�{?�y����!kI��VG,�5�kz2da��i��5�U�Ob[� �Ik�
�d>�
��E��z=��~<�\���$��� 1)qrY�	;2��n{���Ck�&϶y�x�f�����_bϵ�xZ�Y���<%j����1A�#�a��i4רf�^6�/���?5�0VG7�������a
)ϭtZ2�wJa+���iWeC���9QD^�/yl��P�t����ӹk�������#�e
8s'PI�������pjzP�ޘ\���9h�RV�'�Q�����S�A��vң���~�奩�KM)0�� 3w��ZFq'D�ӧ�p�n.!1���Mε-����Mo��l������B3/���c��ǹ���J��?�,�j���L��)�&��-y�91�b�	]�s-<\��5C�xk3��oH�PE�֬!a�/�mܭ�_x�>[Y��wիNB�e:��b$��W6å�����7��6�Ǔ#��2�)3Tk��m]�J"��hz�M��>��>�u�����ڗ�����f=����"/%�8x�9��Hs��}�%do�3�B��#��hj^Q3��ά�[r����$%��1���q����^�� �E��w�G�*tg�N���z lnŭ/^�<w��͖��4��	�:��=@�!��m��em��ڨq[�G=SJ>Cv��NX�A��u��{kq_�t�X;LR�O �uk}x[��I��M��tc���Z�q����
�QEG4��6����W��E�d�Bʧ��5��)hx�?3i oP���Z�,``��rj��k���L�i}�e��(ۛ���>�ϴ�;��I�PP�(<����լ�W>(ԃK=�������޵��*��ȁG.�aYךT/8�u���9���.�<h��.!��D�k��`W��w�����_����K,~���ؤ�%1�6D�A�S�72SV O9�������cVᄜ��������8)��3�&�W&�If{#W�i��]��d���6o��X�͚�@_Q�������NG�Zb����}?�`爭�=�oƮFğ~#)��Ҽ�I#յ#�Y��	n@ꞹ�戶	�3h'[�Gty�bKX��Xkf�e@v���*�PT��F|h�v��%��L6��O�G��/�`?��)rOy'd�e|�ʙC5I�)��Ȑ�P����\�멽ޮ��cODSK��Pu��C/c���2@>��_�����8��yt�U������=�4Īeſ�Y�������z�f*�p��XU�<,�\vw�\�@�wD7^7;T��f�������x��:��LL���D $+ъAZԉ����֊�)�V�'f��_#��=o	ji���CuwFz�� ���y�e%]��U�>��Լ�o^���׉k��ES������T�:s
S(a�֔�ׯ�X�xY���IO�[�D �5����¤�Vo +�W����Ė�s_�����z�Y�ne�S��u[����g�s�R~�!'�j�7����Z,>��>�)�fotˠ0h�ca3M`��+be�m�a|��ƒ{k�F�bۘn��J֙�|~U҅�b������e���T��<8��ɒ}��ጌ�m������"�]Hd��`6�"!8@��x����gIf�)H���OGO)8���͟�rT-%1�(xS���%/ǘ�UA����5/3JPzf��i3���ƌ�n�|k��)^��lG��w �;O����a��P�iZX��Ys�Oc��9S@]2���v� ���tj)iB���x�L�^\0���z^�y[B� vԁ}hE��-@�zaG|�Zj���̢eʬ�nE��m�N�
� Y��Nq����h:M%�>h�v���� ��A����!+��y�e0��W��*���K9��Av��8�w�4��9r݇��p̯�%��¼�#�c������ڱ5����iߣU͸6�������&~wŦ�?>g�P� ��䢿�M���C�\�q�Q/�����)����@:׉R�}"�nZ7�<-Pj6��:���k������ǀ-LRr��Q�� i⸅�"B('�(Ow�&��<I(�#�Z�����wƈ�M�e���hдߊ�}*��Y��~-)B{���s�KhY��-PoF����~D���Ő)�o��_�0*�����nlcv��h7 .�"� �ۘE����f'ox;�'������OV�eBS�B~VA��О�7˽�uUY�Θb�~�Θ !6"P�4������a���A6R��t�L�%���Uf_~6�D�`=b��pt!��<Y�J�+��2�����P�GZQ�(X�[��*-�l?~4������g=+��Cƿ:��ڟ�q8{c(=l)���b�������Ns�p�iR�hB���N[��#ɱ93��a�r˼#3ZI9�F	ڶ뵃�ׄ6��3���� ~fV9�T]���������
t�qn�h>��]+�lg^��}!�"�q� 1��`PIF��ʷ��m�gG�bM�*�k$�v�/?�*�I�D�UԱҞ2UN�P�I/�U ;k��qF�[-��5�K̴2/S�j�.�ro�,��WR�'��H5#9����X'��ָ݊#�<���/<�B�R_�b���'L������C�vg�T�Y��(+%rǀ69���(��Y�Ղ,�љU�x�ȑ/Ʉ�4�<���1"��%��2��ԙf�0����
�NU-�,
[��v]m�
�Ꮮ��Up�rPN���a��d�뇠�
n#ZD�#8#g8tX_�\�ױ_p�`�eL]��k�[1���{z�r��J��/Qx�kH�
܁�z��_��m��5!�V��7�7@�Í������-x�|T��	2�.c�`ף"��-+�#��'aP��H~�?�&�ʁ:�cl|�E��ѺU�fo���n�X�q��&_�����u,��dQ{���C���z���<�p�2D�Ş�\���cL��&���13�������&)�����Y�w~���Xa��ﭒ�㡳�ip=N�R�&�nC5��1Q.�K�����Њ�$0����>�Xэ;��(Z��0�H[���6,�:���Q/V@w�����Lɟ��%ָ�AB+(FZ��|M����O�]G�`���ε}�t����z��n?|p���/���ͩ�Hi�$9��<A[�Ш�2t%D8\yYѪ��r)5��/Jd�na�u �� D�=�v	�� c�yv��'��".C:F��!HϹu՘e�� ��Z� �:`fU�ݺ*��ݣ��K3��"O+�L�p� ,3Ӵp��{���n���J^]�C��-7O(C�i�]��#�O1`yf�3�*�]	�����&h���Si�<ctw�6��6sR�)������4���$����=�vs�զ����u?���ɑ�*`�yF%�L7�����M}}/8�����GG���-H�L���_��%γz�O@��lOj�e -:�LE�3ѓ���{�F���4-�u���k�X��<��*�gκ�ۄ�d��2Wr�j� f|�[�_<ݪ�,��="A���Ł47�����[�'��g��s�eJ��U��l)�5�.
�%�����8跿��8��_�:��D�%�p;#%m g���o�_�Ѷ3�O��F}{���E� ��%��
﯄#��s�o���P.�����5�8�u�@�-�<�4�{���1�/q�W~���a��|,o'�h: 1�X��*���D}��9�Nc���	���+U�pp�� RP9k��r���豎�ā�)��n���ۈ��Gf4�����j���z\�f�:���VP��[k�\ׅ�A8�HHF�@٢�<�D��n�ۛ�4��x���c���Qi{t���Q��\��س�	�B��E��왶��Lu��@+�i�织~.��IIMtr#�sæ�p����ي��d�S��<eY���m^u�`���&Z`i�����'�F�0��%_����kD�dK?���m}D�fq�I#�s��i6
�G �a�y�wb��:G ���iw_�)�@��$�W��%��K��%�]�5�����2�V悚/�5M �����8A�%c}АF���t�!�-c��\��rSɨ���r$���.[P�H��R]�j^T��p��`q���S�@�h�@q�K���@�~}�����WW��ӷn{3A	t�#g�d/��B_x��}�aDW��;�*N�cAX�(�Av0�%L?;2��h4���0?�m (��v�Aw��9�����KA�+k�� N�f�[�^�[G���-;�3�@m�kH�Y&�/�� ���U�i��/j��W*	0�v��h��T���V7���-HÖ�H�n4�s�7�쎌"�6k~�8X�h	_�Z]$ ��+�%B��Ĝ5<d�%����X�Y��@�U�����S���nz'�M�M��ǿ�D�3v��,/�A����Ӕ5;3���_|��*tn�H�Ht̅�)��]BP�MK�S3L�־;��iD�q�e��yp6Uː���{f�`��L��v��T�$;���	�5�]�D|o�r#�|1Ͼ�V4/�fg��"��S��i�*�b,y��mK��ϥ���iF��x_N�#�PC���`���q�#j��`0h�B�Ζ�;R�v%�0;&s�:�|b-
�.єG��Q�<��ё �Y��:����X� L�ЎN����m��cE�PȅEeX�A�U�=��ޜ��V2�K���H'����āJ��Q���Ƨ~�Þ��.�����'g?��r�{��>��$P>��䢙C���Г?� ����b������5�sу�+<���l���!��*��dvE�k��~� �L`��r�0�\�6qrB���.�Z��q��(ݭDQ\����@�+�� ���T[�~���u�/X8��"?�a)9L�(����� J�4k�8�mW��F��(�Y"2F�N�IOG�-�E�Mh�������^��~�3	��`h��/u��ext�ғ�d��4�\+ ��ʒ��q��t$���	� X;N}��  �|Ϟ(MI��ǧ����)\LUr"gO���F��֧٬�
�H������X�d�l��l�������%p�80��uM��y5J� ��^c��ю��.�VѨZ����\�$K�8���R5���˂u�ܲ���t��]���~>��,�F,B�ƅ�0aSy�Aisw�[Ul�!d�����
WB�?)�&�N��O��z*k��l���ϋ�z\�b[��1\ � )>�W��h�L�$�446>:u�͙�Ü+�B-��	�����X�V���/M�{�.�8R��;���4˔���ZOm�h�`����1Kt�J5���Ǒ{��㌦U7Û���� ^��BtWQ�D�����WJ'^D��ȴ��u���Y?�	\d��{�5v�t	��*����50���8��Պ�@씲��@��DPˠ��B�?`������U"~ѳ�'y1���"�]ZiI�� e�a�﵃SǕ�m�z=��;B,/aY�[xD3X�T�6�#W��m��,V�6��W���p��'� �U�pZ}.�c-٭�|7���'�Q@�`��6K���H������/���,jo��{A����m��ʦ�`��n�-��R�q]_�#b����/�Ͽ#;t��U{ �|��'��+������Hh25/RD����$�m4���<?�ة�'¢G�ῒSL{	���~ M�}�` �^%8v	����q��oԤ,�(W,��y�U���}�5�{�v(��L�Z6;sM�;���}Ũ�5�;v�8m�6���lU�J>�B	E��Pi �F���:�TK(���h�=Y��x�s��6�q���-X��rMLC	�ߛe�`0v�i[c��̣&���]�B�p���1�3�k%2P��l�����S�s{�l���m�=O�$'���I3���ȓy����
l�%(�i[������U�_���eů��f���q���mc|ߣT��p��̺2?@a#�މ�2�A��^��j�NI� |9�+u ��_���`���R.�dY�k���3�8»�� �Lf���UHle�o���L�۱T����"�]De����_�$^W�@f+�e�ꗏ�fl6>���BW�� u<ĎC���R9#�������5�ё+ئ�<���!|@�1��P1����|^a�P��a���O�J�l	C�w���ط4�!�F^r�y��xA��R.���$fw�$��W�kW�
��8�z����Qi�B�"}�7qSOp�nm���q�>�:d��z���--(���g(h���+�]g��W��&�}�$�e��]�X�,�xL[m�d�ܥEm��c���PV�e��59ǭZQq�]2T`�l$�����L}O>�������#a�
z3I��Lp��X�/o����w���u捞t�N�{���6���e+�����N���>�M��˥�^�Ő������/x��4���%gVl2���[J�~�C��!p!�� O�w{�1�ڽ=�p�1X<�3���#*�����<k<����U��G	����$$j��̳E���Z��a�z[��}K��Z������%����QI��L��y��q|�g����A�a�2��.,gM�V0�n�E.��0%Pp���~T�u��z��h2��� O���
U�.���A�1�?��/�bㄸx�#9����^��aPnI�d�c�2-����K�3eA+`8�׹�E��'Y6�k���lA2��϶��X�9/�:�v��!3���Yo~K�$�+)�k�ó�
��W��Ҝ)���!e��Oj���&�?g�9��q�N�կʚӃ 2�}%3S�J�U��V}���s�g"�Z�j���0��M�*$��C��v�yIi�5���~�[�D��AZ���!�$�c�)׈�-2��}�T�3Q<�y��`����Y'G��1x�g.B���D�����`L l��&Rߛ3d�ʕ�;��9�?R��2����uJ�Y�f��4�l�26^-(g�Y�F}��.����,�V
�b:��g)J���Cy�`�N�F�y�9������7�G�c����"�[�A�������O)fz5�������G���x_���X5�Zߨ0�G-���q�]6�]�*ԩ���ۢ��j�4������&�&.�FϤV{�-,��'yr�˜<�O��)In�ZEA�`���-K�}�6�������\��z�7��nW>Dg6=��s�#���$�A����v>Y\�όS�X�ܺ�Xrc]/�����q�o`���D��:�Ud�y�?e���l$��>��ɹ2T<dV��F&x���]O	�""����p��Wk�n����ż�t�"*(.p
�"!T��tQ�v��j�=|�c��a�>b�@e���z���&���{	�ŖJW����&������(�{��V]�ګl�~�P�B�>%I��T�$�y-\%T�u��c^=]�ڛlM�P޹�M��ƪ����Z1r4� ��mpA���{���'��s�E��nIS1	-[S&��o�m��v��_9#�.�B�����<�	�^�r\�*Q�W�C���D�V�趌����|�J+�S�����;����`rN.��(�/NX!YF	�ݰ�o�w���e���Y�&��h����C��JY�� �"��g~���/��k\B�$X�	���_a�U`Bo|�ܘ6f���MYG��^ �J5cd���>}��ngB�4�nWK�#J��ҭi7���׉��C\�6ݵp8꜂�o=\�������k���{%���+�&��u�v�4�����)�nSKaT����fV��G�/�2�2�h��HW�=�ZX������^��ȵ�Ln�"w��Ӻ�f�}�_�r@>�h�ay�-淔�_{���p��^��A��ʯ�����ݜ�u���o jL��P��c+�`�T(���꟪qѨT}f���N�����!KyOkiJM�Β�a���>ݩ|s.r
�؇�l��O!�cRi$	pltN��/��Ӎ��s�.�Qτ�\��Z0�<��>�,1��ʄ簬g�쐧f,�#�8�S|�������ږw,��	�3d�y�궫�S���8���<��"n�d~�s�p�9���ÀZ]�{Ϧěx�f���Qի�~bb���pT:�Y��m�ہ�\`DR�Z���9�c��\�Z��+x;4�әm[�g�Z������1TeR����jH��g�1n�Ze(�s�}g,vH�|�x/ܻܓU=4Z�p�����!�7��Q��,� ����Ϭ��!?\��DTI/cCѷ%����@���.H���ȇ���S6AC.�1���xC�D\U�P�����8*D�[}��ɻq�ڂ�b#��)g	fq��G�����lu��6bܔ��f=F�����&�F����Ϥ �n�N��黾R.���D�1���_H�xG��:���ٶo��bJ�|�r W k��jK�{X��ޡq}��J���������:=��!��~Z���Õ��U��m��Ǖ��UGn%Ƈ��9�"��̸��v�P��a��A06m�,Q��/�U|�}~�1�!�&�c��[Ȃ����@0�,�aA!u&��arl��f0���/F�/�:
����u��k��<Ohn%&[�R�"z���̎v\u_[C�����ΐ[]�L@��X�	����ڞ�T"U	Jv���������v��c#�K鼗Ac~������>��Atry8)�Ò-8�^ͷ��_5�s�w��zF�+���9��%�̿m�V�,AO�:R5G��c�gB�!.�*�b�폖��UO��>��yWB��٠}�Ay��03G�������ʤ|�iz�)V���f}�x�_�������	�E��Hڦܭ#�v~�,#r�C�q){�l����6�3�z�;-:��3�	��Fe�m�~�U��߉%��ַ.D��-V��@������r�UiU�N�	7A rNS{�0M�����6�@���}���X<�R�|�Jq��E�w�7ۇ��ޡS�r����� �=u2X�L\j�sdU���2"��g2W����<���8(`��S���D�4C8e}�&��.wD�o�C8q���80ߩ	܉���c@����ǛҖ@J�n��SU��Z����� ���-֙�#�ʭ/��G�\v��-�.17������V�ģ	8�-J������=����o����	�->��z���#Cf���k���A�0̶���f����&թ[հ�&XG�
+�|_ޯ��2Ř��rA�Geü>�$�K��?� o��:CX�O�A�]�2��(�=��T`�~x��W�
��3�]n�bضr\�=Ͷw�ؽ�������qY���#W��D��;���!�rG\O�i$`]�'�ڍ5��G�+�:v��G�Hj���f�@u���j���X���v��n�}>B{yx�r� �w��I�E�;���Dn=1�u�03� ��H�.P� ��c�8�q6P- ������S�!MO�t/��\ȇ���CMx5EP4[D���X�ö#�&!wL[O�� e����|��u��о�p
���O�j�9;f���{���������hu�űi���0l9a��;���Z�(���W����[,S2�6���R.�WhN��C����?�F���1C�����3����z$��d7Q.О���?����_�4��_��A�\u\��o|�c�,��ҟ��@�Dcu���/�d-!ni�ГX�7��)�� x�&a�4 Y;oC�j�Z�8�y���0�+����srL��,��¦�ѕ��9ҭ�e�>�_ �e]����]���7�l���^�FǄ=�����twЬ�L&�k�#��s(,��������l����c!�M���+$�Z�P�H�N�����b?%������{���N6�}'Ab��Lf�WϮ̈́=-�0qO��f�4<��ھȧYm����=����TE�ī&�w!� u�@�S���j�uW[L��xXS�2P��a�/s����3߸$��l*/ؠ�]�<<�� xf���o(4ݝz؝.�qG�S��1�(��v��X��������7���+�V�h�:��sU�$c�H&$��9��������� e/�P��M�ܵ���Q��(�fb�2�I^{��D��
-ᬊ������|F�Y�Z�j\�$0�|zgD+��?�DE��o˂9:�|t���HdQ�ƇU�;���<c>z	�6:X��+-u\��O�?�d�`c��v�,��h�;�Q�UIw
zcp�[��	ObBrl�,l�֜�J�YpuT�"��T���Y��;�@�ձ`�`�!U��X�B�?��]2�&z��y5��m8jL?iѾ�b~���V�ي�`�/�X(7AB���j�_�z�ܮ�r���ԅ�B.�O!��Zo����~�E��w�]WY�)�p�^�������{*���)�P�JHb�P���E'k$�����^�b��C]�t-�~_��)!^��Bz�s�;�]�^�h8zt��1L	���e�G�'��ͣ?�m�.&L�q���x܊��pd#�+V_$�]=�g�������m;͆�ޯ�η��3L2DA�ѣ��_d���Y��x�8�
Z���@³�q�~� _��F����Φe+�0��=�����R��Zw驢��?�׉p]�ʭaCG��2�hZ��N�חpCx��� ��}��"8��J FMc�B�$�!�s�н�U-]�K��t�£$M���?RN�rk������GI����D-���yd�%����`L�E�c������9�A˽ü�^�HHL�m��İ`�HGǅ��%u�������#�����o.KF0���v�	��u 6�>�&zӑ��fTI�J&+�I� �~j��Lz�u~g���H*���a�8 Y3|5�wAr�M�>����g�؎�pNݾ����@��G[��0�o ��]�
�Vj������N��L
�u⬩�Y���4n�ɒ�5���a��dY��K�\ՙf��Q	�`�f�,&K��y��w~�Q�_Æj�RuԹ��8M_V�̖��t'#��ha��!;B:�I��F3��n�@`�D3�w�l"D�v���Q��JR�Ak	w;��S)?�;�p>�sc��Cm������É�n � ��
��\,���'��y�1��a{�ʛ&1|)v$f/�,��zU��7Jg�j�P�zZ����xr�b�d���q�I:ŭ�>?ݶq�Wd~���K��[Lko���M�,�G��Y��P`_�!*� ��5�&�6�ݢ�z�8�p��u�8!f������~6�-����Ӿ�rsC�D��:�\VO��tt��
�I� ��s���Cj��P��6�Ȱ~�#�u}���&�b���6�?D�9�U�P�1hd��F*�;��5�n��E@Cm�nA���IHf@AW��c���܎`�E
�Y�.��!vZI��4��0jL�)=��&�������UFn�)W��g&h<!IEٵ���
)N�7�e�4��2iFeۉ��ϛ�/Ć�t�ٺ}ҳ�ާ��J"��$�������p|V���VtTn���8b�>7-����L��0)�D����զ�z��5fޢU�X���_}2|1�u�����Y)@��|�Ÿ�M4ʐ���Nk9��`^*���J$Uw��ӏ%ө��z-�.�����_5ڠ� cʁ��8��Ij}aP7�G����W�Tfn'"�z<޲v"	t��a|5����bti5x��k`g���d�Ag�S(��`��#�L��#�3��k^oH�d�.r��CUǕ�xv�*q��[ay�r%5S�i^�X�'b�=񷆑IŇ7F�1N�AH���-C��&����P�9G�����m�(�gЯv�	Bx�	�yÖ\��.`J�|q�;W�qH�"F�I�����	�p)��ԯĶ��yq<l���{�l���jm�G��a*�s}�*C�=�`o�	M0�Z���)OMU�_�Bud��{yBWQu�o�>[W�h�K�:ATjx{N��DwK�)oФ���Sn��E�R�Q)Y֤��!'*�i�6~�J�U-��l�.���7��SnP���}����yQ�`���O�����(;ňM/�cM߭�-��3/}*քF�i\�m��Րo sE�w{X�}�j�7�_2�KDg��Xœ�f��mz��N�47Z�g��O.��#���l~�6�~��8�S;4hp��X��X@K���c���}��֔P�1�mװ��gW{�M�Dk��!6k}��r��w��y"Ǯ���MaDZ��N���?�p�%�A���hx5
�@���L�g��i�<\�2�0���M��:_�r."�W+���>>K��^�t@K��"�"!"���E���|��f��5����L��W���k��h�ʣ�f�@�K�CLɠ�=�V(�~N~��ˍ��Z��0���iI����JԖh�^��헗꾡Zd$K���f�g�[�6��H���> �L� �U�_&ʬ�vV�{���.���
��;��jV�Ql*�U�k)a�aw<��ˉ���|��$�	�@��Ҍ�(ή�����|F�9�3�ҭ	{��B}�`/��Yd��k2l'�����t���9�>-�!�B���Hj���%lP���F[���E�Hp�e�/D�Ʀߥ��(Q�K��7���60Ԃf�ؼq�=v*���6�<�ݼ���v���Js��G)��?n��4L�x�y{��u#��v�el��1�[�D
�H�m�ҡ*r
��VS�92'��;Lq+�9�3QCQ��O��(�B@�
��,��*�c~Ӈ��Gbؘk�����Z�G�R!���q�t�6��e�5yIQϸ�-Q+��&��gE0�BD�E
�|ŦW��? �.�x� ���K6�m���w�d����u�J���g�&�q�ۅ������o����M#�� ��c��f�1�G'�/�vZ�ɷ�L|0��A�{�u�(EGb5�لb�pǚ�=�.bl��Aq����)�Pf�I{Җ)NΖ��x��"���]������`U��V�����������_j�ܗ�l��#�G֭`y�L���A���ûuE\Y�`��(�H�o�֋���z�����-����� .V�����A�?Uφ3>�c�7����~�]��o���_�k�j7��>���F�a�Y��7����v��Yx�߆��^�S�M
��P�����>�7I��]T�jE�K��'g���[�F��/�Lͣ0I�$�G���c��S@���@��}���[p�[q<=�A����G^�)h���w	Nd���z:����':���B�g���t#(�x��;��lm�~�ǘb�Fa�&Q����*
�}Ȱ% K�bM�x�B
끝U�_˼���k6�})��9����6�����s,��=��f��6xo�rr�Y+��ޱ@��A\(�`˧����O�8c{=�h&���8q3�]���..��P�@��BT'���V����?z)��=)�ۤ%[��T��Qߝrc���;g�R���w��ŘR�Bp �5{�
��
{��o�S(��������!��]y��,���>�J�<EpO��4�Kp�QC�ż�Yg�/�QUO�I�u�]D�5�<	���[m8t���&��-�sgi�� i�߶t�� �>�K�q�}V��$�Y~'2%^/�)d��*��%��l���Ɲ���c;�K7���e���a�b���������ad,�|
!^Ҧ�#��ِ05M�BJ�`�ڪ���ur��#-��wM�xY�!�2����'��!�k�D�+� �G�v���{�lv������+XY�C�����VAR+��#��m����2m�Z�۵l'����2����Ċoo0�|���Z9�cQ�� #���A�W#�v�i�T|Zcu�6ZI�S���-����Q~�</���>Ny��Hf�7%��ӛ�33���OFO�/W���V4*�X�'`���<�*�S���~p���8������`�6x���
-$؜ߓ�S~2�C��t7�?/ӓ�j���^�k ���7�{{ j}P�I۲[���i<$����Wt0��LR2hF(��u2�,�b�Hd�+�Lj�P�+,��oe�s_Zk�����Ё�:�S؜j�r�r.���e4�=��[q��>�MILWK0�n@�L6xi�	�2��5�ŽZ���^���Y<�E#x\"� !�&�TF�ָ�j��4�G�*���<�qZ���/��Q�z�?�M��*���U�axv�xWd0��/��8l�,	����;`mQ���z��oj[��[A,>��_�"qt~y���G��]zd�L���+�>�3J��pn�¾�V�]��=!��1ᴁ>���o�)�l�E�"@���¼9K@�Y�9)�8��Q�]ൖ3�xy�m%Y�W5<p�^��L5�/3�W*Q�rn��g�a�����(F����:��I3rʟl�h��{�4%)�>&G�6��>���gt$�!��� �R7l��t��}�<F,��,y�$e��4q�8�:�d�X`	_�~o�a@�D�a���r�_����}
2;E�:Gm�������5�2&���ڛ�~?�S1źکK������'��2O˶JA&kh(����o0Xv�����_�묅���������킩4��YȆ<s���Q� �.h�lD�75se@	]���+�:3������ �mϸ�sRq!����T�*!��F��(R���9��s��/��2��*���~,���$g�dlϘ}XR=̩�_�s�2H���h�a]ƛ�Pb��6cdc#@Zr;S�7�6���ѸTE�in���u���d��sO��9��t[f�T�7v�[&��0��<!d$,���Ґ�/�3�%���)���Ĺ���W>�Q�[�3��������7+U��S=O������[1�Į�-U�7��6EdX+�ˌ��\���>"Q�����D�#��M��\��ߞ���m(D�Y���z�R��G�4O�:u�O���Tڜy��9��.@��@���gd��[EņL�u�B�-�V��!X��h�	�
�Z�mP0��""�$�;��@D'��`�/��6r�r1m�ݩ͹<����Ŭ��:aؠ����!���$�r?�c�D�������/Ϻ
�D�>~�o��i��UD��l��)J��!wx6���e'S��s0RSq5�0��j�b᧲xv�8iw����3;�y�T�q��k%�W�B�*\)����M���^�k��4p���ľ�]օ1�%Q���]��[OX����4z�����`���qP���v^�9����l��B����`
��24�;���V|.D[ɍ���������)!��k�����!��`F-�,�X�n��0֫��z>;"/0�\z�S'��έ�Dˀ��/��][�r# ���~�Y V3l�2x(�8Bt���ϟ@�5�a��pJ�V��O0�ي>јzud��d��@�c6㼀��
a�l�q�v�� 6��H_���#��"!S��)�/t��ܲ�S�5e�4��9|?��KC�dN���N�+��B�<V���C�'7��Wz�)P��x�� :q
N�,\YJuŸ6sY�±3{у�〗
}����V��b����%7;j.��'�� �����-�ou*�*�{ϖ|�Hp���i��R�e� p1��S��
g5�y
�Z��񌌹�!������TF�{G�e��<�����n\DXBA��*�s��ϖe�9k�3��qG�y������W�FN+�7��l%=Jw5�����:]2�4�|��^�-g�lgr���shB�J�K��0����"�װ�g�^e3vj#W�~ j�]#9�TJjx�� ���U�1+͏�"�H�1Lh�A~��Tµ��1��M�:0�� �)��vv<��2�4vl%jx�iu�N��@[8�&�m Q��f� �Aʥz��BW �X�Ԕ0�J��%�rs%�������RQ3�Y�H��fJdlW�F�|~��[�\��$������M^+`H���K{��:fe+��Z���VΟ{.�P�X��PK���cd[I�~vږ�n�ϭ�~C	�Kj�OR�Y�}��$HC�J= y���������U�	�^��k�=Z5#�S��������FR� j��>����2]�W_�3l1h[�����h'Q�	�넙K���9��ކa	���4�y.ӿ^�1�
��-aU���:)��ܮ��2$�#(����	)"dl�)
HH��>��%��Y�uE؄�2�`�i���h@��~g,de6S���J�댐Լ�qOHs��Qd���ZDN��g����W��Q��lf:��!���蹗a����i��JM����E#��+2�#���� �̨^i���	0D�c~�������vew�l�s|�#tv,V/3�!a�Z�����C>�ꚪ�?l��6{4D����&���,t6���:��'���9��ʼbD.��������or�k'Úv¶Et/�"�|T�������X�J�2M�^�f�����W�ĦQ��%�Q�.ꡜ͠'��і�ؑ�_�mhّ<��sZ���r�73���W�,^q���[��!���`	��Z_B�&tJ�uv��D	!�^	� 0��'ā�8� ���Ը�^��]4Q�ۏ(��bc��=���҉�vx1׌�`_��WQz�t������vѹ~9��G�e��!C��Su����d�
t�E��d�!Dy=�"N��ɘ�Ŵ0S*�C�-�'���~1�ܭm�ۊo��:A^��)��?�Y7�/��Ռ����?ȱ�����+�i�P�:&��|��9��Dz.���t������|=�Z�a�-�+V�O����|A�UH����RV f�v�]=y���%8eX7�����c��T�����95� 5X��$R@�4�t}�(� //؉���Õ(����I%��5̹��1{:��v$"s�V7k�V��.ޯ�ȯ>8	6	,# �0�}a��h�����
_i���l ꌾ_��"{TR$Arp�)�7X�Bm���l��ܯ�M�{m�Y�O��P��^�w߻������@��|"�WGi�ׅmU�z�g*�t�"��ĸ_X��
�/q���iE����!H�� r[Y��w�!�6q�3g��§eo���h��[w8[0�+�� 1��Tm:�-c�a�E)$�8$�iV�$�z����(G\!3]+L�a�M��]2կr}_�~~�!+�����ZW���~�^]�%u�F�".sKF�H.��Uؐ������\� �����?g�s3�����zo3��"�)m|�J�Ae`�Fε�(��,6_��j���I`�v���}�;ԍ�f�H���V�0P��x��a�<��o)?�/��si�t��p�搿t�)1^%|�?����~EZ�5<r��HĸUw�#dw�b��Y=�R�~����[X��{�Z#1����O��� Ihs������
u�l�����Zeۀ�{5G�@��g���o��Y�'̓�8�H�({��jBv���ĕBc��~,_k&�{O��P�~x�*�!��ɬ`�@0�4�V�顏y��lbt ��B:�����PHg;(B��#��)���"��p�]T�;��_HųT���S-L�E��TpD�~����)��t����=.�~��q���?l*q�f�js`6�]��&[O;����lƫ �������P�]�OV�ZK��%W~�S����X�m�R&ua5�:y2}���&��
^Z�S/5��B�M��wa�a�KCgeP=��V��'R�β����IXA�B@��Ƹ���ڎ*K �C�様A9!d�(PZhi̛�b�C��	�k�����N��K��Xy��tt�*�S�+�N���m���V��7J[:ՖX�0恒g���ZG�԰yY���Պr'Fy�D�R��y;��)�*��'��̙�yP�]�������� 6�%�kR��8��wd��t�,�CW�{ ?�����AU����0��az�����U{	%:��o��L��Elg9uq[�R�m�g�����K�*�`T����5�O������}�E��"�s[���{[*4��r�~&��rQ�n���$s�s5�Ը�7�1�f���{�����G
Q��&]�]�ʌX)�=�Y�R�L����-�Q(�b��)��ܽ�����q�n	��떯��U6�[�l�,\�IN%�${DΦ^^Y&e���@�'o�`UK��[����m��=���Q�� v�&��2�9�B��m����*V\U$�]�ʽ�.0���W�IM��D���P�e�$a�y[�O�d&B�CƋxf�txC[`����W�M�":l�����#��Ah�bB��M�+ȪB�8R�0&���pb�wN���GA�{��Σ��P����+�� �9ކns9��RhBw���%��5U"B��~`۽^��E<�,�l�#5�f��ў7�N�U;����n4c.��i��\'5n�'��a�^M�K�Ə�>�(�}�>J5¯�V��/�+��p 8�����:a�{W[_\,$Ii�����aO|pv�ZS��$y��&e&𩥤*�������r���+��{荑���[	�3�E4FH��Fbpş`�Mvqڕ��PYA�ɸi��_���>�&����d���aA��%���D Ll�'�W�V:Dn�{߁��g���@�S����Ӊ�Pn[�`g��Ƹ�J��Z6�ı{�s��\�d���rh���)E�׻���~��ߩ��&��:4V6��Ԟ�� �jT�k��K=k�p/v��� ���tKPD�tU�#�M�й���j=�5_z[�vٓ�R3Buj�$�6����iz@=ͫ����ğ/(�&RO�s��àxO�b����>�Wr��V�"8�6��$�Uc�Y��JM�ʴ�eP�E&��ь_����|��c�������~
�@Mׁ�dsL6�6�Nֱ�&�vkӏ���rQ��F ���Q6�Q<VXM$\�/VIs �⒯��tV�#RC��q2�Kh-a����g��Xr's�������0#d���,�y�;RD���_t�7���R-7X��Q~��=(#5��2�����5�s9���o�	���xo��`s�s�����+
��y��J��J�p^�z\�Z� (�2&A�	3� f��$�I8���c�vyy�j���b����݇Z/](
[�g�'�MR4��$�-���U-�g):��S��@` 2��i+3?�a>�����ﻎ�����|&�$)	0�F/�~'K��j��n��Q�W]92�@��E/>�Z)*��'2^�.����aQNSF%�9�I�N������D@6R��΁9��9���C��z��]�����Y�4'���;�	:�7�/\��$+'�60�t�����'�tt>��J�`R	P>�|V����}��-.T[�m�=V��G�}f���%+��Q��`�F^ΰW�J����,��vz�n����+)5�]n����,�A��*�m�#H��y]�Fm��淞%4b�FT%wgYӕ�mH�̚���&�%�_Z헬r
_�k����vZk��Ƀ:rC"N�֋�>��lOvME�a�I�F*Ա(�4Y��(1��YtH�ݍ�y��q�;�R�ah&���5���e5>�^# Au��ho3^�WPR�l�B3�o&f�b-a��l�������fqI��!��M�9��s�o-��$1�̕��ol�#5��&�������m�3I|r�3Ϸ����Y7��?C�뭗��9���w����!�����H���������ކ�����L6�͹����@L9����h����[�p�6�>ȢlOnq��!	�z�2�kp�	�/��6��!��	��,�c�d�.@���&�x^2�ԑZ>��oì�FxG�!v��!��-Q�5�s`�����&+�y3LW��|�8oi��w�L���	��c5��UM����9�2�?9��s�j�灸�N|�����M�@\�j��Tm_a`b�X�Ϋ����t��4X��4��S#�[����)�&?ٕK�˷��I'������r�Ђ�`�p�ˬ(L	�z��z妘�Zo7kK�`�;��1V�|jN����%%���k��U�Uk�^�g��~���~D�f�5�[7�%��>a��*�<�>:R���R��2���Đk���V5��b*�y�t��o8z�y���Dd�f J��� ���+n�������S��
MUё�ru8��W��5>�vm�T���I�D� _`���_�m��ޕ4�{�{��e`�&���.�kZ5*K/ � 	*W^�/6��5*�^�na�q�z7�܁?�#�lK3�-6�ę%�pR.�c��]Qe�[�@c�g�u�/1���<��z�DEƈ���·�Cos�>�ڊ6��j�"��� $��a^I�6h~p�S��z3�m5-(H�K�%�DW�*wjFv&! ���-	"�9:~��}�ֈ�Uhՙ)��Z��C@wą4�/"S0a�l� ��L�y�ͤ�g����c���쵍�?��0nl�^�O`�mf`0�V�H_��NH���4�J�D	�m���t�?ED�'�Xї#͹�FBt�.��E5�k��SB6�ߥs��r�O��J�@:�@��2U`'�����C��l�H����RL&�-�I����D�D9�]�b�W7�>��u(��o�Jq��|���@!��#&������
�Uj~�rt�8���R�Ā �{��u�@91'��ڽ���"�>	�@c�x��,�	�o�۵	#y�ܾ�����
[T��?��M^����5~u�؋���bx���no4AeU�F� ��(W�
�b�ֈm��l���O]�0���� ��H2.�_'hU�_����V��K����CHÝ�Pk��%l U�M]��������#�	�9��_A��rQ%l���а�q���T�c%c�(׍�<�n���+D��5"]���B\"'ϣ����언	q�s}��*R�ybb�(�E �f~��e��2��S�a�Ft}�4�T׽�b-��LƩ���"��R�Fl���Dqz1jՑΟ�n�p!&a����l�ަ�Ŀ��=.:fRVm
SN�h
w2�Rf�s]g;�C���O9 �C�`�l	��(�\�onif�X�S%����O�ѧ�a �ؓ��ůW:���Kw�q~|�0;4�����5,P��8��T����5��
��� ��|6��x��{�9/�\N n�I�n2�ԋ�{����M�4�d�Eؘ��[�3���S��pG>�B���	i�=�s<�d�6.���x���Jxxc\����^���l&�p4/� o��H��L�z�k��D�|�y��~�D]p���&�����4"���%���!���A�@<B�������j�7��Y�y<�pC�����!��YoxN�񈬹�ZXPs4��Z�zʷ� �]���ު��
vf���f���L�]~8�� X�ȌZ��n̚���D�SQ����QR!;�J��b\'L�T+�����k��I7Βv�c:r�l��q'a�@�tI����U��/%<�#�^K���8��iG��+p���v���ANCΏvt�Cq�:�A�>7�|<�6�>3>��/��|�y�<���;�)CN��,4�|�/���|��-f 3�h��yY�t�'N]�î�G�c��0�|e�_�\���C� b�Ma�(-@�Y�&�Oć_��Cc�ř��,n���Sv
��]�)1a)���ktC�H��]9n�MH�zd�u ��P��;D �b�Zi<�Z���±P߿�Vn�X���,�Y=o����J$68t���W�SW���/�I�_ti$|x�.Q�mx.I�d�{L�Y��S���A0:�e��R:����uJ�l��"�*��H�����@��A+�	酀�\�Wj��a\(zZ�l�qA�8��5�M�ڢ�"����B<;5��햕	�(\��c�Z��@��A��u�u��U����~��������AY�#������N0O��$oV��=ͬ�=�G;a������it�X'#�l=�\)�7�����Ljf����>C���_������q�.�$�.����lw.%^5j)�=�SH�ґ�/9�W�e�7ns!%��V�x�L"]?Ȑ����\�3��� k3�M$M��Ij��?�����2� �Բ$���]���e���(R���}�L�_�ݏqIs�up�� ��*��g�dH�6���ކ����pk?��N}z�y��k"D@D�z�'T\^)ȉ:v���Uj �1���ę1�H� �<��Q0譨��A�j1bNA���Mץ�KUQP���}#��p�(�
]�]����>�؝;=�u�q76���}c���$���a1�L�-'1������nY�{����W��Hj�ٞ��Ecި������=8��ԅ0i����m���!m��,>i��b��Ho	&�j������c�FFoa�����<L76�Bc�v�yO�gG�g��t�����i��v��C���^���j0�ܶԕj�I{)Wg��q:�{����A��'��c!�Tu� �P�g�#{I���ǻ���=��k�i���v'���Zh/&�Eq;�H �[��C�n�c�� t5����n��*4��́�a�*
Fn(�>|�(,��^x X������B�Z������b�+0CQl�C�M��Q�%<l��rN@�:�ZYQ��"[`q�j�H��z>Uڟ�$M=�R	��J�8g��x6�Ţ���o�հ����Q�&�t(�'Ϸt�2��V�)�ӰOrx�r��y�J���X�]�o<�]�*�T.:��-+�.�:J~NMԳt��,$��)�]�tRI$č��cۿ&9;ڼ��B{�����H����P|C��;�(;�b�!���T��e' �!F;�wOF�6Ypс5p0�P�|\ *��Y�E)�v?xk@Xy����ё�0C��J��˵#��B��QI��ai?�1�~����-a�^7�룄�g���;�d�L!��kz�9;M��C��a������`|1����c��u/rB4�����j7��ر��Ȉ���?�'c+��� t�"��A-��n��Բzi��-���б��5�d&��B�N��o��E�Ǻ��Oz*����Y�4�A�l+q-�@�
#�~EB���mO���� �5�a�Xy�w����4 R=c�G�ǵ]Up��uE��|��!4��iQ$Ξ{T�_�>"�G��s���.��q�$a��v�Qރ��}�����^�(ل�%),<�@e��oԁY�o�t�è�v���4n���f�עP��.p�3{�����T�
��)�U����!>5�5��l��[3j�F�I�
�o��Yw�F�gpk��0Ņx��@U����	��4q�sl�頒�Ւnj_�k	F���T9����~� �(�PÚm��]m�a!/�<��y���پ DCb�b�/�g#��9��"��n�V�է�Q��
`.'e<`��#���8- A+\�L���e�A�����`����*�O��޼����"e�(���_����Gs�:��f���M�x�Q[+����س,�YC(����dw�ǊI���^6�j�&�� ��{�MC�r6=4M��^;i�&,�Y��?���hCʍ �?�F,�>��%���^����)^�{�\�4���bR�Ҷ�wf����oy�Y�<�u5��@�V?��(�.4Lb�LՑ}�3��28���K=�R�H��4<�ω�T� �&<�R��i�~�8'm3�.��܁����v2G~=vDW��S�����J��M�Պ�%��R.a�s�?}\��
2GRe"!k���@���`ny�������?����Y�������y��OQ �3���F��-j��t�z*<o���s_-�JYnJ�9�y��عLD�6K�����6���m�5�G��/f�����N�r�3���?�8_"�yf[�+!G����oV����+ِ�0�.�7y
ǜ�3Jc7���	�uzZ��K0ʴ��2+v�v��u˄������Ǉ�P�����Tj��I�PB��+j�O��<d���_�PF\�$�$�eLHr�8>{�5r�v�{y�h���'3�@�3v\��=�����������4�s������a�N��-�j}�ԣy��[Tq��8�����mC�£��N1c�)����?tl�lwv��ňEz���Z�������S�&&Yb���3C2�����a%����;j<�fVHiH��W)$�9�uPՇ�k��' jص����妃6bC���ǽ��E2@J4cխm��� ܸ0���JI���� �G�{,)��[�F�����@#\�[I�i���Z����f;U� �q%�"�up�7�	�{��Jќ)M�/��_���Pm�T�z�2�4��mY���x�u��umz޵ yf�����|ф��[����|���͈�L��[)�~�
]�{
(���z�2�˿���F�Q��J��z�;�[�d��aI���5g�i��9E�-�,
���K�c�֫���#������(-��ݵ�]���EO$��Ӻj��68}�]c��#4��e�k��"/$C��"�?�Z?�Ur�2����l"��q�xx�(m
̱p�Mm�nx,a�F8yp��!K?�bm�Ɨ�?)GA/���l�4��]L��
�*N;�^�x��&'�<>��#�;�w`�\P��ҋ��XL~H_|TU�%(5�vÿ���e�BQ�ޮ��b��`�����9ڵ'2֫2a��o5T5<��� �w}ʡ!���a��H����oe7�l/��ۆ�i�T����v�!,�uq���~}�C��um�Ր>�d���YG�p�m���<��<�|�"Q�g"�ɞ��-o�����F�ǲ���.��Y���0lq���m�������f�}%�D��N���XFw+ih��74͙H�j$�S��P0��wٮ6�>FS�S-n;���2�Γz����-�\��1gB�ry�����s�VQ�Ǆ �֤�:^ש�?���b����;,��;&n�h����O8��Y�S�VF����Z�j���B]�3�-L�ub�A%���I3�#��8\z ���'�{mLI|չJ�y5O�V�wj�#K��4'I �@�|c%f܋��5>-[lS��4%���	P�?)S�(���Y�X"uy��7�ʥ�����uS��ʝ��OX�a&1�m��V���R`=�% ����[f;�G������f�f8�4uv�z��/$Z���&�*�.i�gɒ~�b��)*��'1��-Q����8׍��s��ΜM�R��˕c��W|�
�2���l���S}�����ZKD5���o2_偰Y�Z�@˜��<gU�	��=�J�Y|�� �2> ��L75��F��^Y:j���U�ş6�Ǐ��o��R�2[��5C��1*
���5���l�"�P��-����r|.Ҏ�񾾡�I�����$R��QC��O&�M�e�n�7aȷ�)�۔}��qy�q xN�g�������Н�d��Fi&�8^����R�}��0Mҟ/PY����6IϦ�$�VƟP���gR<�N�;6!`�P��M}�lOcKS��|U���mp(���i����O\��
CR3=6�0����ش*^*Y���̤�ѽ�Z���h��zD*uk����~���Τ�S��}����CU�<���gK�N�N%��ϔ*lP��V5�j�Y��e�ľc��P�qIC���al�*}�L������T�qD��U� ��Y����ג��/k�u��X�4��͂ra�=o��6�l).e [ִ02#ܒ/�Ɉ�OgL�1\�s~Md��3e~O�X��K}�/g~ˑ�.��E�9��Cb4L}2*�X���3TO<�s����� ����������z��jR��rJ�t�!E+�O�����ݜ�{%5x;��5Q�p0s��ς��� W�?B���2�a�#dR�����4���X���*R,��_��3DI�EW_���C���\Ϟ z˩?�|��GN��c���CD�| 	fJ�Le7���l�Uc���{p.F1�1�L�
�좦��m
�B�7/�|�ל��V�Yج���_=�z��n,*	z��@�Ts���X���"v�\C��TM��� z\�Z�I�:�&.0���0EG�i�)��r��>���K�i��͝�`�����.��0ߡ�to"��X(j������Jg�z�J3��rv��W�i��%V��NK��C�?I�j|�T`4tÎ�-UHZ�p���$�Ъ�N��ƌ-dC���ZN���rࠓ���Y�a=��Q �����(��)�O�iJf>ͭ�p/��`h��p�*r�P�ě�_V���Q�¼�x��2bO�Z��>X��P�^%Ay&%��-m�\�$tTx\U��4���&��'���o�c�ʑ(� ��y�_���D�wnxvB`(�I@n)�I"U����@(�e#�9�7(�,��A���i�X1�MW�m��n���VmY� @Ү�^���P:r_?�${�\�>��[إ݉Q�<Z=�>���^"�TKa���k�Y]~�h���&4�5��XR� ��t�+�N�!���f#�U
�p�|�Q��X?�䌹]gU5C��9��]���%�A!����cat�RT�:+?'�x�8]q���(Т�h�;�g'#�=9����kq.4��i�#]O�F!�	��_?�J�%k�	��|m��T��+�d��ȱ��<N��)�4~�1x��k��6�W�y/@�-�WlJл��,2�q�k�8:�	�;�x$�#U��8�O��G�dsU��ʦ��!O�k�ذ�O�i}�x{K�3G�ı����}���f5RDi?����잟RB�<��]�P�V�)������z\7y�t��m�)����r�8�`3��̭��[F?����S&P���Z����$0�����cF���-N� ��o�7�y#|���h��#A����z@O�j�����I!��݅J�Z��DJe�HeV	$F��	���,��.uT�:�	����!�?>e��s#ф|ś����G"1~t���m��L���%쵹���Tr�G��8�a����Y�����\�]����eX�N:0�l��pr�ׯa�}���/vi��#�ĕp���,,�<�UoWן��D�u�p������-?ki�P6'��C����YBKH��3惫��!��mU�t���f�aW�G7��8�'��"9�f�H��Eq�-m�W�9Zɽ�|�'�����(";���o���U�(B��t^S�?R�A��:�+ռǹD������6t�Ve�Ab���@��G߻��|7�{�) �-��8z<Uʃ��=�੷�h؆�;R�6;\�]^���|��ی�������S���Hf�v0fVi���x;�.!(�Jb�k.#8d�A��;0����W�C	ژB��������mCJzo��r��B�'��6*��>{�j��˜�RXf��I�����A��<#<��rϖ��F���s ��
���z�g#VEı/�YHW��U�p�� ��cyG���_��؎=/'C��bt�{�ү�i&��'�u�5Œ�z2.5.�����_�%tn�����;�ॆ˛���-��qUFW����-���Ǩ��i#Sm��B41��/��Ku۹�{e���ZZ,<w<�	��u:[�yT�oi��dh��h3b/�b6����dAf�1&x���S׻�E%
���IF��u�UO�S4}���v�̸
�����/�t���p���*L�K"4�D�Uʇ �`=a�zc���@+�G��K�SUr��c�^��?xiASy�t��Z�c�r��=����y��+}
�z�Z��E��мx����0*S����xb\�3��G���qO������o2s>N�E�$Tkr������!,Cp!?�s�(O��V��V�ձW)�i���d mU7�?಩��Jk�r-[h1�-E��ux�B��M�q��e������/!��ag{����A�u�LT:O+� ��9Sn�+�� �#�Q1��`��bUa�,c(�$�!�ڿ&:%�ƺ3�L�s�bl�d��FE�L#C��1��:��n���=0n!�z(B*G��9/lʬ�m�5u�@(i�8Sz���+�#'��Y^��_tPu�2g~2nG�1g���Q>-Z�w��f:q@el�ޮ~�G�; ,h�1�i�1e8� �/N���z(>�_���|&�B�J��rFV�԰E�0s�F�AT^�灛^q�Tk$�����*���lG�E��ڒ�}��ɏ{�����c�.�#I_-����x������yt0`��Yʹ_�󏱌���0�~(p�$Z�,�ڴ�-�{ �� �)m��i�ɀ	� ��|�_�&h1@p��o��2�i˺8�/ŏ��
�VS��2�ד�ܾ���T-��qܿ���?��oiv.�>�A{se�@�1�W�Ts�� ���<0�f'�y����wP������IY�q�g�5|�D�.��L�*+�b�MLyC�~:c�YMu\L��q�6Y{X��CxY��`�ĳ�ra��6=,�tЯa�K��˯�2,�:�0<�wq^�$?��0c����d��^X)�3���4�z�6��K�b~J��z-�P[
-R)E��Q%\+O�u�PIE�9��8�&t�P �Q�˟p�lTQ�e3N��"r���ڮ������K٣�+C˒ӸPo��vcK#F��v��9�X1-%�����{�x6Ɯ1@W\�>=��'a��Q��=��J�u�b�F�[A�&/U���\��G
1O&�+�@
E�ۅΞ���kS�u��^qq��i}���S�y9��>�@>�`=��c�9]�ni�,E�cNB!�~��xQ�dwt��:���&�p��f`�fs��S��ņ��z�K��j��"ٰbC�&:�M�k�ު�,�&���'�hq6�w?c���_G
�a~���&��A��)=W1�w�q܅!\�Y6��.u*B��qq�� n�`w1�Qe�U�����|�K����G\�����Lr�ō���Ti�ɗ��r��]
��rg����$NR<�fʻ�(c�ݶt�z1+�@��f���M�F�U0&΃� �C�[�oc'���a�2�'bd#����$Ƃ"_�b@-��I!���Hl��^d�/޹> �S
�_X�!94q*J̅�D��~!��l��(���.���otɉE�uz3�������Xp�Y�$}�s&[��D{\c����l�y.�y ^�N���Re�hQ��+��Tz�WԌ^�B��~�9�ˌ@�$�U������Gk�YO<sl�e��|f<���ֱ���Z�K7b X\D.�E�@N��d��.qB�!�W1� ſl+8��z5�К��4Ñ�����ק�O����DeQXf��zz�a���͡�^�V	$:ض���^�c[~� �%�k�~g��r�/�㨹�#Ju��f�q��.e��ņ��j�����6z���N����c���G���JQ��"���`8�epʺ<,�Ph����O���WczP�0�rz������	_�>����ؾ�rE�L�FJ#7@T}1�؄&�`�M�T8Dυ�>�mv�`�3��p�1��LB��٣�+-.�7�����p�#�jN��l��(��X� �pC�,�,��S`�=J���Dx��"�5,V�%�I���e/ӻV��>q�k�1u�x�]B�~�ӝ׽�����/w��z	/U �<rt/��|����1��m��1��
��hv��Iݡ1`nv�CL����nɟ��Ⱥ��۳]���	��:�}��{"�P6A8vt�8�F�~z�z�����^�}�v� ~�۰C�iK��n����,5��E���Ӓ\�^}r#��_�q��χRƈ� W9a>��\LO0�>��� 5	Ԃ�C���X-i}E9�������;�qm(����re�ΔO$5מ���B߿������U�E��m�g�ؖ�4P����}���}fh'���=��ǙY+z��p���ɖѿ#pn���݅�	���L����!�����p�9K6�;�=��%��716��(ph��d����)����aC�O�T�N�P�+*�AgF������M����?g,������5�r�x�n��@�U�9D�"�h�V���hLrPi�����ߊ��j����;XW�㗊*}S�yh\x���07�ȋ��� av�B^]/X��T݄����Usa�$�w�p:��"�-7�wW�N�g{�+�½P�T.}m�
E�F���&����Q=J2xxkm>�p8�l�ŗ�bw���&��J�r�?[T6?�U�ƅ9یv��5IU���iO�^��_� ����4��[�t��#&_�������7��#O��d��W�{
v̈�<�r�dx=����U����%X`ٍ��3��B�doDw�$�J��B�I*o�_^�C/��Ƈ�M�RS����/G��/�<}�|	���H�!0�1�t� 7R7Bٽ.�e���ϩe&U����є�V�R�w�_�Xf��ֺ2HB8Q3�uz�R#q��.E�ў"�6.'�l��k�����ܯU\DPj�uxi� Y�҇�@F����)��ѻ�22J$����{�)t�U��凉��������X K�g�g���3
��J�f��};C�P���&,ZG��� �$#o�Bg�Q�@(v����d���d��$�]X�YVb������͚,ؽ�=:�_�r���]E:��,�)S.�`�:5T�Yu��RK���'Uf�|\�r�#���pq};��q\@
�َfsj�-�8�SE�q7aA�S�\Ǆ2�C#1�ǧ�v����ǧ�;31��b�c�@ ϔk+Uo �:#��Re��M��TZ\�4��"��U]	(�{j��_M���d"Kf9�ŋ�oח����mSF4�dHz��`T,w��VE��/�Z�A�5�^�f��M7�]�7UG�"��bE�Ek_Ѧ�	��Ú(̻s:r���_��HG����<�]9RqNS�nC�9��o�r��ͱ��O���>'�=M� yy�H#s����-k��6w�An�v�c�NB�W�,�e�e�"린���??a���ЋCXȈ�H&g�
����=X�J(���O�*�bc%c�>�£��������mA?EZ�쨃�`#�D �.�-�vs09�T�'�^�X�o0��p~kț�g1�LI�3�m&g:._�����ަW��u�8��N�RG @�G�0������gX�0O��Q���U�	��I�Rُ�������5�S��:�U|s�����J���N�0�ۼI��Hx/�g���T�!����ą$$������?�Y]��K�y_;��飡l� �R�����
\�j
fĔ` &�&�p|Ac�PZ��Y�eS�X�Hq�^�3a�B�V8�����X��3���f�������o�|'�t���/"�C�k���>�{!�|�ӨM�~�҈��!���Q�HA5O=i�b�m�[Ī�dn�)S��b���ղ��s��I�JQX��"uC��`c:BD��-�p�{���&����YR�Ff��	lE�Z�"y�E&�N�$�����^k���0�FG����c:��_��y<�±�7� _9�`Z-��KZp�f������RIO��i�$�����XF9�^�\��{�S����	�Rp}�QM`l��8 4�o+{z�����.\<Y�b��X�%ٌ��D�1�3�L�\b�M�6�e'��5lu��G���٫c��o-��z��[�]�ay���I�iE)�'���ۍM�|�q��(E:�Cܫ�G`ӼJt��W`�TIӀq��Y_�^xj��͞s�m��]ڵ}B�F��<vdz�.�&�G�?�Rb�Q��_�81�(Ы7 ��UAWf������">͡�M2
^ O����*s΋�[k�d����J�̭&�o���T�7n9t.��F��������j��sMZ�9y���l2���g���� �o�]9�[�����z`�,�ʦ��)�V��ʾ y	��zp��I��� ����+��=����{���bF���W����#F4�Ʊ��a`?߁C�"��V�o���Sޥ���P<��ن�v���}��O���Y��@�ǻCyLAB]C�C�����E����Ew¸F�m�9�+ %ϥ��=���\3t���/d�$�DA�e�k�%�{��x�'C%�"X��|'�P%,���0�2�c��i9��s+m g���rz���3��|��_@���/��+Z��H�ܜ���SndZ;�����伕(s:Z��eٜd�g�d�ЖSzZGJ���}��|M��j ꐑgyŻ�t���o}ia���;h)©n=�j���UW���^�=��7���|
�x5�v*/
'�A-?jS�qn��5�d�.D%�T�����<UePf��5X ��p������bӄ"��^�GT%�X���4��kM��J�gA��8Od$�\,�N���|��D�#(�*�k#�� ��F/`A�6�:�M��B"vN���a�������YO�EN���	�=.(Lu��Hg%3geޙ ��LXS�6�^_����m�>�����~B��a�ö!?��?G~oҥ�����N���x�V�Umߠ�Ԛ��P���>N!q�9��#��
jɶ�4|�š�~tGf�p�a�.z��O���l �l
M_�cO'춱�5]Eڹ4��N�`�9XGMXX�w��cy��ό�{��>&�̈́t�G��-�S��P!T�3���� ��\��M~�S̨�=d<B�Q�K��5�� w������?PI�p%��n�o7A֌;�/yHB����j��]|ͬ����jǻ�ֽ���N��Y��5p�ls/�q�[�wPt_���&Reb��G�����1+��6�����"��(��]5�'� _�䡲rȏN��*![SD99���oG�寕-m}��G���k��ר�u�N�V���;
���|F滒�C��Y����[D/�tUz㊎M_���� ��7-��b*�q�V��Kߑ�o	�Uk�Bf�6��4w�W�d�вs��f�����O��f�
�=����H_���3~(Nd	}xɵ���Y�;���,u_	���7�`QWX��S
��c�e�AoE'�YP��7ȟ�D���;��_��l1�l&�~�U}-�=T�E����t���&#�dB��P�.�����	1���y���y�
�������*�(�r��'Y����ן���.	>��M�.>+�7Ҝ艚I��/�"4��r�]#��p��Z���L����Ø�����SD�;�Ԯ��?+'m��t���*`
�����w�~�Ռ]ֶ͞�2�y����f�V�noK{X���f��G$�����X���g� �1&K�#::��y�Tw�%aI1^E�* us`�k2Ɛ�&"R}�&{KP��.�+�l%��x���P��<��U���Ǥ"Jw�ЗVԫk��'K�y�����.�
�K_��bA�&�炅�r%>�CzB�1ؐ�(������9�q�A�J�Ӗ����j���c��>���P5S����S*��)`ي{��M�~�̓-�(1QRZ�Z7=_�^����J�)�/����ws��S��Pq�x�� ��V�jb����B�����c�J�4�bd|3E��LF��jj����?�u7�=��!@�\c����V�z>`�+�nhU�Aܺ���*^n�:|�+��/É
��r�_�7�U04� )���m��J� �f��S}g���V���&%���B�+C�������l��hu���wh-��'��qӑ�5��Apk_��Go$[]��E�O�mؤ;	G1����,�oOPǄ�y���e]� �G�Y�'�7�#g�)�

��ӓڵ��^��@�"�������Ef�Gںs���D�\��ȳ��-A��k_3sk"��L軻�.�����]�~�a�D��Ǔ��er��I"pG�,����1��E�_m�3�ހ�Mm�o����vtn�\X���sj߀��א�̜\�T����6�6i����?u��S7e��}�y7�+��X_89](��4�4将9/�����n n��qI��QY���B��h���k
ZNn�4t�p^�7�T�#�*cZ��^�>�B�N
�]v���Q�T���F*�������I�ۑ�Gw�����rY5�~�N���������Dl=��rR>G�Q��1�����)ܴ}��뎁H*�ƫ�[�TL��1�x0M�]��7e�ٌ;E��L|͠A�K1҄�ܺ6\n��#_�%!�X�B$;K䅧X]Ӡ�CD��/���f
�k�߈��y�y���e�"~ ���]����I�-�<���t�r���g	�����*G����E���� �ϝn�*��ՈW�o�<2�d��9�D<3q!�,,���3����=����C��ـ�~8M��J���q�b���$k�S=�tf��{��)���J���!*q��ժ��f�*���K�Y��n�#�G��
	�+6R��}C��YAW���!O!�b0;s�V> ͶO#%܌%^r�̌�i67O1�	6�_�zF�m�Wv"���S�Y,W���k(n�bi�1��8cJi-	n*j¯���������'<gw������v�T����y`���s,��/�!��|�Qğ��(�Շ��u�i�R�I`QVeh�?�L���P��O�/} �<9m���h����7N	o�
F� *��)�~��}
�IB����Td�m
�A���ޕjBFN�wcD/��u��#����z&º��-[;��5s.4�l��;|L$BUy�?�Dj�"��cg�G�7�)d�;]j侕�8nCst�T�0?�{1)�6uP�q�d?6��{��VQB&��a,��z	l�ݦ
��v?,0���z�}�<��N�6�Z~L�; *�G}vao>�P(w��(c7�l�)�1��u��Y+BNL^�$/|Px��5N�C�4Ҧ4:��Q�1�Q���~�̮*���(\:� w'��=��p.�z����/�T�0qF�3��Ss�y�@IǷt�����u�_�p�����c���MšЫ���0�3�+3	��`�W"�,sx��xt��R(�Rr�W�Y���͞&��f�z�����A߅j���Z'���s0j��ﶴS�k�����	�5/Ε�*}6;J�̩�SV�Є�Ӌ���a���͈݃4
��3�/>z.����U�- ^M�~CV:5��������{�9Pg-����6�kh�Ext��/���s���`/+���-o������ ��r��##=^Qqfvh�x��4yvϒ���ۏ��#�9��5�j��F$3`�,K��b����p�S0�1~]�164�D9<V���7xJY�%G�$5JTP15dk*\��G�n��;�{T���+2G�(�**d�t�h��p�U��
%��Xxo��QlU�B��"�mG�uQ������TI��s��þeZ>��=��n��k�Ȉ�Qv$F(I
��}���9te�7)���|�Y�}Q�?���dyj���}$������KO.�X��i�*�q���Y�\�<�? �h�8,�,%���=ɷo9�/��%?f��ƻ8��ϫ����0�Bw��W˨/Ȼ��~���	Tg��"��b��:�ُ�eU�Й���Ih��~�
����I����x���t>wQkA�q�U���X�����3�:���K����qF}�W���u#�W.IH5��#�a�$ΠŶa�_GS�*�N�XY����,A��ߍ�t�<N�?|���>��A��5�Ӹ�Au�ݰ�������>RQ�vp������t���g/����w8C��,h��Dg�]u�xU�5�0����L���|����G� (>K��\�Q�����:1�,�Y1��e��U�oI��9�q���1� ��ޥ�s�+���t���|����H�b�#g���._�a�C���iFf�f�.�����dT�Jz*f3�E>��=rRrK֬�ɦWӯ�f5����<�1Ϧ9��#6.���p�M\5^��n��a��H�i�A�9jD����y�э{�d��CE�`-V���MrO�.#���7�n���d�ˑ�?_�g���}�mw�6�>X/���� +)0o!\�̽D�!EI���y�,,p��p~MS��^qM��ʈ -�۠��g+S����j+2k}���-Z��c�+�B�#*�1(��?)-������!:�v*A�y�!��C����s�x�GJl��B�>�����S~�F�ez&��T���4�ͅdړD����\gY���\�i��L�3�eQܣ��l���?���\�&�����G��c!|o�#u���u���S�K��g ������s8���Y�Y�L���z�:��1�_�H�xDz;M�V�Y��0� �� �[����!�Z��Ĭ�$���S5�X5����p�@�S�D������]�[1a�~s�'�ޯG�����ꆜ�1����S�k���{�j�s�q�>mQ[��[��V�(GM���վ���2�`��섭|�jU�>�K�ω�dP�4<��*[�,Ъ��׬��;<{���/)��^��v��L�,�=}�!$׹}&ʀ�5)B~3v�{�2_�5CXg�Ly��<
�4�:�S��W�%O���\�Z�����2j#�t�n12�e�޵�4�Ʋq������)�%W%�D���u5�#��h�;i����8�U��P���_���~%Ȩ�e�玎�kQ������Ǚb!�1�,�3�9�U��,9I<�����g�c���� ����M��#��sY_|�fѮ$���23�
,<�1⠔ͩ�UY5BJuI%S�Y�����v��C>QY�&`{�$!3Ǐ"�QՖ+d*��U)��,0wҠ�x�I�Ԏ��yq-��U,��أ�2���[�ɕ5N�/�Eeq�G%�=���ߪ��C��f���I��p�\��z[���f���%�#�nL�}�b&y�B�Z����RW��W��e�l>ɕo
f^���'����Y�����tn^:~�&(���v�K�ڴ#L/�ȏ��}45X������݁bH��2�(W�v4���负8�}3�_vzvS?/v�'H��8�S��ss	e��z�_1�m�p{;*C��\�ˋd@����]�Mۊa�8?��{%�[� xo����tiw�Ȝ�H(��E�z���C��px7��3KLA��m�+���T�¦��O���9��F!��S���}�����o���	�ݯ�dO�W�S�D�����Go�9*��0$�W�9	����^��kN���;h\�+:�B����V�t��ͤ�:o��Վ;)|BD��MEJ���v�0�Kt_��x�������݂���7�tIq6��&QYV�������ZDR?�\��=�5m{��:?:r��Ȥf+ b�����yϪ��2�K�x���Y��E�%�	��t�x�&�V�ʪ���_�<���U��F���o���k��kCV[��t�������Ȩ�[�5��TxQ����OJ��-#Dx꽍B���v��U�e��iǥʮa̾�0��N3���a�4HO�gG���UrJo�t�Ζ���k*�m쒋�.���??��-�3�)'dQj�F�[��;�u(��c�q͌��y{���1�R%U��]f�砪�8L!���M���QJ�D�Wil���p+�b�[���!Y��pZ��i&Wҷ��.�떻�T�!�Ef'��:�/�9����N7|���w�+]?�K͋� �h�WTc�V�4�l�
>���LG���i!Pʀ����h*����`�Q`+��g�\�MQR�#��Î�>_1ט��Fׇ?��Y�y�� ��Ϧ֭�~hX���S�zi"Յ˚a�U�����r�%=���[zk	�vS	�c��N�6�i��2Riu�%��#?8��/'ߡմ�Ϣ�tۍWj!�0%y��<����|��� 9�䪹�"'�jb�(���_���Df�֚��	�i��2��M|WSn�q�	�+>�۷���vHB<.}�?,D���'�<��d��z�J�>�;P^]<A<B�Uq$��`�5�oX�"ء3:���Þ�|Y�2ex��9�.��/z��K�޶�>
�W�ĩCL�G�t�X��8\sWr�����K.*�ݰ�/
�����k.Y0�H�7e]شق��,��f������?g~PJ�z�U�v���퀗?ߵ��:$�6��M�; 9z^o�Q%��f(�[� ˙�p7���vP�۽v�������o;��\���"+&EZ�MX�䳕��J���
�t�4��"��@憑R`��+���}�$���Ly�ū���s+qZ�����C��]f��!��Ίy`y�^r��G�C����D��^2��᥏�:���n&�dh�K�ؾ�q���ꝍc�b��h��I�_�v���P����$"��~�GH�Fۅ���C"�4�r�3`�k��w�^���Mu�h�_�%�9��>{.��K���I����yͅL*��\丛���n򨴶�n�EԚ��,fd�q-�楳�rϵ���كZߝ�Ul|���Hy~�`p<����+�Y�X8�Su�����odd�@.p�
�)�T����X�5�j>
	im�ڐp��֤Rs�*�ig����	u�w�^Kb/T�S�\�n�r�@3���v�"�����v<�)-@3W��CD�=�����k���;����V^'�����пj��Kb��\:����2� �d�i��F�Q���:��a%U����X%ژ�8�!B��gn|`�7��I!(��]!"nU7�<t�M�����6�%wK���H�|"b.���\R%�%��btӬ�cЄ}/�O���SUo"�	��@
��[Ei
���yI��. �4���٣A`қ��n�!D>����X��SM�E��q�����fY�x����Ȇ������*��߰ �gY��J�	�:�Ѵ*��LOF�U����@c�=�N�L�)i����6Ә�f��@b��/&!Ï��fF
s�?B��;QÉvE���� <��D)־��ʲS�Ec6_�G����:��Y�P���ޭ�ά�����oU�H�S=������R��2��4���}��~6ڝ�#��07A	����rl���k�^�"q��z�uej�id�r��I�p���-�{\7n��q���~3��(㖜<�kw�q�3�g���U9,(�CE�h?����.�R	��C"�G�ȏ9)C�3���V�����a�=\�D,&�-�&y���a�)��\��Ba�ҋH%���r~��>
��Z� ��;�F$ ����9�A{���D�Tć�'�-D��Ҝ;}�-��X�++��<���S1��b�m>�B����h��{j7�1��m�RҜb���\�����Cn[d>7�͆i�y�)�
i)�N�U�����u�S-���e&�-{0:�&��4�48���62a�Y�d;�(M߸¨�c|u���#Q���}Fp �z<}�p�´�B�H�ZU,r�����<��
�}&�5�_�� ��[ߢgy�C����`�.p�W�S���/ON!x��h:e�"�7�ZT�͟(N�ST_ �I����>7́n�-�' ��̝�/����,IRi/���έWiak�7O|֡L��=�iF�MI|*��]�9�"Y���Y�#�S�5qNƧ-��=�;&D)تԺ�j��r���^����?�[���/u��(�Y�g�j�j�1���I�l��6��a�2FГU���Z��Ftu;�^�¿`��#T;���3�B3��aq������B�2��E�xD��޽u��+]I)�1��H�'J[��%��U�R�o�D �֙j��:�����-�yT
x�G�ǶK@�Ք� �PԆ�S�M��q얷\	#��=�^e�!�5���&������������W��k��u%J,�`��Q�FJ �_�m2*���7+�dy�GO��6�^������~=��Ph�7�,T�һ9�c����`H?�"�=f%�]eNl7�2=�+̖S˭7�x
c�W�.��?�,����ۂ�Ʋ7jԧ:E�=�1�8����$.�T�c+,�x�X�ƆC���.��ϰ]�0(s]��;��~�>��b3�}��9���d���+D���rCR���U-� ��i�.�mW,|��p�e(�tP���4T�l��K
!p�\QA��CX���|'@��.�����7�Zņy�?���� ;�u-\o��)��ǺnN8�4`;'0�}鰰�����\��G@��;kz3u4�ZA6ND�����I�!^�Ѿ���F8�pd:bJհ��nFx!��h���Y���@�B:��b���GsRI��s�����LnF�o#�����)n��jAߘ��F�WŲw r�G��mD���׭��=1�'���]+����;!\�ϲ9��wR��#� y��Ա�e���j:a�@�_Iܚev��Z���k�k��b��ؐ�ٌN�[)'�O v��=�i��D�aE���m��wW<=�b�§�O.�O"����ΐ�ǳ�]�ۓu��f�-��*��'.b���uFro��0pD����k?o�:h�٘N,��C���ct�)�kA����e�c(3��h���{.�N"�]��5�ꥣ��МV���894��*�Kn�F��~��vȚ�����t�]�KZ�@����x��d����В��ݏ�#��̷�lYO�ap_=�Zg����bE]����F`OߛZ�����{m�~�>W"�U��/��p��i/��f���Q��a֗)pj�2Ƈ���w���(���_nE��A	Q�Z�|˜�Jd��t����V���w���g��
I�[�/����~g��z�%�zżL)4������6VTJ0g��A�	�1�AiIj�����p��"��Hk͎nq��(��]��$����T����e�j_k�i֒ʷ5�R��Iѡ"�($��b�̦|:@�����`�b�>�k*���.aR�h
 ����7���tdN�d*22��B��3!�~������$K�jO^O��ߵFϽY�(%g���NB��tj[��� ~`���#����(>�_�	)��"�X&�ְR�E�@��ܭFIY��:؜��Em
���U�c��\�c��B%���*d ���R�uc�u�q2+� ��c��#G�D(������Y���Z*^n��:�t����ލd����Ԣ��:.>C6;SE`Oށ��X���.F��K���#!�t�J��Ϸ8�Q�Q�bLKpI˻�Zm8kN�la�.��"�nq�@=�n�8��qa��X�v��`�]b��4�\OSyp8�Ȓ�0SB���I������Cc/sEO����U��+�;VHA]}TrxV0�/�l|$�.�*H�Y�Di����_�u�9�Ï�V����J�H)�#vH���ᗍ�l�H.���<=��,m�1��[�������iH�ި-F���det;�U��#�.�dm���C�2��p`
	F�o�4�9W�!��мdnO���#CC� ��"���=���*�w��|MbD���tS�ck��D��ݾ�Dzvw� ��ǆ�3��ƞ��0|�xBX����1����<��9�#ȄŒ���t�M�M��)k����fs�U�9�n�;릞y3!F	-���a�O��$Ʌ�t���@/��:���8{���S���]:�x�
�3�ҕ�A���K�f�_w��>n6�G�±��-���w���E��`�x�$x��a;����#��a����0t�lǚ����( P8��k�h.7��=;�2c(�*�ʶ���Cj8�3˟��hAۀw���Y1+�8�|�<Q�p8�8	$gA~,V]��z>�������t� $:�0��Iօ��/
F���v7!ڄ��MD64�s���g_���r4#�n L���Sg������`g.�M>��y�ph�G�X���Y�Е�Y����[^	$U0�Sٓ��Xg]3�^���1���9l�/�D��!������l�1�m���{m�6p�C.b�gC�O�f�9�@��j���!�����B^�RCS���fn�Z�w��H����;>5�	��'|K��`W#O�WF��0������oD��H�����r�<��BZ��6��:E�AݏF�JR;u��tLs{��!MJ��b�� /k^ r��:W�����*��5�0sJma���P#C���J� m�m5��ݾ�%3�qy��ߍ���K\o;��� _���qR+�ea0��m��1.��R2 $�)�4�7U���S�4m~�"�<�!|X�R��a>�nH[����F�WzRR]��g���_��&<Z�j)z�h ��u\��&DV8���!��IM���ۑ��b'n;�Z�?���m�R>�<{�g�;��r��ho�!�j��(�����w�-�MCӒ3�t@b��:��;Lmx;P�1�:�N���݅�=�2��0+�P���P���`W��ue��-���9��z$�X��_���� ����"�Yn�?{��16�y��F�8�2L����6�e�Tř� �GV/]�W�R{���	>�Z��'�~ѱr�\�;����U��|�/�r��0�TOR�Ib�|���4qsČ��41�?#C���vU��_MR����5y5d��)"��9�p�4� `�F��d���X�Y����bI\v�ٗ�޶RW��ppMˌv�%1���!UA�˼=˨ az��lֳ�H"5k�rH��{�Z������6m8�u<'����H�D���(�F���H/ ���������~X��3B���6?Vj.U�Hg���X�D�k��a�:�[��v����	vbÂy���Z�3�,	�S}J;I��$��<f�
7:��o *�FA<_��a��P�N�����d�>��?	H����T�T� 6eHv6J'u}��@�+W�'�O��o'@gD}���N!	M=
��VJGDGf�YQ^�J��of�ws�&�����T2͗���#��'IZ@�g�Jr<B�/A��W
����*�d����X14�;��V�i�Ap2�q���kt����DU��=�����e֏:�̧.9�}2�m�V:�-%1�ёorZ�[&��
�j�}�,3��ٛPy}*{��N��× ��J:��g���l���Ǣo�m�r�ZJ�;���Я0�@���ԃ�O����7/���/�ߥ�͋���[�3>XU�����Q�j*2�
��3o�S���&GIU�~��$R�� ��A�(�om.���@ja�x�;������t��v��M�=4���8}�Hf�#�e<��*MJ�#C�C�g����B�d�u"Ȋ-�4E�י:cǍSh>��<��y�(�������sJ�`���2��ԝ��_�C����@�Q�i�}������d�I�Cr��i� ^�U��{��/�*vR��H��*���+�U6���Lȸ���vau���P2��e��!�S�Ú�aM���[
 �F4X]B�H�0�5gj��x2����<*��J<�8o��U=���W�IP�.n��Ԛg�m��T�d���-"�b^q|n��y �p n$&~�5�����!Q1�C���@�b ����B�&v��n�A�)��Ș:��{���W˘�N�H���hB�9x�"{�gEii�l�$V��蠰U�d�Nz�12�)o� �����h����c�7qq�Y4��O����:��[�͟q�TS3g�d�i~�&���xd��C��1�b�NHs�a1oL�������e ��'��L�n7���N��B_x��3�V�´������W|#Xk 5v�^J��To������������cT��{!�������+�g��l�_���kؐ��vZM#M�O�b	Fr���`�\ܠm��� �O%�+��HŻ�=7T=�`�>ZsqiG9fC��J�:�Љ�?Y�E��	�﹃���c���i帏W��\��� f	@4;�a$�N��?��Sp5�
:��|�����7��.i��@�+aT����$�k���q;(�W�"m��#5�9,�y����n$��T%\�ⱃ�C���K(� �D��(<^E ��ޝ�P�Dc���(y����L=%�d	��u.Ry�X�4�i0�|U:A��'����`G3���S{C��ļ����ʌ��3��Ï�#��h���2�5}	�ƀS����Sla���j?]��m�������i �l��>4C�c,�"s�S��(��뻩ɹy���*A�-º$�QK���\�
"�h��7$�ӞQ7,x��-�RG53n`ǽ~�� ��K�Z���o�A"��<�h�%d�J�O�x?��s/]/h{�=��	E�����{�á���%?�Y?�*�&��"?��\OZ8Fa�X�&W�p�={���{�㎹��Km
��r%��[@��%m�`�XwF�(N$
�D�?&`�G-�&��-�Ʀʑ�,��cn4���Õ �dn�����S:����V~��2��v%�ޞ7�'^C� y �Tust	�X��K��#�����8��ד��321?�(²0�����X�
F;�CTx��>���G�F4'1U��&�.& -���O/0?���g#n�SA~�%�*ˏSp�N���fx	�)�t������#��Tc�gܮo5좕��������]�L��*�c%�OWJ�F�UX�0M}�1KN>�.[�+�f"-(6,�#>���S�VT2���i���§���~s���,F�<��̓F�k}}E��w஥\�	��T�ν�ü�Ò�;������n��Τ:aG0�:#� ~�g�d4-�H�����C���]�%4$���JmvlA)�����7&�3p4@jU��k�T�\MS���<�|�����%��FP^m:\�B�K���e�@�e�E<�e|�  �`�S���Z�v슌�@�.�/��mQ����<]��/�::K�&�	G:A����G*�B�����ʌ$��ȴ賾ɞ�ëOMN�92�r�(��k`�ϔ,�D�eW5]8+����zDQ�<��ţ���v�]��H������;�	$����L�J�c�A�Q]��� �࣡	��H���4ѯ�o0��6����ew���}�ǙL�b�8���p�+��B��g'IF��m�b ,9��[��Av=��^�`{˸�.�!��-.G�?&	L��n��r�C���� ���r#��дs�o����*Jи�tO�@�B�5CD�=�?Q�2<h�q�����B�p\�0o|�r��$�`�_����{�f�B�yҜ��`2���p��4w��J"+��yҹ4�[�`F�W�
����:8t&� !�E&�����M"��Q½������B!��O�Y�q����O�z�$����b���?��!��2����S\���%-<�H�E�{�wBQ�A���̩7�G�_ʗLLDi�*��.d���:2�U���%4A�"��4��H��1r^��*�Ȝ�n^!+��%*����^�_i���%H!>�[�m]����@���*�&����K�O��P�u��L?�~��@�K�@�ѻzܠ�.hͻ���9���M�P��U"6� ��(d�?n�cl�q�C`�l���c���0�!TX��q��C6�j 2��H�Ⓦ>1���*�q��M��o�5�w�:��V�˒����m�qPH��O�?1������8�{�s:h�R?�����	\�]G�T��\�'Mr�F���XJ*��bT��� l�?�]/;���_�_���2�!�h���ĬIO����z��8|�9����a�}���N�X2�E��ĭNUUlE5�t���'�n_]es�I���N�S�H-��Ojn�-���lh�(��[/%��a?�'\G��t�Fz�aK��r�3Uej�;����y��}��L��j���v��7[�O^#��w*�e�g����v~�>s��,�dVPL��2�ca=�|�
O��rm9�E�h������N��u(�@��}�3���e�����]�w��(������O %�k�=@�w@��­�yf�ђQZ�SjL������Z����O_�F�������X�B76�����y㓓��s�3
��ܗh:�8Ew9Hv��4LG#O_h��+�"Z*Sd���乿<|\]��۷�Q-l��Fi���~��aNc�$l�8�:{p-��~�>������X�ՖcLgܹ� �&M��{O�¢C{�.FV�}9M��4�.)��_g�H�=�o�n`�.C!/�z�������,�9e�:'���܍$��i��hi��ƛ�1�}G0�=�Q�|z�{����n�]`���=�-Naz	�ZB� �&,X�j|x�\P�AF�T�rvE�~(�6+rU��b5��[��Pzs�\���=(�F&xz%���j([|� ��-1�="/��'�¶%5M�]�À���R�CG:�_@�.��V���a�e3j�n6!�����z-�����޷t��,�_o��j��X�e�7⮒��*�k(j���ѨE*vh�a�p+v��7wABF���qQb�7��S�7��c#>'6�qBõ$g���0Zy��<�l\���U]�j�*�a Ra�^�3|;G�CP�t�F�,
-@ide��,a�-�39r٭a�X�wҞs���H'�o���7{��L���L6�����Q��Zq��eխ���	}��gaEP:�{nZ�����@]@L�ߤ��ɾ:��翂V/�k��!	�U��Bd�pi�oϯfB=�q��$�Sbl��ڡw�[�xp��u�.8!A�?1aj�{�epN�Rv��s�ܠ��6#���XؼG.8aY&(�-]�0�\����Z�DK˻�B�eC����g��0ֹ��l��=�q��u�ci����>��K�?�zy���z~P���߳�����y$�u�ʟkl<�X�fxB�0�9`ӈ�
Q�	6Y?aO:c�m��8�r� e�z`U�.p�%E��a���w���_d�|?���� e���F_2�W�{�z�'�>f�M9�t9B?:���R_�e���~�*�_[Ȍ����'�Â�1���c.;V�"Ƹ+�$�v���r��v2s�i�a1B��\�q5���Nh Dg��'.\+�f8���j�V�q�k0� G���Ll=I��ox�E���LDZ��tϻe�ȝ!T��8L{���a�@�'����pG�ْ�&��8�+��#+7W��G�`D+[; :c��`8Hn
����z+G�;���~�^x�Q$Y{8���0�ã�/!�\��g�!����k�16#B�;�P���s�~��}�c�wydv�Z�����>`K�����7iʴ���,�0rG��P��dS�(��x�_|,�A�h�
��A�$I�D�j�|��:�E��bk)��~�kIhD�X@;2ϔ�+tq�C�[������=�陯\Jl�E��N���q^)�����8�c}+���;�߿`䱊p�)a�vS�\�C������Ŝ�N�M|D"7"3�TG%ϷQ�NvY���9�����f��=Ss5~a�Ro�nN���)�*:�4�����u��=s��"�2����X�w�15��\�~��s���MPc��<
��O()�e��L]��{Ɓ�l{A�g�f�s<0��	�2*�o��Շ ޵��u^$��VV���y1��]ȓ%oL6�^R��ג���m��_A�ⴽ���f�����2�ʌ.P�4k�jjd�ş�?�{�=����s�`�Qa�qP�4��Hj�K�_��*g�