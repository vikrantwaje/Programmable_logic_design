library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY LAB1PART3 is
GENERIC(N:INTEGER :=2);
PORT(
U:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
V:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
W:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
S: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
S_STATUS: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
M:OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END ENTITY LAB1PART3;

ARCHITECTURE BEHAVIOURAL OF LAB1PART3 IS

BEGIN
PROCESS(U,V,W,S)
BEGIN
S_STATUS<=S;
CASE S IS
WHEN "00"=> M<=U;
WHEN "01"=> M<=V;
WHEN "10"=> M<=W;
WHEN "11"=> M<=W;
WHEN OTHERS=>M<=(OTHERS=>'0');
END CASE;
END PROCESS;
END BEHAVIOURAL;