��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#����f�RP���J/�i��/����� �� ���!+$A釿Q�ex���֝�[��!��3�� ւwx��;
:��R�Q4P5�p�!h�X(��ݥ��Z'cS˨5��/�;O�=߮ҵ��R�EjۛW��ӧ��w��4/p�y�Og�*'�\�3P�Ӝ+�9
_�؈����kx�F����'�"�p0��dD����	s�C����eNB�u�z.{�c��WzT|��,�f>O%d�^��j�[�zw�ζ@�&�ሬA7[�T~u�j�B�

���T�M^-�;�X���n�L̂� �0�2�S�{B*�w ���}π1@׭&7���Df�E�,��T��Bݚ��z~{�(��sUs����	ߎ\��� _�����%��I���s���P�{��o!X-��S��)܆In=j�}�ÐP����������I,��%�A"PѴ�3B�ʑ9rӿG_Bu=���+{�5�З F��K�mU,Ĺ��r��<����Q�}�]����u���yZ�c5?�6 ��;��"*���bd]��߷l�D�&u�I���"�x��D�:\L\!��X�)8�ϔƣ�c�[F�x�(�7���˟�m�~d�/�O�GMs௵V2�gt����6^�#�u򀊌�`[׌ׅ��b�Cϭ$�"�Ƶ���m�e���-�	Xė�N��K���O[�p���}����JX>%�0e��q��qd�M2�)�1T�g�Ӽ3��~���_NF�
��S�4Am��rdnց��B ��w��+@xʗux$��Af�ת��ۛf��6����~�Tٶ�~����V�m�j���&��1�[�C7;�'˕i�Q�Gә�r��*B�mײ��y�S'�4�<�ǥ��i*ԺY�.����t��K:x��qa1S~��h�7���m=�94ctE�lVlU~m��)��6�w�B>���r�DQ����g���g�%@)��ꓟK!�d^��������e�7���#��$fx������O75E�J!�S�����.�3��Qe���0��t�Q�!���ː��1~��P�h� ѱ�]���_cC�}/�*+:�����������*l�B��	���.��R�z���JZ
�o�::������fh�"�rϫH���S�#'�����RS@L�r�x�qo�_;�|�{Lm�Ǐ�����?�'y� ^�[4}����j�qe�Ϫl]<��H���އk�Åި��vy���r��]+�?M��"6r%����W�\�+�Ē�{��Yql����i�bn=��H�_��R~|����UM����k�a��d�G�������\h�ޠ�5��ܣ���~ k������決R��F�q�J!�h�8c�(�m�)�)D�\\O�z��2/��Ƥ9�٫y�(g����r��I0UO�$C#�'��= ����C���.�	]�jɫ�3:�L*��OSG���*
Y��Ҳ�15ֻ8u\��֞��=Y'D����r7�J�$��%����^,���� ���j���G����i���Qo;�$�9��B$���RU��Xwt�
��߄��(wܩ���
���/�|���,���@G0�.�{h0?~B��'i�;ǉ(�VC*�z�&��\{4i�!]|4C��F���w���$R�J�����|��V&J$Eb^�xaz���g����C� ,��� S���.x&6�{�X�ׇYA��:윤�%H{��u%s�6���Vv#%�-�����S��xo�6S�l�n��k�Be�Ѽr�7�CC�S��F��s�̃�د֗�CZ����cs*�̈́j]�] C.������`�M��o>h���ǠLw_�Y���˚��������tɳ�7@��)g�5V
��Df|�S�n!�����]��#�!�׾���߯�wջ_Ex�6����z��#���Dp�t�~*����as{]``�v��� f�Ĭs[QIys� �\ې�[q�	�5:s\Lhe� ��s��3c�ŘV���Z����9�96@�WD�}Mu���ۺ������o
A:���ߍ��Ɖ�a_s��	%��n���Ęq7䅃zdߍ`�/Jo˛L^��=v����o�.5�X��}tQd��@��y1��{�Щ�'Ͳ���}�/ѩ��I\�s�r�x#��<����"�_ܦp�4�Zg}9 �ن��)rM���|j�Jh	w�T�������!��uu�ˈF�Y�Zg�cܡC�J;����?e�?̐5v#�P�C�U�ۍ=d�/y �g�W��Am,������f� x|�0��_��?�h�h
��*�*����*�*}� $��<��
�6�$]���	��n@4k*�w Q	��������	�S����$��K���(qG�!X��eE݆t�Fl�Q��4+U�����g$�$C��@b0�%̈́� ��+M��*� ��D��.��}���
��k|�vL�X䴓-"�jc�0Bw\}z)���Mu���ɢ�z{آ�[��
X��Գ��,��m�N�<53%���dC�|�Ags�x�"��/��\�������V�^I�̼�C��IU�E`+��0���:M(L`�Ƿ�+��ky_�}31�r1��Q�Ɲ��w��J�U���u]p0Ư�%)5�eS(�Y����w�.�6�1��n�?�_U��:��^�;���"C�%�v��rpu�����Cy��X�,���	R�D%�Ki;X�B��L�p����PC��Uʨ�uW�v<(<C�+	м��9	E�����!�K�
�D��<������-�	�e�K�45;�b�/ŦA�D<r��D��DN�+����E�ƞ���Xzx�j�Kzʱ'#�7H��e��@��H��|�K0q�Kjl���J���K&:�0��xFB�X�Jڜ�aY#��w��ʚ��&�0+R��0�(F2��غ`���Ɖ�W�)�`�/#��I�N���:��0�ZM���k�[��qNF��͌bne��Ѱ9<��I�X�����Ŕ�� ���k�Jl�t7��3s�����{7�|������o1��_��Rv靿T��`uX�CCj�jĒ�^$ds�(��K�Z)������et��Hz@i�	-FQ�H�=wyv�oP$73X�vp���ݿ�Ʀ5��^�	���ǮN�R�1]�h�Lc�t���>#GMn:��e(�诲7DzKc"���HZM�Pˬ�q�E@(���P]�R�B5�̭/c~8<��%�;蝗�e��T��i����!��+~߆�3	��*��~��ߥ���߉��C_�!�py�H4S��<c����x)l��XWu�a�+�ǥ�_F+S��JA�J7�:���J����R\�m�4�C�O��~5�|Y����ӧ�q��a���nT!���.<8���8�c�L�Yg&Op�����V�t{գ��=`�z��^�K��	�G�5��W��åԙ����`�HuA�	�L��e��O����^}��ﷷ�U؍AU�d�>��!����[�^�8�lR���x��{��H!�ˋ��sl痪������h6Q�he(lQ�ُ��7��%~zkԂ���ο�N�9!�5k(B|�F��j���G;.D��'�
yV��д�l��٥?ٰ9��q[�f�E�`s���O�8F�NC�)��muI��v
�=�_#i!$��K�������(�$���7�¼7Y���^�`oy��
�&j�!^ri��g�ظ������.��\�(��Y� 5�^rEs�K0�@IcL��v�-�A�SZJxE�*U�9iո�\�Ot9ÄV��� ��D��*D��9/G ��ܜr�>73�X��	M��o��z�I��|7ꢟN���/~ɔ9�Z��T��h�jD�ԧ�o��%",�������7ɬ�}ΰ�|Tdo��Hnu�e����ի��t�Ch;�olN�'��CU�Q�}��0ڮ�7�vP7��J~b��T�@�"��z�e_ތ���e�;�6�M9.eGj�� y�\vU�-�7:��$��®�W��d?�L\7�)\��5��kf���PQTT�,�Z�h��D�ct��Np����!�0w]�.���y�7��I��(��	�Al_�5>r�y��_��9j`ir����`GÂ:�������P	R($Γ�ߦ�k=���� �G������|	����t�/��?<�,z���+h����ؚ?7K-R)���4Zy�z�b��/_�J��j\@�ݕ���lP.v�Z��=��F�������.5�`0����Ye���e5�v8�|��@H�Uό;�	
��OIa<^�6ņ�~T+�f7m+�r��h�,^D�E�t���d�,膟m\o5��ű���\�A`�Z\�����#_U��P\�O� �� �tI�S1�Iho̵�������+_zѬ���Y֠�,�e�n���o:�f&V�HW�����i�ߋ���s����C�/�$�|ʋ��B�Y��Z�Ge�L�<���������m����p�p���=�2��%��| �1��&}� ��H���[�UYӥd.��P�����e��?L߾��O20���Ց�J���� ��+��r�}K��\�C%���X-�u*��m����[�5��D^���刷gpZ:����o����U��M#{��$~6��rγL��H:�[��,v�-��ܘv/+�2?�NM����y���W�E����-E�0͌!'�J��墫�h`%��{�Oj�7�f��ų��}��!Yc��N቉PI��T���|���o��+]L�ì?h4�r/��pZ��S�c����=���G��I�LF2��p7d�����yNB�c�
�����ә�b�>a��D�~JR�\,�s���L�����!�nq������߸cl��"JS(���&C��Z��j�)�o	(�{`��f���Y<�7�>]�c���k+,jp�P���R6�@�|7�u)��ڶ��@1���Y�����:G6{<���ݘR�0i�f��N'��>_�d#geן��37j��9����sQ�����A�PS��@9)Z�w��Б�p%V��Q�u	�g<���my���熾��M�c�d��Sv�^��3��s���G���¡WZ3��v޷H��+=X+�]
XÃש�[�G����b�n,�i�{بV����:��y����	;ó�o��k��g�q.�Fީ�/<z�h*�j����4�~�(1��"i��^"�� �SOe�EJ�<�i��_�(���Ԏ���4X~<V����(g����у��$��R��yk���e��a#H�������*s ���SR����a�ps �Ε�8�r1�!k��Z�r�������x5���y��_;�7�e�CS�u��u��x�01��`w�(�9�� �s��;<?�����Ăd��HB������'^��y���Ĕ�ͷ�c��UG�d�\�S��̥�TB��r�O+�k���?h����5��Ƀ���A�����������	[~�/������Un�o�ۤ:"wp�7�i��OMȔ���9�Z�c���x�8\���>2��9:�~���m��	�.1;�\E���}�'�(,�4�N�J.�s�+0�)�rc
�s��ʕIx�2�04Z#��xL��Y���-�7�.�Zy5�>����(�ޚMڕ5���!/�}�:�!�0���r�� �����s& "x�DR�CԽ���0��i 	��h�o=LZ:}"�*=�W	/cft6�g�{���?]O�ͱ��:QG�,;�w�o7�n$<��B`�d֏��\B�d�-���s��T�%+D	��d�
ö�Ƚ�Q��}��>��lJʁ�Uhyv-��]R=��&
�I_hp�C�="�����Ie���;9�<?r�L�O�E���4-�	J5�1mCyEok��g�>���WD�&t�j�4����gD�&���-sr�r&4�#�Wk~4J�
E������K�jE��ۃ!
@��#1�CDR��0��{�=��P_�>��ap4L�͏"��,��h�u��l�=��[�y���h����1�??�[�+f�q(�7N�?>��ӯ��am��{��i��FiK��@�^0�!D��oc��.'YI��G���_:��#���9� �R�@��r�>�?Ԯ��m�i���i7�����
A��'�1@�f.��{���p�ޯ��eU6���8����"]�
2W3[�6ba�X�����}��I6)�����V�|���^�A�B��!z��H)ч	��MK�H��Ì�'A��;��tmY�x�-���n���V>Ţ�n�����W��)���t�"~5m�^CuJ���aL�>���ѦKౖ����,�'Qe���0�"�(,kt�v��מ�O(鴨���/�5\��]�y�����u����3�E�G���N�u�-HDmpp�j����۶�?�ݛ�A�����s�?��t��-$!�U�i�{Z�<�-V^�<ջ$���7Ń���V�/t��������r%�]6���aح�H��q�A��eY��A�𠤉�_��ߢ�%
*�tD�/�g�0D2�	{Zqu͟>�#bD�M�P�kj>f�s�Ѐ��<t�B,ny�Vk�@
�Nw�� ����Z�,#(H���"e�W��;���ʭy�������~*c?�x��*W}:�2)R�7�E���o%�������p��i�{��4���ks���Mu��Z?[,�1�o"����5�vN��^8}�6*51���{�AH��t�G#�Kֿ�g��2�]s8^���t��x��"n8N@�
��/�Mn�.$�
zlh�Eϓ�0���J1i3e���R�?��&, &��<�Z����(w�W��	��w�MJX3� M�������PVk�mU�/���2z�|8B���#k�36Ӹ���zA3�q���ڎ���sT�+�i�vR���mvov�� �����}ݓ�+]]|S!�����{����-�e��gQ)UE^-H�&�se6��%ե�漁
�U�x��z�3��d��t�c�>[��[q֬����Ԇ]��A$�f %eɮ5�|��y��,�G8�� �] ���*�SJx�E���&�t��ê��V3�Ɛ��[(	� ��n�r�Kg����
W�ݽ9���jT-��ibb�a�x�p��s�o�t%�������nor[�<>-���Ǩ��r��b�aXbw�kɏ;ã�)�/QX�h��[���x�_rͥ	�!��V)�s�B�+��%5qD�p�O�=�ϖ��P���*g
��?�uC�?{��l�����\���Ɣzw�a�1�y@q�����!�֊�R�F�%u�e (�:uS�&���I7��Aɐ) Q�m�b3�$���e�!�Fj_	O_I���/��"r�T�iCr���Ⅰ�@�q��H!Ǳ�����W~t'��P�w�"�n���ϔ?dtb��k������%���~�W+U�p�@I^��[�"��J�v:tB�i���\������ѧ�
h�cE�~縃�8 ����4�eXڄ�0mA<f~+QM�9OOCN�?d�"h*F}����V�܂[w�tK���~WN����p��97�J}Z����)�]�9��qWu{~U� �c����h��Q$���DPԸ��ymw�����D�░��,�W�l�m�\�/��%�A<#T�T�H�';��������nz!��/XC!�or=��ٛ摮a%_�|��k8��P�E��6Y۽�+�3Ѹ��8�l����q"V"mC3���f�����7��{��Y*1b0��[.#��:O��w=(�U��lH�(�[�\�}킇)z���ݑ��LV�Bչ#������\-��t"T��p��VV�������mҬl3��#��T���zG�7�,뒓����w4qw�k��/�����q3�ţ�6����Iأ�����1������S9�`�4�2��d�UW.o'��?!�y�m��Նǉ�s�䩮��ܛ��e��L]�Y.�>���+N��{�_ˏ̸����#�m������(j��(�z�P�A���o���r�C�Z|���`
���7�_k_sd����#����W�8G��8��|�eB`��p�E�~ڗ~�2��w����ӡ$	����m"�e6�`��K�����gP�s0o��`��־3��e�s��T�J��|��
Q�v��,���p�-��qz��O�2���յ�b�x)�H�ֵk�?��cs�ē��|���h6�kZ�]�6����O��"<1�l��8��eǇo]1���r��(�Sa&�u��ݒ4;NU��ͮw\J$��8����UY%f��p>���8�Z�H:_&,�#fz�c������� ��	�:�S�a�T���S���c�~5PrW/�����W��t¡k�j/� �tC�)_�$�s �K�b�����D��B�ƃݵ*Ҙj6�萑�F0�uEƮ(����0�9��d�b��f���ԣ.wh5�\�k��1�S[U�Т�x�Y_T����Jo�ٟ��c*z�� *��֍�6X�;��õr�=.jӒ�v,��X�S	ǲ���� �6��֧+9��<t����$��v��ե�����GI�B��?c�3"N��P��fVY0��F�����ҕ�ƪ݇T�*�ԗ����b��f���底F $1v�V����j�`��L��Z��OOS��w��4�9&�x �e�2�Ȍ^�S+�V��\�{+���)30�	]���z�$��-��-o�"�Y��i��n�J�L�3-�|��jVQ�Y�t�Knы'�C��M�T����\�_tՈ��P�Ԛٕ����\�swp�)[ຨ���'�'|��pͪ+عİ�f*0>T�ݒ,7�eK�3�-t�$�k� ����a���ݿ(����@R��oj���rL���������ۡn�>�W#�`2�9�N�(��� �����on%��̘vk,�x�?�i��Bv�!Z�WLt�LEEۄ���' U�C�#��E(̘�l�uF��3�:m���o�-)]�8��py��� kW#�It:R�2��g�v��դ��umv�X��9�N>틊��H-x��6$��9"_�7]L�pC/y_M^�K}/�D'��V��ֿ8�ɍ��C�W�%+��9�*�-�P���U{�G��;'tI�s�����5ꮢ!G��X]���3�vK�v+)���U����Hr�R=�eW��箙.݉�r��k�,�����b���i�iJ�����Vw��k<)���i��d[^x��V
��� c�}�'ɘц��87�o��'e���D�qob��<�H����7��d�y�c�9��vSi���ONh�$�9���IsďF�B�*���E�Y=I�.���I�����|��5�Q�q�]4�����_�Ε�*��94���	�I�CC��ݔYMY�<�.(("_3C��+�Eam��,)�0�'�9ck���+$������"R,ܧ�%lb�:��,�8���M<��Rd4��5c�?��[�T�5C�YF�p�K�/�LT�8�iFpw���
�@�vqa��:)hYw3�{9���c*���'z���nŠ��F�e�BCMI��M��ig遈�e����E���2&���-��"}�Y�8����.�R-�>�-���f�#�L��&h��br�B�W�.n��N����,�(s��g]
��ᎈk���P�E/����u&x(2�4�E'���g��$��`#��#�`��M
��&��g�8M������l�� �0��[��@�}T	=�*|x����{q�)��Y�1>�"yS���Â6?g��Uh�{&00S���b�2!�'�Q"���F�Pq[�w�1�`m�/0~-��{�i8�$�g5�ֹ t���B<96��3H0�D3:����׽���~�g[�7X������n���7�EK�k���m�����TT�������11Hp�%AKy�+طy�Q�q٪��嶯ɯd[d�&��z������>��L�,��06 0�n�/��t�\p��yp�Mx�r �?��h�|6o���ԯ'�R9;v��FFI�U���w��D�x��m�8�8�&n�:4��õl3�O�����2�i*�w���	۵�G�F�S�����I�TO�,[;�sAK���E�>؟�}+����7�����w0�z�z*�{!C����;>ߤ���X�e)e�Ћ�����u�QKj��{�*�-��[r*"8������?$>�b��|i}�oѷ��"� ��z�$��h}-�dw8M���)|�����3I�9���;�.�nX�4��M���R�y��(��5n���M�Ɓό��1f�6'�'��(Iq�76P$V����F;|<?�DP蔞��Le,#��$W.���,Y
�Z�)T7���6�_�UD_���\��t����,�%�(�L1o�|o����7�X���%`�$,f�l��6Z@�����t5��β�������5x���ǖw9���rt���.�����*g�U"�0U!�/�� U'J���j�����"��f%'�V�	�tRt�/�[a4W6�������u�2��c'�Jذ�����������9'W�&@:o���.R ��{�5
��@�$���7��=��*���?���[^lL�����l���R� J�Ș��_��8w��)�Q�[�5�јI&)XD��߀��agC�7��;B�H�0���ӽ6�R�H������KdED���Ёee2/��P�fL�8u���l=tO2%`Ί���ڕ�4���%�����.BjF���b���o~>>�?�����?�ہ���e������5�1ԐX�,c:wNECS�g]޺*���`�/qy���;�U_H�����g��*�����6���}_�aI�O��m�����&�ʹ�=낒��(���rl�W!���Q�l8[�W���b3�
Z�_c���H�\H�)-[�nU��^�v�}u
*G$�3>O�ͱ솙j�M�)q?q	����*:�2T�y��[]��`G����(6/���K�`�T*���t��K�l�r��eE�_G����8���ы�f뙠���lGmT�=���⼴u�w�8�l24V�uhn���S�4^��̊�hUg��!�<8u��zObV��X��t����+�0�����ek��-[��E?O�p�V](1!{�t�v戫sGz���W�e�B~`�d�'"�rwlܛ�+ϧ�燏i.)��c���X||��&Yp��+�'uY#�������á��V!���6�Ss �Q�u:������N)��ʱaa��NL:�y�z��_��e,�Ѩ���g/�9�$�)u��u�1YK�=�:��$��j�c:��w���	�/���N��|�!k���y��a���k���؍��a��q�8#o�zl�}�b'n��d���D�W&>F/s1$8Ʊ	D�6�Mc��Ŝ%�]|��X��_#6ȯ]1 �0�X/J�Z哦٠�7��Qk ~iDV���!�LB�IW�a'�=)0Y�СxvǀY��nj�S�H^F��@��%����xt{�%��y���� �f���j�H) 9�X-�H��0{L�V�L�RǬ`j����v�T,ʊ*;1����� ����ac�m�b3B�4kx�`���2���t�uI���-�7"ȍOt�0Wt���,�k-)mwVч�-tHLM�e�z�Z�ȴ�Y�T��}#2fGَ���@v��1!�w�&YXǩW4AI�����<�a�`�S����0�M�e�`;E�j7t��芏��[�;'�)�G�.K�,�����Tw�u�c�:7��֝Z�Qop^���A��Փ�3R��n���=��v������:�J�n��+#��rR0p�8�����n����E��?���¢�p6�2I�ܛє���Ԧ�=D����2�m"j�ɹ�	�)Q�{3�Wm�,a�?�*�;|\�;������0:- z�G�u9�q��+�I&�*#���I�6Of��g>����~���o#�'�R׊N��[V���W��	�XC�1R��9�pJ�U60�U*��f?��J�w�:����{l �y�.j�}D.)�vQmW����f)g3N�����V�nLX�_n?����{/A��9^�XaZ��~h~�6O������q��޻t��I�:��ZY� |�W�ZĬ�}�0jM	Š�}�t���u��s�
V$�rq�aR�^�2".MO��&�P��"��r���k��R��O�q��7բ4Qa�����j�j$	'3V�:�J8W��\S���&�'Vh%LdK{��ƨ�[�2%�za�M
2�>nt�Pu�>T�U��Y���&c����?����s4�/R��T�Wa"zăY���74̕X��r-���l���Bx^���2����rh�rV�dן���t��fJ9Y��0�Y ������c��CB4l��B��/�O����ɮ�L4Q�@8�h��L���ݡt�3z�j�o"�� ���/������p��an����b��|��j��MP��6&,v�Sq�I�d��0[�z2�ǰ�3��n�6zM����m�iC6��8u��	�.��9���������6a��v:��ˇn�>�N�T�qS�1B���r)1��5(L��,0�=	��m�X����ZOH�z�pn�)���	T�
ќ��ϙ+����g\�
\�[ʤN���X�O�%!�&_,�\��6\�o[�Z�0�GP�2)!H��Ǣ�K,����˓㛬��Q�5���M&d���8�#��n��K��L��.?��5���\��-��]?�2����,�nG6�>;�����0���zetS��W��#=l���|T�~�g_��ů>��9Cf���K��>� P��a�eDt�	˒�j�u�':D5��E��rSNwH���VaB�}2�VC�n���<�c���<ݺ �F1��$b�Ib�H�pj1�j�y:���ö-�ac��ED=�u�$G�!�����<�FKA� �������c�ry��i��D:bq�<0!6���2
 E8����t�Va-\�w��mK"�f�&�a���
�� .����ԃ�$����ʖ�H����B�Xrؠ-W6Fe�=�S�o�WN�tڜ��T��:��Hi�Ł4|a�eu��539�MI�t�o7J��S`/�A�=üM���QKK�%��G�:ǉDfo+`���FBv�k�F��3�Xk���0k����9G���DƇ�6R�� �������#0p��W鎖j0h4.D��2�q�Z� �]�eL�.�WU4�=_���]�8)�p޼���J��c�(�����u����M{��+�Qy��A4�8c���ċ���sg��g�\���i�6g��DS�ǍD��v���P"�uH5Tg��^,�׋��C���_��r�ɶ���У�o��U�X5+�����]-أa}?섴�`��8�K����H���9\�x>�&}�������J�:Wp�PR���}C�ƣrĽz�K���Cj���O )xQ:�o���&�@	ϫ��uϘ�j���̔��W2L!��UDb�-��Q�.]��b�g��/Ш�b�d�/GE��׺��x-ZYA\v;�z�gG�|<� `*���6�z�iz�k��t��7��T#�� x�f\.���ˎ�@�W����\h��A/���z ;R�-�Q�h�S�]'C���!�1�]��f/H=��ggj�GM���`��x�y|�krF�ԡ1Ɔ��e�	��`v�sGב�Rє�g��!�8�s1u+�ƕ7)��2�\̕��XDPz"Mɑ�G44���W�]a���E�"�0�]�]o4��v�����q��WњP��H(�C�4��o�{���|.]�j�2F�CbB����%�� �7�@*���8�_���\>���CN)rdw�K���Cr�
e9�-�B�!�ʋ�2��x�PW�;�:����Mo�߃g�w� 2��֚Eb,�A�q{"(�B1B9�m����N�RLC�٩-4}���&_�;��@�h�l9�h�a�����b����Z�ƃ�{�Us�΄Eݹ�-1Zk�i}���x#��c|.�Jf;�,����t�����{J�'ʼ�=�d�!`�K��TXd����^JP�)X�M�h{{�Ga))9́�Ie��q�V�e��y���:w�Gt���1���u#����3��}��4�P]� �O�<����'����gH<��:�^u���s�f.A�TrB���T�$��>�c�`a�F�S>�n�)R�+��U��L�A����Mw�:#B@ PG��s��[�_/=�R,	���"!���Ja8�
�F���SQ<�����Vr�fHE\���_��ܔ��*<+����O��	i����ӥ@KMz ���ۛ��Kϻ���17(鄳��5V��+	t�f|�)�,R=]�TAR�:F���S�an?������yo����&ϥlL����z!�vU5�~��j!#�J�g`sCa���/lô�B!���Y�z%l��Y�M���F����ѿJ_b8��OͼGT튆d��x*6b�A���cOBp�~E���@ط*�W���u�X��	��� �����4��Tn��Ъs�6�2�
SL� fHQsz�6驧�b�YݽT@yUHٛ�&4]�p��O f!������Sr�Z� ۱C���6)<]�k������%$c2��Çٓ�Y1*ҿz�D0�BI�g��$��8���.�O��P��6�����
��t|�r�>�3�&��^��-D�/%1x�"O�@�u��mS���D� ]l�,R-8^'x$������M0Hr�Ѵ��Z���<�QZ�{i9� N�yv-|��S�;�2�q�
h��(��Ŀl𓿭I��؞#qZF?B�a��8�ȿ����%��S����?��R��f��]�Ꮉ��м9�yx��r|��Yvo��O����3�,֑^ ?��\N�<ט�$K�w��u�o�UE�^˙zJ��LSA��:( �����v%��ΰ�J��:�Ƽ�o���斩H�R���r�����ƸVNj�9M,w*���Z�&¿/{�XO>r�V�0�D��϶BU4��-���k~BC�Au+��.ҵ��vg�d�*p*�K��g���}���qd^D_i��O�o'����ϯi]<��!g,�o�%)������K��Xm`��������$M1�#�K9�m����ݭ	j�b\y>�C�d�[?K�ЁuB���>/�,�i��6�����p#�yR"|�&�XKhv�TX�g۱��>.�ʹ�
=��7oȗ�'�Xm^<c�P��`̵�1̼~�Y'���lW�a eĤ4~�@]��'�$E޷iT6�5,ͻ�1��>aa�k^4�FA?���7=����$0)���?RNY(��M.�������c ���y��]Zo�n��EQ	�����o���R��GMɐx�ԓ+�//�>�u9n&�E>UY ��Ӑ!�5ڰ���K�����sA�R���8b��v-��43��gB��s����]?El;j����H4PƆ6+Kz�QV�ؾ�]q�gC���t�CJv���^ ��>w��������7m�rx���9����?S��_��.���<��P���1n�?����Z���n�m/E�⊪�W|G�u�xhP�����k�@�	[:ϯ5�`Pǀ��?�d��~D`�f��t*�������x�����X&��]PS�)q\��HZ ŏV�7&X���Ht����7{�c�:덒E�ܨe���/��QC[�j~_��!0��vz��J7�gB_[m8q�%�����^64^hIe�:��B�B'������-��,�� ��Wf�$�u9�ܛ�K��*d8~F"�F�5�&K����/^;��։�!Ǵ����<��D�(&�Ul}�ve�1g���R���=�Ϛ�V�?�,r���p��k� �'�zS˻��G�jNp2�? ��o���#��;Έ�X���L�����[�َ�Q�>LQ�{�	����њ��%�Ϳq������m��
]��X����Z�E�&����3�<y(1�^��a�k���)=]d$�6OA��|:9�=�	��C�r�d9�\�Ӗ��;k�F��k�'�h�JX4J���=�'>0�D�d�#(�A]�`X�޿֍��n��R;K��h֏^�7�� ��~J	}6���ǁ(Dzs'Ǌ`�"oRsR$�H�+�IɌm�+�czjt2�E��\�.��ۍgQT�+��{û�$�nLS��|0i�k��]C|6�8L��v��fA15��XL�Jr'�K��KQ�1Y%P(��a��P���wuB)�QV �dWzȞ>�߮۾�M��h�#]���bvҒq���&��{k�����)ڒ���X �6H����Q$��⿹�3)�/ ��

(u��e���@|�Mc��<�����Ϫ��7�0g ���3�L/t(�C�m#B�X���h��S|o;=HA��3���^�z���4��.��C7Y�����OCP.�
��p�45Q���8Yd<l��yh� Qh(�&;�D�9��C�F�q�bI�D�!2I(�~�J�z5;�U�0��|����ǈ���;P����Ϩd���?�)o��ޫ�R��8���p/]H/�5��6��O�I{	W޳�Fk2�OAh-M��P�&���%W��;�NvGN�B�|������GX���5��Ѩ"gJy��nVӣ�
�Y� �E��Bb�����i��[F��	K�+Bb�bՑ@��
���TI��te�0��$]t�p0^c�� /�$P�VUV&m��H��̕��'��3��/5��yZ~N"�Mє�jQe@F�],��v��t�e�,�
���pe���N�R�R!�ƫL�\����i�	���1\'�/�m�M�M$l�����Q�/��_�B"��K0�O�P�Z�+S��E`��)�Ȥ����Ie�"2��qc�bЄ��^'g�[�~�"s����0S�d� 4�${�K"K�o[Gh�I�_�i_�y�{V��cx���R�R����@��k/T�� ���<�$�<��6�UW������z����5_RӊJ���`�Q:�Θ��;�|���t�e�P6�w �.:��'�B��'�J��:� ��@����ҿ�r���2���̓��*���/��+�ss#E(���U��1�E�=Ag���F�u�D�1/�|�Gk1�l_�h��3ib�מ�>�m5�͕s�Em�K��KyLk]h���}��(QKb`[<K)j���m�m͵�N�[��l�&FK�ou�0���9k{��A�M��i���Nd+>�(n����Fl�}�0{�"��VCX�N�ۙ�" :��VOi�l�^o�O��^QOTm��"���L��r�Q7C�K�!��K}�A$2r\���U� ꤣU�؞E��0}ԗb�S�邽��2����'P �>���d�K���x����O%��R��:|���E]̡�~��I}�st��]��L�H�l:�#^<ϯ��30>��cl �+�<���K�h���}i�]W���{��cʓ8�o�.�|��y	�5R�{���i���d��H.[8�]� T�w��xx��^^Olq��z5��!4
	H!��R���͔+��j��]��=��쑞U�ap���d�#"N`î�$o�bk/�f�r������y<�B5oj^�*�0Zɖ���ý��5Kc��A^!�z������ �g/M��	#�s�/Ȉ��o��A'?�J5�W�$: !��s� ���M}��0��1u)��J�C��J̑��|AC��0�[�`}e��z���+�=��u���M�6B�i���ۖ�E%W^�dp�8�?#r�p'�z|���m�IS�)djZ,�pu�����v�	��l�㏩�=t��C{����/<:0�{��B��1��ћ���m��wV��%���<+Mn��O�)��j뇻�l��"�J�+er������\�yp�!�-�dD�g}��7o�t-�		��QT�.M�3��I���$A������N9�QFX�F�zLhI�;�+���Pr��)4/}���3rp�ePY�}pdh����hj����\��/e[{�#��ʁ���b��-�+,��F��d3I��WK���N<N�����:���SZeM �M�qꛑ�\��Kf�s�lJ�[���F��RmU�(qX���/_�Q�l�V9�o��YCSR�	�
*m����1�����1�^L��+$S�Az	��-Iy��?��H�M�tL�p���r� �n����,�0ёB�f
�����d맼�ˬ?f�)�����O��Fڣ��Dp��L@��R����O*J?W{`L��Zq�9�ݸ�]����{F�Bp�l�� ����������$�"��_u��?ħ���Þ�W9��"�껟����ƴC�*?<'��5�=��y�I?1G�]��k~���E93�󦓆��!Q���-�a3�6��x�D2�p�V�<E��ܡN��8
Z��ڪ;W��D���	�/ܰ��Y�SH{�X/�6�lc ���p�Nؘ�|Թ�AH┐ӂ�S}�kU���E^t�J��M�wF��.�2�y�;G��c0�A8ҳ�<jF�r�^��d�Q�`ܽ 銟��4B)����\;�((�����;'��w�xVK�cC��x*m���\��U0�ji�a���`]^��@��fدV]δ�ώ�צ��O��Q��AE�Ef~����p���1�J+*�N�y�o��z.A �m��6�r��R1	=�����c��r%:��ͩȨ���h��T�Y
sOe������oP����נG澧aEۖ Sx�r�0�¶���P�.�ڝ� �� ���U���?��A��|�	�w���ʎ�-ǋ�jF @�%9<�5?���$�Β��B^��2Փ/#f_��~�{!
bl�ա�O�����/r���4G@��m�Ku�����REƞ/��70,tD���w��H�����A��z�OT�g\kض�x��\��sq���YT�3nq:�+�Q�؊���e�,�y�_� �%eF�>��	���;D�O�O������\�C�$�V�n����n�pu�$�ޕ-Rc���
�<1�:���I�=��t`T�E2�bW��C(%�,4Ay����/p,MMqr[�����P@��k��:�A:!S^�|AB�<��rWF"4�a�0WSێ���K�=mƫ�F����=�Av$Z����\��T��Φrf�;	����g)G���fY`��������R�ԛe_��W�
ՠ0�c��nj����e��/%��Ǎ�����a�2K����R��vc7��a�F	��d�|�S=�*��槽�k1�9N�f�f���WaSiL)��i�0ϵ���N��Og��bZ7��|�vK���mq$&��5N�椣�ND��/�6���}��-6��� ���x�m�7g��R�����uRH_��)*�H���H)�+GX�������7TmNVv�v���v[4X~�jbr��8�/�Y?l�sK7�иPw��㔍����J>���Ȟ��X�U���<�8LVyjYcm�z�+/�-k�4~Hz�@+���qL������{�
������e�&H��8#�]����\$��yK�h/�x�O��(8�E��I���`Gd��Z�G�V�g�Tb�>���Wb��y��x0U�J:�09�l���| ���7��zwo��6V*���X��:��B< w������\j	�N|QY��;w��1���#v�Q6�*��m���@�Y�=�d���O&f��E��A���Z6���Y"Z��BIFx� �A���v�h������Sɲy�7�-W0��6X��j]:7 }��t��2_M���8�{Q�l��E�yQU\�vh������_���9��,��WU+��v���_�iLbՊ��{�ޯ�!&���Ai�	5�`e�:����H�s�4����I�/JV!AlyxT�Nf�B�5�,�W��!B8���"ak���#��v��<����qs1��Q4'PV�O�����.,���n�L���/$D5�
k�n��������O�C���MJ�N�#�mm��>�4�R^F}�)bw�p����[�A����� .���;�'�پm���a2RA�&%=��|�#$$���C�sn
�_1�R�%��=ўܮ��* �6���s��E㌰���������f��y������
Z�����鬢f_�����UMk��-��F���+?�D���'V���Q�@�:;ܙ�c���1y�qBu F�v�䫿�'�UNvu�֧�� �V	��i:��&u(,{'ZCY���OR�m5#��͈"��me�cx�^Q���F��v|w!BVL����³S�p��Ү�6�B<Z���|p�S�ZIԈ�t�S�\��x��H�6���I�tBJ��(sϙ���R�v�k��6z�Nɉ��DZ9R����=��?��#k���9Ղ_V����W K�M�Wk]o��;���Ռ^qiv��Ccv�.�?2�=6CP驐��imb�@MCc��(�/�+�ҋ]��{{��Ͻ�D��$p���������h$S��p��8-��K�~N��,�2O�s��^�=��F��z�h����	ӯ�I�,M����0���Jp���`��Z\#c�դ����S�;��b&��5 �F�K���<B(2U���YJv҇�M�Ϻ5q���]<ۀ�c����&�~խ@w�;����O��<
l\�����򪥢�����4�ߎՃ�I�{�oQ�&��e������<�":y��3����+X$�2�&�$�@�����#���^��/?�hb��(��/����ǭ���Y��� T�<�X�JIyHv4�mLM"b��۠���mP����5s#EJ�\����i��˯���lV9W��l3di.���6?��/�"E�\�[�b��B�G|�c��v*-��Ԥ~���0���=G�>����N��	.��U�iR�;��ŉ�Bń	"�k��B#�'�h:<�	�x4��+��}*����y�-h7���?M��Y����^�Q1 ��	���+s�${����=}�J�u�}0��@��>�nT���U̠V�:�?��(da��d�,��btyi�h�k><�1�<��QVk�L���I���:�h?Y �����H=��/�i���B�����/s����3��$���6���lZ��q7'��*:�����_���2��x�.�*�8{O$muQtLv�l��(��M�0�.=�#(
��Ѐ�0#}�0���#g��7rF$��P�����<��6��=�uL��*^��[�gw�%F1�q�%��~@^���*,�FNߍ`>q��V×�r�ѐ�K�L�Y-|���d
�_0�3�e?�~�d�L�ͫ����o�ג��:��:�R.���-[�иmk�@v�]��{�E���L���W��8[;V|Ap�T�w_�o+�� �m���C�
@ّ�R��A�NQa���ʹb^3�ܒ�Av�xޑ�L-����
O%r�6���v���������a��N*���J0�E��6r�zC�q�]Nڤ��N��5\���h�.�c���ؠޅ���N��Y���;Mr1�ˮ��qh-]�8��Tm��^�?w��㕁ud��~�S<�=��:\;�7c�C�󟲨ް�m��V�,pt��]����JU� �����+F=���=/�V?�3ªh���|���Y�d�e�wن����ľ�i>ibvRs�EfD����b�Ə��cm,�֢�x���{�2�p����Y�)��7��<����)�}0���yr�fv9ab��M�<j��a4��L��-�V(	������Y*}��+��l�ȿPRJ�|_U!��8~�y�rv��	Kt喌Ϲk%X��\�M0��Y��W����Q��t�Y��[�����_?�Q"��D�n��>����T�,@u���g19�ɞ-0p$ZSz1��\��>t`k�v�rW6C�-Yf�i�̀Q��C���S�!�8��G�*0����hZ�|�ԓ[(�'{�
 �����9�����^:�d�C<��D�|��"����K�4��t�i�x15��a岝��Ǔiy"�X����⚪��I�Wq��T2)i}�������v�f�l!����7J��`�2�n��{;���!�