��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#��gߑ�2�E����hy���a=��cy���mou�4�L�R���:�ZM��'c��_�T,S���w��6�r�u��%2�p�R��+tR$��W'>���K$B�-�"�א�d�H�4׶kZ�OC,Y����	b��32S)��ޡD^l��V�ߐfhʣ�I�X���lH��\��Q��؏�(;�����˳���H����f�bţ��[�W��+�I�"|���� ��15�!��u�A:w��N��g�s����v��-�e%F��L�/��8�d�6 p���7Fj��`ȧ׭��Go��[à��m�T ~��ϗ��M��D"Dws�'�ބR�D�S�Yz�-�ͣ	"v�Y���@��7��r�a���k�p�ɜy�Ir$����L�瞍<\~'dl�V$�v��T-k3U$�7�A������c�jٿ�0��J5|��8�=����qtc�E�E8��!nq}�i�Y)Z��*:;��j�h���8�H�C�ae�Z,=T���rw�e�d.���S4)%|�����!�4�RN�>����)��9!��u��z;�5�|ޕXk�V5��/�E�s��J�F�Z���7\���R���|B󵳨j�߻�Ip��s6�/MQE�GP��ʣ� ��	�$:rMZa��	�W���lk�q~�](�������VB�RP��C�c�奬ݹ�[ьP��q:��N5�gg�r��ν�EdK��'_��W:�|�:��d�=h�x^Pz�p���,�
�&�}I!�#����/Y% ���Ǆ��B��E��#�R� ��?��> t�#���(@�.�س!������Xh�O��2��;P���* �cH2$n�[Z�`��mB4�c�5,�V�`|EY�z���w���ܻQok�M��<}��7(��7ϫh�ǡ��]���w2������N�T�,�9��c:�\�C�솇�C-2��b?�G�*�_����{���q@�V��HF"	���\�)b�H�Z?��M��p{�%5ޅ��yv�Eu���ڦ ��1.@�q��t=�|�Z��*맜��p
��&�ӹե��Ϭ����_�	��?(�|¡~柋�E>+�֒!	���j2����en�k�8��@\U��,�)�����+7��yn�x+c���d����6#d�*) ���}���_�1� D �9-`���u�si�	G����;-��zAН��wDD�׎g��)�Cf��v�x�r0�_s��Y;W#�:�y�������?Q2��D̏9������In%a�}W�a�V��S5K�ςe���M����r�����h����/������Zk����idC�c��/�_JN���bL�(`2�#�I���u�@����l���q�:�h�߷�S�W�-��v�*^�����ɂd1#湀l}D�2x��E��'4K]���$���@����ƛ��hn���D�Lf� �.��a�"��צ�_ È͋�7Q���Rr��q�˼��o�k��"�d�L]�SWL[�ߝ~ǔ�}ʱ>$O�;��9�x.���6`����������MLEY�?/��|��ߩ��CO�
�jL4�޸W}f,���礤O$V C��0p��i�=��}r�cLfSK�%���L�oDlgN�d�8���i���YUJ���*�����$XL�B$�R�������9݁E��Z��W5�����
���$�B>�?�ܒ2��	����4*�*8�2��l�����������/8V�gJ��e��BO$`L5���V����D�D��ó������D�Iu���勂��B+C�g��J�w��4"w�rL{Rk0����5��<�ek�#w��C���^�Ȫ��s��/�Q4^̟,2G���2=��������p��}�������}��kr	k��F�=곩�I�Ѡ8�6�7�M�z�&9o��k��9<قZڊ�r�b�����jh:C��N¤��o���ɉȌ|H�Uv��"�����s�;��t��w��kFQO��J���0�C� �/[���u��>M
���\Ӕ&�����pr�P|��]g�eۺ�`E�LX�����n�Up��nv� أ��L)b�Ɉw�o�pw�;�eC���zcM�ڥh�N>�����w_�y��o]$�{��倇f,�o�A�Va������z\U�"0>4�:g�Eq�� :�w"�n#2��F�46d�yɻ�R���ap]���!@P5�sQ��ݧ��'��3	�D�����X��O�_8���Zm!�B��D)P(tB4$
օ�08��`��C��9@J	?��<���A���h�>y刘�b��-��|]�vVD5���n[��k��{��#ϕ+�(^&d D>�?�a���T�Г06B��w)g�����ӃH*�UH �ςC�2jӴ93��U�NmQ�� 0`��OaA��Q���������w.�RH�:p�E��>i$�#�÷'���ul��9��d}� ��~��#g(z�NED���Q��|D�Y�%�^Ep��і���.�������Q����) �uo�#��c��	F2/�����D��u4��`�G�����0eG�vbA!gE�*W��;�m��^K��G{;8��N��,�"1���J�R�=�J�j�h�?y�s<�ԬN�|��=܆%�H��:$���'SY��+�v����U�k����T7���^�2�_  o|�����Hc�~�EZVR'�e�Һ-�.O��ۃZB���Ac�������dnn��+Q(EUӏ-`� ��ô�UA��a@�jpB�<|��4`FDP�xs�'ґ.��t\xs��W����(���k�Ch��#�ݩ�=hI��Aʂ��z�EY��Ld��Ũ� ¡��3=El�콪HLǟ[�pcT��)����|+�O�$���n�b���T%9���u�+�&�Z�P�=����Z�'��RS��u[�I�����H�\�������������f)}�0lH��#��=�A9��l���R_��%Z�4;w,ҥ�f�|�訾Y���G�3_\6�5|�'�hq���>���U�ώ�Y7���J�Nk��|(���L��T�ȕg	]� ��+�K4E$Uh���:�����m�/N����'^����0#� '�N=aOb7�A/�;�����z�a����T�a`�k�A�������z�yl���:�RV�����
�R	i�V�U���	�GD��5#���;d7Q](.�4�C���O D�����}��9����
�E �ģ��zqg�!�1�!#�%��&�U�1���;�\�Y�?6��7�^($�8�nl?[.i���Ҹ��pHS�y��B��c�x���U�,�vQ��-�N��<G`�������鱲�_��µ1']1�u��tQ�
�LJ�|u�
�V��q!��,R��ƞh>�;��;���fP��}���*曽�{��RsN��W~~N���Vx�Gϲ �۟�9��C�:�eAc���p��o�)>�<�Q�w5��2J�� �g���z�̂a�Ы[g0ﳣM���<�&2�a�Gm�)��O:r]����ǩ{skfA��G�;� �Z������T��#�(�)�xD
|�����V}�S|.f*k*9+e���^} �#�L��J�4�~����CB33����z��""e7<�B���\�ע�'�ҤP=bb���m?l8���u�����Z�D���쩔�W����H[�헜	��m�� ��W�Ȕ[�|m�ߘuo��P�v���(cfQ�Ѥ��e���O�d�H�k���Fv�l����^���&,	���>P��S1$��x�܃��Z8N�L����tdXs`�)O��Ry0%�꾟��q�	A��Z}�u���o��ՠ��84T��|�ΠF�^�_\��1d�N���Ѓ��:� ����Be�1Q(7�L��eռ�xh#��{p�Gr��7���"cE:0u����x {�t�:ˇ���w�gJ(i�*���T�E}� �������F����p�*��+;�h���鲕j
��E���0��$�1����]�U{�j��_��ʎ��k"rXFos��#�q��J̺~����s�sv�*[<�a�
��M��U���s��@��r� ����6�^W�-�6��9�B��p� q��w�m��Nt�1P@u�� �4SLy�)�Gq3 ����T���)��F#���\/�CX�?�:y2!����$4W��!�������cɬ(8e��;��ʇ_x�wv>��:@Q����xx�v���.�5j�r!)�R)+\�ĩ~�� $ߓL���[������s���}6G�qA��F!D)��q2u;�+�loU�"IU�B����T7�j��*l�Fjm\�e�����J��<�pb��@t<�f���Ծ���~V�$�Y���Z�A'�U�7fo!IE�T�_\��mP㗆��z����"�f��Z�5�A��8�R��ј���C�����A[�5<OG�쏮�H�R�5�F�������A#L<W@e�R��D�_�2�[�����`7��@ro�[>*�;��5!֑(C���>���� �Z¼id�9��/�F�;^�b�֊��>V2?E��D��������V.��Q����h��Jr4��A�_����Tm�	�&ɺ���m6Z:�'}6�=��qz��/�t�_)���$Z]I\�w�]���D�x�Brm�f�k�4d��ϝ��~��бO;}#�;&�w|#��=����k�t�z�4&��B��)"\!�i��q-")�֜f�=����� &	�^v7t���J�%.�!hY�V{<e��OW�t�W�l���:��sI7�Kp����j�)݋@̝�x�bg��J�[��v��:@����c���Jc��2&t����א	���0bG��*������y�#h}�Я�_c0!��e!ؐ���G�O
2\r8?�����ZA����?�Y8����=Xs�6d�߶����� ;��R>b�I��|#x@_��Ӻ���>��O�����N��_� B��F��P݈x�S����էP��Ze�Ґ���TL5��Ճ���?F���������N��4�V�- >���@Ā���8Dp?mYN�>�W#����$x��+C�	Ϗ\Hd(�F7NN�|)+ܨ}�`�^�=#D�5^D��<��i�]�z[j$C��� ��Wx��2O���p�.LYM��2��z� k
?�U�d)(��ӫ�Sw����J���꜅	�6Pvrzk!Λ4�O���
�@�������lذ?݄M�tz��~+[����O�q�2���{�"8�"$�#��@�7��q��� dۦ6�>Dy�_>��{�8�P�b�=����@w�j8���S.|�5����F  �j�7���`l�Y�{RRی�.4�k?����\���-C��mT#hJ��*v�/S�h����An#s糱�E�ЩH����)�ns��n�=;X���N�<�-s\��n�DS'S[w�=�	�S)�xDʊ�&�_�? t���\C��l��f��/�w�xE�7���+�-i��x�7��:��'�$��OW!<aj���S�����;�۠-�Kō�i3u�䔫�B[�H:�79gW�������|w��H<L2��s���Z&�%g��F�'*�G�ո�������_?)y�i��2��Pp�����j�.~��f�'�|���%eo�#�a�f�kA#Po�j�&q��L���p{'J�㰏�h~�xeM3��B"��p'��w[�vuR
y��� ��=�zT��*�3&�B��|"� tZ�,?��<���I�����|��f�ϦE&��,\e����a�R��Cƻ��1;��_ܥ��Y�v#u��+j���Ek��-!~�3��4w&�H�U/�}6���5��.�Cy��;Ok1�.����@É6g���Է-;��h^��YLV��
��sRP�bp�,�4�	�ά����$X�W�od}� ao�|[1���Q�̢4�G�2�{dʭz�a�$g6\�x����h
/�VB�gx5�a�G|��=�B���g� s�"/�q�;�.�m<���G�Ʉ�V
x��Y>�.߳G�Qm�#sGKny�(�y	���9��u��;��o#�[������`:���|i�� 6vQ���s���^'K��JlV����ī@��(�X#ܣ�5d�7��>�eX �Vi�~�*�����hq���Kn�^�1!�X�x�l��?��WE�t���JZ��8����~�`�������,�i�.8��V��g��z�u��Pε`@���]㴔
*�6��eG~E����uNuW+�ޥ��uJ�z[��0�`B:�Dj�V�.OJ������T�ȯ�{)ya0���+�^�'�~�Y�q��%����.�_9_�@���j0l�L�rmC�~Ltb1PBe�8������޷B����ֈ��wMm�y�
 ��C ��_��YK����`�՚G�g:��u)�+nPi��纙��w�M�2MzP��r�Ϩy�7�pW�b9^�E�8���Q�_�}�|����g��ͰF��H#�P_���P���`��t�ҭ�1�Jw5i�2�k�վ��h��融�C&Nn�TuG�����i,�����>�m�'�ٝ�9����W���J��#���I�99�L.�V�  "�?MK�1��Z7�0&�	orA�$��)T�8eR���ڃ���@-�ahǥ��"D�ȝ��8�SR2�
�gK[��6��[*�5N�¿�ⷷ;�$�I�q��R����M�}�9����TV�8z��ͣD�%��S��n�� ^q=���+��0�)}^��b��aQ/���4����=�-�_������HKՓ��T�F]�K!u>L����Ph-�.ص��	R��P��{�'(<�����5�Bj0��{&.'ip`E�����GqH��^�xa��Q�'#U�CH1��������u#�T��� E�ɣ�R[3¬f��z��h)�[��5x�Mm,�e�>@=4�m���hb�����eX����G0��[b��0~�fS�D�/W�	�J��U`B�?�𴀝dn�흩�Du@3��%����$�F���HIm _x�����"e�L�;Yx�D@���c�!/YH(��v�cĒ�
�l� �7u�����E}]{o�O:5R�f�rѥ8T�<>s:~�4 9}����e��?�8��o>Z���ϲl� ��.?md�IA;ޟ��ާ���tˆI�r����M����1��n�H��<�y?V0���ȩ5r��(ð� y�B�Vl�"�O�A�Zy�c�*��p4k�ȯЯhx��{�
P�D۱&-��q�l���ؘ��Lz�(
$�d���5�U��t�J�p쳢#���X��;7���N�E�>��;��KO_<.-�!|�|R�5ټ|w�*��-O0o>;p}ӷ�����w-m�Ͷ��]���a�����	�����j�M��Z��������ޙo��W��s�ذ�-� ��8�����A��㗧�Wv�j{3���er�5����ί�ޭ,a���K��	˵E"�^^^�d�n��[4���v�);��a��W���$Z�n�9$pS�+B�.��������
���t��H�E��ҿ�n�L�;�#J�πc��I�Q�(K[�1�8z*q�s��Z�+�O�xH������l�S�~�]K�O��f�lsMOi�����WS�����%�^�WW���&��a2��)�)B��E糺MHK�M�~i.��@�qܞ�=>A'���K#��(Z[�	TpJ����G]}�������Ї#/)�G���LԳ�_�R�B|je@�ߊé9��Ը�S:��%�f1+^)c�k�t�푸��BgQ[���,,�5�>XE�����j�n��{
Ջ�#y/ϸ��羆�_�ȩ�o88ˁNg�B�$���������m�����T<���v	�܀i��g%�8P�oؕ�8/�D=Q��M5�F1�������l�S�RlI�M��^^q�Ȥ�V�@郷��i���?II�cϣ3���D��@�	v�GXZ}��
	���!Cq�&��]���'���y�����+��� q��+��v�TEc�!;�Pw�|�,�+Mښs2u`���l:��+Я%M/� ����F�L?U<L����V��3�Uد�V�nj��|���܍n�A����v�6�<R�kP�^;"�Q�}@�d"�jFG�e8Ŕ�p>��NuCd:�GNN�o�,'��B�B+��	�aPm��@:J���Ǭ��� m���V(�H�u�=��P4�SȻ������@�ҤM��A�����>��z5eb�����K{��Sxd1."��ѩ����m�J�9�X�˥?�O>��Ŋ���t������6�En2:�L�����t��9�I��ȁԁ�(�ؒ0S���.�,������'xv������8&0f|5eWnz���C$	/Y�H���1�R��B�sʃ}tM��*�������"������Qjt��Y�[�g�������
�=�n�[Q����q2�#r���脇�����/�O�9fy��lyS/�x��{�1���L��ѥ,�����'a�J�}��fKx��Ek�y��Y>J��ƚ"��}�B���w�m�uh0�9�
����ׯZ�I�җ�I|�Y�K=I����S�O'���:\�v9��=�F#{\Fu�!R,�����"˲+��&��g_+��M�jt=~(!Q�QO�r��Q�RJ�č��l8�.*u#��J�U@�^oGL��Q{�D)s��L�)��S*��E�����01��#1�Gw�OTM�8R��Yt��#�5�v*|ad�8iY����2^�Q�!�sQ���lX~ڙvQ����a.&L�h��{ĸ���L&�P����l��ϐ��M!j�V����t�XO7�*�M�Fz8��MVBR�~���A�́�WV|�.7m��*������&�ٝ�='��q]�z��A���^HFD�~b�DT�{O:�š�MCW��ݕ�zn$0o�Ozz��ޡ]ڪ�����x0EP!�X_�e<�����*��m8Y`�_�q�li�pF��]�z����V����W�#�8��CI�h�Up�����Z��I���d�G$�N&��Y��5}�������F�������=c��r@��ߙ"��g�CD�(1%�ޠ�l��� l��e���Z������.���"��ep�8����e��<���$wB�^l�'�^�0%�z�9q���v���q\����!�\�L)"�������Z��V[�$0�^k�<@��4mA�4��JB��,��-�-�-��4�b��ܴP�����n�(G��
,�x����	�p	kG��H:�a(Ff5B~��[q��C/}�6o�8�lw���28���Vw��Ȳ������/ǒ��D�!\b*Ve>��I�'%t�e�N�g&r�N<��WJH:�������F6�V�?���hisٸ�"W;��@����Ԗ���7�x�m��)��\|���t�S����8ft�h��v�ʈ�p&�8Z�\���E�V�� ���f&�CB��`F�#ߙ���i
�O]���A����� 1�0��V�L*�n��O���� �y֒�YD'��Y.*\�L7�I�r�s��kZw�@��8.�}�\���ĳe�.H3p�)�cq�taoJ��f�yϖVCf�<��$l�����tm��:Y8���Ҳ/�N[��Yy~�x�C��[����
�ٴ�`*�eT~e�:�~ǍrP=I��%�Q���;�A���D7wP>��*Έ
6��Z�d�}W���>b��"twX��D�AQmIp��o,G�S?9M�Jɇ��E��c���ձCAݠ?��<a��������Y[�Zt��l��N����Fu\��ǣ9xH�p7+�Y�u"6�¡W��xa��\ ��쎹�|:/��7�0;�`=�զu"4d�