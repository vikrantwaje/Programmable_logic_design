��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#����)�`�7_��H1F����%��]��Y�zt�o	�x�Ĥ=M����X0�����������#�lwZZJ/y��b3��!�Yy�J��[��Ŭ���� ס^dR ����*O�
aG��~B��d���Вvj#^��wP�K�LK��*�d~N�垑U��/f ��&�� ẕ�|�BQٓ��;�d��Y��Z|���;lDYqi�\QLw+�����6|�zl�����Y�d�:�N7Q�|�(���[ٴ�k�9 �y�����V�j��ʃ�`�s��2� [|h��Y�!4��*�x���/'���p���B���&h�>P��f�䠎G"��6l��h(T">@� @��B}��ם{�@9����qS�^�T_�/oڟ�)�@���U3æJ�jm�0~1�Ԝ��"t��m������[~(���K��W>�j|�����Q7��[���ｻ�)�	
��d�4��k*n�p�iss�W� tt�.�l�
̎�TY���m�A��!�����/y��	D�C�w(I�^�x���/��%�ڮ��9�~��!Q�G#�d��ZA�i���v���բ�J0�`f`�� �)�-����P@���|x��"��W����HI�&
�G�y�N/x��c����SJV�w�X�vl���,�2m��W�rn郙��(GV̢;H���d���@�<��c_ #/~,[���|d��ߍ�.�t|	�q�V��6�Q���D�o�	&m���yి&�g������͵Ѕ�E�ߟ嫔͍����a��n.� �R_������Jy������X-�
K�[��;E�	���E�ہ��S|�7|�<2j��~��g�ȄmO���#�1�H�����q�G~��.Aw\��)�f�]z����&0��:��l�,7�Z�ր�o���1���&[�)樄b��s���S�,�!���	�Vrݷi��L��h�DiJ�p�S��i�� ~l�7[�v���`DwTkz�����G_&�D׈0�����P�G궶������/��3��p������/�n;�m+?�s^�T�d3��jU2����oI����U4���&�r����O�\E�>���?�]�I3�_9X���iV��m�/K C2
��+P�� :���{c�A�M�""��r��m�Y��R5r�Fp�+��Z�ï�	��ЎOD�a� Wja@;Te�o�>�;?B#�v6�ĸ��-@N�x�	��
m'u�\7��ש�f�Hv������l��@���g7�E�:[�	R�S���T�R��pC~�p���I�ת��2��P9G�.�!hpaɹ2`:	66/sE�����Ձ+��7ޠ�]���A���+�h��`	�ٱ��ќ��Ygr���:�";�����iNU��+��L	g���d.m������Bb�&y'��j�"�{�G$7
��꽔x#x�Fm#�PSA{o���l�ǭ���=����-��o��Z�b7o��~�+���+"-�F ��%4�v�I����]>�WP��H>��	x<�氢L*�N a�^��W�.e��Z�=~)��6�I3�$�Y�h3����D�Y�'�ק�9Vg���L@��P��)�@洜�����r��|ư&��\��6��U��M�~0��������I[���Z��yg�Upy�b��� �a��%�����543c�Z���+$�UIf<�a�=�j�:�}���gV�����(ƛ����#p!$�}$��4@�h゚�8�78^��;�����#{�{3�Ѿ^������ph�Eѽ���y���̲G�`���_���Dt��������ݬ�P��ߠ>��]V�04���u��+Egw�8��1 ��(T��1����V3�(s��K?ʄ�;_)3�&��>�M���W"�5��\C�O+ԶR+����ʂD��[�;��������1��p�O�Q�3�=l�ݚ�9� g�m۩��T�H,~���\���a01	=��4��4|�grE�x�.R��j1�<���0Z5�C����g��&���P�����M�fX,F��
d�6֕ȣps�D ��,��D�c��W����-n�
.��Y��J�����I�������Hͷ�>���I���!譼Z8Ͽ���.��H�z�q�봝���3�e6E�}��>����!]}hW�CG˝��w�t�hrh����&M]٢�Em�h�.�(G��#�?5��.��s�Z��W�;D�J5R��%����� =L�\�n��r��t_e5��dL� �J4{0M,t0]l�ˣ�}3������n�[B 4�	X;f�$�K�I[ܞ���>����]Ԃ,�:��VA�2�y2:�z��?!���|�[���)���א���A>�E�Wd���o߰�(I�V�N�EsT(>�|���f'�-�gj�F>��`;�	:���9�	��vxX�MYD�+f������ur��􋜈��w-"&��+BM���ωs���;dg��yK.�ÄU�H�D,\�E�]aV;�dn� |��v	�"�cjG�M���-�����X�eF:���80ً�Oj:yIv��K�7)��,��y1z_Þ�n?Z�(�/�L��(�eF=�Z�{[�q�
}���X12N��e�L;��5H���M���CN��j���afAf�Y�#��g*�J������6�n�cO'�	Q����?S�?O��(="z�"�g.=8�b�K+�ҁ҂;�b�y�B8�w������)@�C&������GM��b�T��(�ZɞN�����ԋ�)j�~��O(�(3��{�%D��T�����L�Ț����o�\�5�5��&�1�X�e&�y�Hr��-���?��i-ۓ�>���4�u'5ʣ�";��9��!�ǎ�5}�#+?~j��u��s�����2-�Ys̳t�����'�#}��W t���bT,��ڙ��n�37�� {F^��~�A��JOy��gI����o���G��˜A�힛9K��HȒs��p��� m��seRv���!��ۗ��mh�r�Ӣ`L1�J��\N�R~��s�Ç��+���m���\�#���6��J6��sĹb��G�U�|��)�7��ջ��Wn]#�H-�G�^-��0�ǀ$
���|f�Nh@NE9®�_>��	�E��k�
�I�ܝ�	�x�YS�E��%�2�&*l�rJ��u�B���ơ Uj�k�������b����!c����͌��ߊzJ)��$X�H��qbV�D:�,*B$��z���R`�� D��N븀��@'����+D��Q�E��"����ap�x���>����_@\��T���Q)A$5J)6��pX(�kE_8�\���&�,�p�AdEfv���c��Ǧ|���;e�&��P��>��n��4V�fD���v��nw�����5&�����(�5�M����;��e��`/Z}K*1g���'����+�ZP�>f�07��h"�O��)�J�>U(��$�K�=ek�����B���s����,��Vv{@�����gksS��	��h�Q�t��:�F��7�^{'F�x�#Z[�P��/3zT�+��t'�p�Mǭ�%��C��C;"�ۏ�S��7�;��!�E�S�)36w�<�����a�7��F؎9�K�Kv^�H_�ڐ"BY�S
-���Y��E�h�6�@\��QTQ����(�!c¬ eRs����y��w6��۲���)I]l-�WmE���78qCA���[�O|	��F��w���7��ƾly+�)(���zK�:m���8� �����+v��=x�ʪd��V���p�`9�-�u}�Yݰ����lY�j�"#E�g��d`>�H�R�Sl�*um�m�O�N�^�}�D��{(�P�4��xjy� ���<��|����^C�W�/æ��U�@����^l�	��`G�."nB�����TA i�8�8�f�@��/^�<Sc5d=�\�?�\9?|_�w�s���w"�k�:*մ�M�vĿ��J�&C��]��k�E���@�'�ٱ�-����;�ٴI4��H�F�E�P9�%�S��|%B1���H=�HC�*����4�Y/�<�L��1t�J���2���RQ����ī��M�~�/�ۖ���_�����\���)ҵ_N��g���"l3�d��F�mK��S����mol���i�i����&h���3���yx�]X�%2�!'şƔ��a� ��ʄ$�^
k&{��J����zu����ѼJX9�o���[�D�,:�p�|����jc*�FC��3�ZJJ���^�Ww!;2��@H��Y�,�޽�'FgZ2'��z�ƒ2�0��A�
/凙������t�L�"�'� 6X�qs�GQ�k�NY��S�� F1C%w�B�-�� �$��+�� �f����O�;EA�	�B�=�X�1
��G�m/��9}1�t�"�?
 "q��˂p4�Y�1�z��Ā9�5���hH��KcQS�a�]�v���y����|�M�l�X�x���Of���m9�u�(��.��4��9� O�i�u)g;vG�Q��?T	��|h�p������u3g?�@/��̰jo��b=p�Y�����
�|�.Q���Цi)�y�L �F���7�\+N��Ư��h[K�D�m�6�� kљ��%.:�9���G��v4��U��������sj\���.�@��5���-4��#�bH�/d����S��$�"�v9w��v�p��{�S�p���+��(�♧Y����t^��S5[��Z�3�΍c�x���3�E}�=Z��I�g-�3�s���N���-�$G�s����C����-F��A��=r���1P��0�������6�O��8t����/�ǫ�d{T�C�E�������&����6����s||�9M����TQ��$N�O���[7b{3-��@��z!�i!rR+�/�@�<u�6T,�h�M'ʜŔQ������zޚ�:��YW���`����0|Y[��x�6�&��8���}��S+�#�9���q�[�ӕ����Ih�{��+��Sܮ���h�&-�;�	��w9���]\Ӿ�����T1G��0�����Eݳ���.>hUf)�� ��F9�Į��$akuy!����Y�:su�$�d��I~}�"¯ U����'V��Ց}l�}�!i�si6��<[�z�d�oħu"5Z5ı��O�i�6;�]qP���Go��3���h	���E��s�c�?���'�S�\�٬g*׎��	������gU�сX���q�%%*&v���l,��$�p_F���?�I��{����j�N�+V�d wl�Wb_�UW����8C䋗���&Ȓ(d,#}w�����-=q�;k�Dϛi�}�,o�(3����G/g V� |g?Z�͈e�:z��5�?��M�x���%/g.wï`�g�� ��Ɵ���Y�za~�sO��N���E������}�hy�I���:�0T ���]�/��&�)|�w??bۍ~���U���C�)�~�AƐ��_^Zm�oz�Xi�"��E��5�󺚕�>~������w��U�;',� P���'�~��}�|��k�4d���x���K5pU<�]��! 7cO��ٺ���Y8t@���(�̲q'�9������s��T2��zL�$п��T(k5#�V�]��������{���2�:�V�->CY�:�7XȮF@+1S��϶r���G LX9���6�C%7X1evl�l�
(�"DQ����eCܮbwyr"�]5��5�!Nv�4�${c\�M�%ݞcA7�B�����fa��L���˔ik��2��:�%�^#�m��)}�S�A<���J!�]�����G�+7O�N�*����#��`��2[�J��z��LN���gQ���+6� ����䢅�<v��&1�Mxn���/�o@�hϺ*��p�d�`�,G�Y�o����0�<��^K�c�*�f~��.��Fr�{	S���Y�e�D���>�5t�=b��^�"�Pcܸ��H,�V���d�ٍ2���VXn~#��T4�9\�L`�0w�U(��$�g���fU q��R}iK�l���CQC2Ė��˿w����m�Z��J��A�*��k���E�+H�y���-�O�6Ҁ��7�z�
�Pk��X�����MAw�m�ϵ@���jf�:s�lj�0܎�N����,�x�7c�g�(*L��(
X��e��ul���8�FE0T�����:ȯ&�m0ux1�Ց�Ω�j��� ñ���?���z��������|� �|��{�cػ����