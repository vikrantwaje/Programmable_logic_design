��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞���Q����90�mU� ���d�ܻ�x�;�-(s�E�^}�-!^��Q3�$���i�x�V���.1��j	iC��ȹ!�͊���;�4�1qИq��S��~�y�:�����BI�F
D������.�H����/Ls�&!えky(�o�go$ˑ�G�ү'����� ��G*IHA�{�Pv�	�@��7�/���B�H��X#�ژy��7���Kրiv���
��j:�^�W�������ҥ}�P�~���ͶF�*UO��,F���iQdY�'f���F�̡��Rv���,�;%|C�t���������������g�nim�;P��R�^l N$Qq���;�jw��g���H�K�._�bB�:8�BHD ���(�w�{�A��@�3��빠����D�˿�؅�/}���7�&IkZ��xw �8dԦbq�������$6�I-���ǫ"Z?"�kS��ܞ4V���\���/�L����1���|=�[��_��C�(n�e����iퟦ�'���(^�pʪ�G��������J۔G�ϛ�b��� $�	C��N��g�V@��*z[�4�a�/�ʼ#	-�ѝL�oy���`6�ٶ��'z�pQD���
}�Zw� 2TH����'��]&t�����v�}4Z�
%�*��Cc��N}SIL���"��6����;�M�"'�f]!R�ʸ�PT�Uc��3�ȩc>����{�Loʕ�Z�V��������H ^��K�����Tl�i���=�5 ��^���t�]�qе�=�4	쎷�)-��|�Fr�A4/�ܖ�eT���!��ئ�Ջ�/�tґ�)�D���]�#��n���ӅA�!�dB��\Rv��ޒ���PzD�8E\Z��պ��{u4?��b�Ԥ�.���/��O2���Q�yq%.�	I�t>`?i��A94gz���N�PY�~fd�l`�a[�Ì��6��5���C�OQ.c�
�"!|G�K���c�.���z<K���#A����W���� �`ʊB8d#�{���"oa@��)���=��E�,��|'�i�^�\�q?E^�FV�=�1A��S8�<�vh�X�Q�9�Dh��h~��N����@�XW�+��FKqf�"�f(����\�ă~G�h���H���; ���9�2��O��&�%~Я#��a�ig�|��M��r�?�(Nh��q�չ��`Q�Чd��
-����� �"񎹐\�nҥޢ��NC�槁 =g<��>*oܮ�tx�V3�'y��5J�0y�_"�ݣ���tJ:�5�-��:arlI}�{5�Q�mW:Y��6� 3���2 �(;����]J���p��[@���,%V�����2�HuA��N��T����q
�"��8���++k��G1o[=�?���m�XW���M<�77�E�n��T2���F�W��p8w�U���/�u@\�-�K��o�����XPs�3����|�*c�f��!<���Y����H�����oA�TQ��'R��g���rD�������R-F����S����	�T��g&�cbm-��x�7տ�
ΊyAc.7�}hW.|ˊ/�����c�{�v_U?/�
�'����"�������<cPl�Ya����M�2�0�"5|S��4���	RC�g>Qʨ�A�qޭt:�S�V�޷~��@���F2ͬg�^(�Y�!��v�#���S��He�����	M3;�5{�&l0,���Y������Q3�����Yo]�� 8e���b�A�~87�E2!P�oG�j��a�.��EP�����r��V�=8)P#�2Ө�A)��4��Β���+����]
[���~��җJ���"iI6#} f)�L`���7��!4X���}f�¥j�tGI{�d�Y�(�����[�M]�PF�6�����G�d�xo� �oȸOx̲V��X�J�S���G�<mT�(m���r��QX�$�D��$�j7��L��w�2"���V���7I���a���)�Y��5}G��Ӟf���.5I2�1)�{�v�����3�$g� B2����#�L��
Q���˺�Y%���M9��"�R�|SG(�Mغ�v��*J��6�%�'��G��hT���:�	��x`~5�=`W��	���F	K{�c��r�f������c���C� ��sX`�35B�Y��'�5_Պ��7������눽4����ȓ����[U�Ĵl��:\��흾'/�+�P����P'�{ri�oV����;ׯPx�e����$cʾ�����t��F�\�$ݔ�n	�U���yjTЎ�^u<��՟BQf�����*����~�E����b��^'	V���O�l8��5"52*,b��7l�9���^��!`L ���LNU���	R��ܩ���vQI�$<VԌ��?�j���1xk���z�ͪ�?&`r׋�&��!=>Uۚ.�H�m�±-�	�9R�T9z��q|jۧ��S�?w�������ɉ�> �m��dG���Y�	�Ԡ3�`^�)yY:)�u-s9����K�1Ֆ�F�\����'��U�(	�p�5���}�
K%2����#ɯ%FL�74gr�����/�*�P��D����:U�dڻU\}V*%�Ts�௢&�-�帍��q~@S(hPک!��~T�s<�D��TH�4.��1�	o�EY"���>-MzV�������_��6�钫bn���،��R!�V\��]���������Mg/Ϫ'�&��V��y�$�t�[CjSK���T�������!~�h!�ذ�%�8 x�"��Y�K�p{�uۉ�Z�L_��@)��؄��>-�D<T����n�9��g/n%���H֫�t�\yF|�wOs�0%�t�-ܠ#���WGC���q���7<1;8�A�
��(��p�Dé$mi��]l6aaÑCv�_j�� pP��M]�1�e��q�k�Jld�oIZj ��(=FU�"PǢ�j��!� �\�k�p�\6�3>>U?��=.V4� /L�f��W�E�ts;����"��y����6^����x�#'OJWT��G�0����L��$����`�(њ�c��	��e�Y�m��^O�P�-�gX����ͧ<����8�^�DыR[�9�!S��-W�%�M���{����M���r��࢔�*�f��t%�|�.g|�'O�qz1���s9�mr&2��+��Kn 2���Obq�d8�L�3�������|l�'���lEs{�h�)_j��=0�l*/~�����o�N��@KQd��" u�$e0oFjZR�\p�r�OP�L���N=F�P�8f@����;�;