��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛����
�Fb�G�f��ۤ`U���oȚ�ufJ���g>U�;0�)�[��[\C٧��Wi���a͟��aoOL���D���Kj�h�4?��n%NE:Yi��b	 ���5��G��r>��T�CF�'�!�K�EƱ��!Pu���jϋ��*bئ�T��V"���￩���[�Kk��$�=篼{�^Wo"��V�L��b�V���.�Dŏ���.���2��n�����)�>i�,�	Y[��>a�׆��"�
�<7Ɉ���m��./���DSBT�pz�
�9����Ǌ���y�r�#�v���6�T�X��mB295ʥ����\|��ӻ>��һ��J�G��*�ie�*oP�;4_4v�j��/~_�lBI�3�uG�`wi�����^��kR��3�� ��$���)R[�ی%��H�Y����0��1����

�M���S�>��0 �2�m�qk����� �{�N��M�ђa
�Ǣ�|���j��v�uS�kp�;���]��=�J��Wo�	Jw� o�DP�������^2T�����zyއսwQ�9�{�IF� i[�^Ij���mNTFn]�!�߳�+�*R�:�x%J|�5RX�ch����q�m��W⏕�+�����]�r�w���fafM��%�J��� �wD3cn>�H�p�#��jv��\�>��o�5H�Cمx0�)��a�J�'���];"V�ؙ0#s�ϊ�1 �@�������~[^����f�����L�|��#[3`�t����H7��vںN}#�G-F�@�肤�晘����C��&B���؃|��	�v*8!LG���5��Ն�®Zjx��f��j`�U�FR30w�m�����ȣ;q��	O��n	��g�PaR���@����,Qi��(p�x�ߒ�g~���p-s�,B�������E�����`@Q�X�l;#/&��ğ�R��1����ۓDL��BW!���5����(E���3ۣ0g�P����@Z,��j�cU�B����`fʣ
#�N��-�\K�5���|~���!F[�r(�/�ߴ�&��LY��%E��������ִ��a���U�3�j�p�����p�c�c9���D��Ibu���P�c�V�G�m�^�أk�Z�@Ras7�T8�$<͌�ծ��	M����z�R����i���tM9Ux2�|Ǩ�������<�MxXz�Hh�v@�-���G���3���On��	�������3,P���t�~� iao�?�G'�]솠���>�H ���WJ�Ja�̸���H7s�^�v���m��*^q���Q��ف�^�I�e��4��ȣ�CEm��C�/;u��ug"[�|u�!\�x���VB���^�_/��h�`�IU�\��)3�I�&j�,�=�9Oj�Xi��Ɛ(�M�qA<�E�ic&/9*��Y���y;�������hVL��"�d�����Sm"�R��֥xijYE����ې{��/D�Ȼ|� ���s8R��i�/
��(��V�K�]�?���_[4��]�U�bh�jK]bȵ��<�^�X���`|���g��j��0l���_+n�/�x`��8��\u~\ս�ĸ��c(�cK�D�J�����C�쬲 e^�3~�ڪ��jM�,��H���C� �tX:j��$��`v�d�Z&���9�EV�}�s���\��u���i�jx<w;O?�� D�Zf�|z�T��e���������և{��X|{xVs��y`f��oWQ U�!��$�6I:b�:u�T6P7�I�[�����Y��b*AVr�,ߑ)Mk(��u/�P�3��bz	��b����
I� 4� vt4�z��D���$LA	\o�F�@��C9�?��&��^B��h05��R��҄�*/�5��x��2����;�YSԦy�5p5~�v���[�(x\��f ���Ua��^�{���JV�5�y���9�+�U�WiAL�w?=1:��u���R�,��F��#�_�m��V�Lb�L<�+��n+ҕw5p'=���N��aVq:���I�����5��`�ķ��3����~�4	�Xi�4~#�ýN����sE)� 2̗Wk��-�q�D���ݻM����!� _+���/�&�_�	�h��'��)��-������ڄe5����S B�����TIc޶��(}ؓ�Xtŧ�q�����J۹.\a��{��".��2g�������`r,�s2_�b��r�|le8�j��������2a������)׷��>���x��-bo�jL���!�? �f�f;'��5��cF�6 Q�T�kQ���x�l��T�aO�6K�Id6
��=����3��8������ ��;�E�n��Ί�݂��w|,�@�0{z���X��N)uvPb��;J_��Tv�\�%�]�4�1@���	_2�t�_-��@?d>T6��̒{��� �<���i$��h�ҷ�NN.�^�G�xI�z7��Q){u
�&#TZQ��1M0bη�E_r��w��]�^n��q�Y74Ls�n�� $0S�h|;�U��$y�������Ș��>%�7�������p����Z�� �،E��ʼg�ߜ�R�
 �42��5��S�τD��BN�'�O��l��d�;�j!�8V�SĠR+����)�����23�G�[������nF�3���1|���fg|�f$ϟ7���,�����,aЙL"��Q� ��H�쬴�Uꚷ��3�ȀӤ�[��نO�ù#?�(�#��������,;�7?�/�r�l�u����%�{�&-`��^��P�^�3���YY�&�r�N����j��+�p��B6&Fl\�>6 ��������D��%��c:+�W�v^E2����b�����cY��������~���,��~�B���]�d@8k���#��$�DhB'�/]΢�Q��rElpSb�:����Ͻ�ЧxK(S���@��|<��Eа$�V��2x1H,��=4~N]J^e�*n�ʁ��"�(.�!|n��Dؾz�m�`��h�O�#���w�G��Ҙ���7���hL�Y��Oa�" �{�PD{.?���m�?.�8�F�k�pѰ#�Cu��;$��*=rh��a�&��i�)��v�at��F�amʓv3���v{sШ�_�D!x�����ʀD�E�y��	|W� -K�����dk�4zU�^v:����ӿ���4�uW�n�t Z�jD�WN�w��9�Ү�u_/Z��L��3pn3<�YJ������z18�hH`��?<៍������`�/nU�����������Y$8��,,�Ӕ��q9P�2BE�B�������km�?cm��yP����%C�iUE������v�'.���uj��1׳~�(��_�����eS�j���|�8���C=��/���@�e�]hE6��h�7�t74�#]�j���o0����b�S��?���J��[��"����b��D?����v���l���>-�����IwP�^�-�U�OI���I�欱�v~ޜ۫����Xc<���z�	o>��c#�w1yW0r��P��y���&kH �����L��;m8��l捽$�R���,zT�z��	�#�SB�|I��I���3;E�{������_5��>���i$��k��/����xڊ�> :D�*)�IM���A�j������䅬��+�j6N$)>������>6Osa��R�Hd�y��~������5;^��VB`n���o0�o:4�#��ʕL$�bϨɢ�� �k.�
�P�p	Mq81u������ XiK/C�sXB�7�4���)T�*���mC�IY�Sby
L�LB�5V���<#,&�ii���?G��.<��gw��1�P+өc��;�_L�z �,�b��{�*���~Σ�[>����ܻ}|����t�᪙��ڊ٘`i�<��^��'0ӖiT&��Y>x/Z~�#SL����3Ħ�^�ϵ�RU0�	�99��_9� :�y���D?��˓���ܷ5z�����]Ϲۓ��~�ZH��A<�j�.Y��
�'��̂E�;5�dӠ"��W��4<Ln�y��1�!Z�$�S�H}�{��z_�z7-����F"ڥ5U�n�(���{�GD�yWY����F�?�W;[mx�3}� �:��;&.?����Zo�c	�SJ}qTR�o�p��GM0�x(�+���L�c�3�����z!b�AH��?��0��"�-q��0`�V�$ݷ/��Ʉ�r��lC��2ӲS
K�Y�o1���������^����A���.���/����x�+3L$�R����8��Iފd���Uc4_-�x���u��ym��}��j��#��'TUi,�f�ߢ%m��h�`,̕G��#I����$>��������8�c6\����A���:;�%� r�Hi^պT'��Rh`g����s���Ļ2�b�Esm�G5g�:E�y�_�cB��
�0Ԁ`�s�m7_Y4S���L�ujփ2�>��Jm�c-��Θ���u7�$�K�eK&'��3�`F`��G����FcT����Ô��k�A�$~���|�sE���*�v�45zqb�ڲ"�.o�H�%��:�պ&�P�FH�������8Wr�e�g*Й����o��,QA��97R�D�)<���y;�@SoR�1��R�B�ޅ�@�=��%��M�	7��ڡ���;ӱ<v[`��u���]��@�RʺQ��+�vyf�R���6�U�'%�����<#�l�,�q�L)�_�6�2f�M���Λ�Aҁx��]M�J/��q��� �����"=��|s�c=�_6t$ݫ�6؈��].���-{FȒQ�ș�ľ�����y��V-���[<Yy��2vX�?R��g?�3zߌ�������t��fx�"�ߐ#�b�!^������N�<�V���=ޒk�7�D�N�9m"�:�3G��˽�>�~G�.���J/����9 ����1���]�����(�jI-��W�VN߬��K:M�=�Q?����r�3�;��y_G�e��j`g�������"c:D��|
�e�Ab���d������5���$P�;;\N�D�}T���A��0�Y���U~���@o>�+�Gs���Y�%oS��UUyo�PWLK�doE��U!ڭ)AWL^�OAV�zX�^�l�vS�����y�`��57�6�12^���덈�R��;�'�� �¬���W��Z��Y�R���c���{É�q���QgI��,�X=���ƦsoU�}l�d?�*�XJŷ��/�0.װYM���0����O��c=�I�/z�!�}��r�?�_祋����/�v�OgU�<��LM�_p���d�v��_���̞�a,5|���*D�;`�9?7��D���XE��a���X�[���i��P�V̅�t�����{wՋ/�j�/��Y;�mg��ޅ�,��+��+M�\���p"�}6��%�voej�s{��yG=�ݰ<�N�X]�rk�T��,�Ϥ��N��[*��mfUlV=�F� �F1aއ�U�_��d��VuT:���O`��
y��N�ȩf:��?�;	Z�?X6����{��YS�y��4�%�2��!��R�����t�۬�=n�1p�E�w0��^'C�Y���}�P�\.a�����
y�Q�Qզ�먲@���������%k�hc�h�\�����ق���D��[�g�=�����s���\0]����1�p�Z+P��0���3�a���EM���rd�:�3��̷�k�),j�i��wA���+��שqե�����;����aa#��kRlY^���"�e�-6%����&�5�n��#�����̓Mv�nf� �3�'�\a��d^tP�҃�j��+h)�O����M���6�[?�.�f}����B��fj[:	��ϻ��y>�}@W���hϲ��΂2�8��#t=�?�1�S�셗���A���u�N�s!6X��*�-|�2sOAHik��0o��i.<�O�*ݑ;_	�sG�����#�h��M�9���XE၍�T���y����
��4��F�&��1˦ݸP�Ե��U[�2���^p{��gr,��۰�{�-V4���3d7o0�����Lm,�ÿ����*;��J�
c��������ZO�إn�e��$h2����F�1t�3�S��N	�B�EiwI��s�=&�;�����j��ҫT�:Ig���l�^����j'i�*
-��@{L��4�T0&��)Y��K�.rpE%����t�ݥ�z��f1D� �)Te
C��n��}�&X�S��¢V5 ��d����-ڍ�ŉs 	��"ɕ�8{-������}���~�?��O��ϼ���v��Ei�d]p�l��ny�u1�����9��Z��褌{W|�g[R�C���\��%�����")7y�sb�l笥��®.�������+�E�
�w,,kAⵞo�B�WV�lk��ѫ+������bBN:�L��n�YQ�yk<��xZX�_��H�$����rJ�_3�A����H�Z�4���S���0�&)}W�߿��Nw�y��6����5���g��m»����x�aUv=Ǧ����K���r�N�n�C>��/�%��C�i�ʷ��L����.�@��h+w��ƭ�jM6�=5t�N�i4��&	fy����@�N�0��H+��
\G>�_�mܪ�l���_�_H�k��}̎M�Uh-7��z�����C�jEL䢁��h�����C��>�CuZ)t��+��$�	���+,�%�-D��wz��s����YE�E�/�N\ɁH��9$���b��]�5�O��"9<�}������2�7�T�����Q�>��^N��M�` ��N������;&�!���&�9��7���a�\�s�8�d�n�߹�)��a����"�)[U����"�Ʊ\�a0'0��ߥt�� ��,J��В�-pT����^�=TKMp�[�1�:�'Պ� I+�r���^֠��E��N���˳���e6�*���#�Kp�}ݧh��v�,��+�0v�Y���i �p�h���R��b�F>�/o��&ss�y	n`�tx�oD%M�^,9��rjb�t���J-�=�lvZvDIwu`$�6+���t�\�Ͻ�A���Xڴ�c����r�����~*�Q�)
��E*?v���J�Ï�L�W'�N=MǤ��e��E�f/�:��ԅ8�Cb���ix��ֈ�訥w�@������bTO�)B;{��<f����/<�t�w�y�K�c�5���6���y
�7���� >���>�0h�~����^�`��2���-�V��[_ɐ�A�*=�y�T��׵��ˑ|:��_��+�
�Tx�Yq��0~�W����F��fC2G�u���Or�����N��)�넝8�����o��hQg�J�e0k�㵑�W��`���H�qh#�0��T*�
�Q����`J��?;�6��xe�v�;Ĩ�/�Z-�Wɾv9�0�[��qˢ:Zn%Z�(6p��t��nv,���&����}d7��CE�jI0:�\u@,mq��s4�$83�f4������Į1�:��#�/��GY����H8�_ٹmjÁw��$�A_��l��\e�����
��u��^f����f�I:~�cg-�N��q>��E�L�(1��uѓ�0�r���GnFK����STu�n�B��=	-C�(���R�1���{�}���sf�wWh��o�KR����˽ļG�%P�OSU}��7�{�8}�>��BN������h��)�_MJXb>�M���E]mb��?8��/���a�*�+G�|��@�?������t����4�(�;k,���VG�R��5R�0��>%��Ә�
����l���_$�y����f9B(K��������m^�e�Iql'���3�X�
d�O��K�KT�hm�jz�d	��
��$�j�1�G��nZ�CO_��I� �z\��UVb}pN����E���z�l�ڥ.�<���│ �¯���+.�r����C��v:Q�v����|�X�]�F	B=�@8{��x<�*<_x��q�Φw撒 �t;�����v���:�D*\:����|+^EΟ�Ubo�t�����t���ж�n	B�W���{mF9��|�Y<���ߞk�i�u��Px��8Q��)-;
����q��C�6�����Ȗ��Iè!��!����Mx���M"`�����x�o���O(w$��ԾQ���<ȟ��� -O��E6��˼�l�3�v����]�N�.��ێ�X�����j?ԋ�Q:j��M��T����%���V�FNg����pO5����O�04�/�9���M�.�}1S���m}��ٚ� !̰�nK�N���%Lp1*���L=���,6SS?&��3|M���e(b�)�3���~`~�1�
��_���Qc�G`oM+RK�{(��ιd�9����X���~�>-s���hoB�g]��KAhO���g��	��Dz؎��Z����� ��ۆ�RJ��e�wD��@�O�k/>ԙHq�5�|��'Rj�e��"�?�Ⱥ�`�IeITJ��C	c��4κ^�& �Q4[��
y�e��G��t<�3��
>�Aszп͞�!�������	�%z�q �	�i�w5"h���*�VZ�Mԛ��bVG���;��f#��Re��wX ;�WƐh�L�y��!�!�y
A��/Y�r���o����{�1$� ��^65��HR�}�~�F)��[�|�d�'�x<"2�)}�ۯ�XLL���	�D�� ����y�s$���'(�]L2X�-)�$�������j��r1N�g�D!&[0��w
�����Y�X�}i����]�}6N�4�,�@�H���m,����������Z�̶hCb�Vҹ���^Zwr%CjN7,�e��?%��BI+�V�]g�S�^a�'��5��^������"����)Y��?k�!m�� ٔ��4�"�
ͬ4�$�#pmI�rؖ0y�o[̖x��e�|��������E�S�Z=+	�Ԋ�2��2�ѡ����3�����;ٖ�yޚy3l���d	qY9���N�#1��m��y���H��C���Z�ur�/�BV���
W���cl�ȱ���4�j����#���?�,�߼�x,@��v�V{�2��Wd� ޥ���X�.R�{9zxk٥�E�	�R�
�����l�u�j9�`���p��u��v��F^���� a�t`��ak��<��p����YGy��{���,q弤5�zl�+mI ��O����]��l*���H�H�z��VXK�٣�&�H�̅�O�Cl�����<r_k����q�}���T���6�;t��+���;8o�z�|OW�ow<n����ҭO�ٚ&3��4ꐵ �&�bZ Թ�`dh�#ύ�y|��h��ܰ�j�[6`_6�RH�]�O��!z@������J4�̔�U�h�����r^1�(�Js0Ѭ@|��؊7�Vh���z��p����[5��4���L�"�ϫ|��˪	�e>�L�n�i�/;#�%䣑2ن4t Ro�d��H�'->i+J�j�dע�t�4)�@�����׮�n
�n��6F�f�!	���ӈa�j"�elk�)��Q����X�,0	��O'W�pR̛�,���֘`��1@�
�iFzn<S��7������ �#d�.A�g��h����ݰ�ܧ�h��گ�2���5�ÿݸ�JM���#W�#|�G�@���5����+�P���V����F6�$D��.z}��`D�f�����z�or{aE�T��o��
.�_��D�DVح�9,��Q\�@lѺ��>&zC��޶�"����6��T��8��������p>��"��9�Bt���%"d��H۰Z������z�_���C0f�����_��{3���/sЉ�6�?���
���*''�u6�u1�ď�� �L�
��u0�8�B��w��	H�*�яP����.��������سb �6�9�>)#ɀ.�>Ϛ.fI��R+��"A�Hܚ���quL�p*A�<eng�(�3��l�)RQ��Q�e66a힀B�X��T�A��J���H���xP"�V�౨f�Ak�qz�t�����R -V]�v��$���t�j�]-W�E��Ǉ�aӎ�/[�D��Ñɍě�Lݨ�X��S��A�)m�0�A��LT�Y�kzÈ�d��K�	�[��3Y&�k>�+�F���s�ED�&b��\��m�:7X;�<e�Jˎ�N�@��J��C`G�lcYH$�� y0��y�O9A���R�A��*>S_�gh�N��$�&S��%+_�)�:(���}5Pu�����6F�k�?*� ��NJ��>�~�?���1�ʵ#�V�W7���<-
��0"��x��4�׺Z��2!rx�A�K�i3�A�t��C]������e�0�=��8Cyh��"顸c��������t��%@jR��=��	�)�����8��=���kӁ�+s1_�_��t�d7�X'D�!�q�#}M
yG��OљgjX	�j�^��qoQO��w+��X�k��
SN�]��3rY������,MX�2����q+�L��qփJ5HR��Ы�*u?�4�	zy~d=ȅ�3;L�k��ȳ�3H.Ժ��9�G�zMP�ЊA�cJ���ԥ/��.�>�*�B�y2myV�3��N�%3�څ����ÖELʞB[���6Ŕ��9��3��&\W�t6�'�>�>��u.�#���R"��y@F�tq~dt�6�>�i�M���^��"3�V����N��Wc��-t��M:W/]�`��C�g���^�7�(y���pf��VB�憠���A�Cͪ�C���b*���,��vz�X�Y8�<�Y�àr�-lYK�.�sF>)�)�E�j���D48_.�z�� >�j ���s��o����qܯ�"q�<��Y�C���[�W̡垚���=��t�tJ�;�~�Rx9��$��m�h��wŇ�W�W��C���&^���
%O�z��f|_e;7|ThC>j�ɻ"�7���X�C�.�T�0����I4e��`��t��z���T⽊ؾ~+�ٜ�(���ń��άd�֭%���G0vJ���Z;�B �^'�EЊ���.�31cP���&o�rp���Ș���<��$�,�J�an��ɘHq�g۴?R`�p��\���$�Qm�o�w(#�^I"�� ����8�̴��a�sY�
�Sh࠵�[����e>�� @O)�	��$fݏ^Jro
�6t��o����*9��k���y�m+tN��T�I��� $��aM�=���U�(���Cy�.��Ufr|�{��x����Κ)N?�	c��E�\ڸ���0�uM�C��&���l��QMC|2M�ڂ��mQ��]$�F��%p�*�rV6�n<)�F�;)���VCG)_����G��4ډ`�����D{!�\��[Ѳ����#�9��\�z�`�1���_ܩ�o)xFE*d����M�EnG��	�[o� ��.X7��&�7��+6a�&$�`�����0?Z�A�#�)sRB+W�{�^^z	�l�r��t���3�ջC#�XU!�$J�/Az�M���V�P�� �\�:I;�W��QF��N+�ɞ���q���ux4�ύ��a��U�w�N�.Ƞ�7�1�&_��]m���Y~^8��k�$� !���6�n�95jdT,�b	����Ҋ@��jg�1���b[	[?%!b-|�2��s�g��RC�̜�*�4� �5�@�����'���AlU>��[({�ƪo?,�+[sϠ�hm!p��s��Îv���U�l��@�=���PR瘭q�J��+�:� �(Ϯ9��8���8��[-1���G�O�C�|Dh@�x|S���6��(J�+ �bkZ2��+hP�Y��:�=�*�сåQ��u|�P�$I���ɐ�J�sT-�)3,qk��#���H ��ѽ��͹�<�3�U���Q�}i�����j1�D	^lTw*?��-��$��0��`P
��*�X�4�C���I��_��N�j���
@v�xD8Xjfs�H�v�s��0����I�|���Bu����#�0Q�P;o-Rf�@q5q>L�b>���#P_Z��|	1m$ǵ�U�r6��gU�����Y -(����7JX���X��4o�㪟�Lǽ�r)�h��vudvD�����E��XZ/﷌�x�퍑�thCPA�El�5�y��w���B��fZ�"��[�D�}�7Ľ_�3��<���l]`�������Y�QӦ�F*9.;L�x��ڱif/�U���&�?��p����
�U�FM
�\:��* �yY�y�n{�gg*��aIw�i ֤���,�\"��_�K}��qQT~�P�%�s��F>��uV��*w��R��1�ق8PH;I7@u��m(6�1uhŧ�v��D����R��X��(�o��Ȋ*Z��V$���~a'���-hD��A^���p�	��&]�TJ�&���OT��u�-��U�P�A���SIm����FgF�s2�*7�Z�NN�Wq�����gW�F��.���ވv<m��c�,�R5�8�u�s�_�����ePꇩ$uc)�N�Id�
�Äe����hR�?��3����ω:�:�a�� �>�ڤ~�ʶ_5'�o���`�'���y
Q��a2F��[i|B{@��sa�c�m=j��W��
�ΘT~�d��\g1sU	��r���pF"�}Ŷ���57G�RCJ�5 �C��O!NB�W$h�����`�1h�ڸ���䤩�}Eek{%)΅-�0u�q.d��r��'�c��
�e��2�/�����?��&���W܌;�H�U�|��e-����}6���An5��z(\X�d=�`��É��i��zR�����u��7�R^�R+�����S��}X��h����z��^ɲ��Ś�	�A��a�2��Q�8e�3���v��0��� ��<X��0�K���݈��Gߦ�5o�}�s
BQ���o����c��
X�ߚ|�E7JB�
B�#y5!��y�iۗ P?㇐�.f�}ģ0��o
��g��-PQ�j�cl{��.Qtݽ].�^�F�L��>rL���l���[�,�p��+��$k�CsA�JG�I���bRd��is<�)�d�Z-�t�1֯'����gK�C4�F�96͎��m��q����O~e,5����Vp�1
r#5�����.&�{��H�vB�k��X2[���X��SPu#�����_�Pim8����^
69i!34�cP� ��l|�p-k�r�4�8��hӬ��Q7�Rٮ����+�H�����/����񖸍x9�n�����f8��:D��m�i��F�5[2>�i�	9�i7�ҿW��
W$�f@�3��X+�e�0�{��WK�M���Xa��`��Bu:�=���G��~��|�ϓ�nG`'�*/�Ċ�����U��"����� �б-�Bt1T�����U�!�N��=Ӷ'z.��C�����ިT�5�$�ږ�������ލ�ہ��nX�İWb�� uzť -��i�9?r
�VjD��э]���4w��B���P*��i';S��_]h���������Ň?�P_���_������s�D�|�,��ea�X����S_}g%l+���Lt��,��V��L��2PDc���	�9�*�b�U�J��T� �[�D_q/�ڨ;|dJ͝t�ګ�|����.��]6r�1%}�X���>;<ա�0�Q��t��{Z1�p����6'�r[,Y���4�o�ԡ�HC^+���ܥ9������܂�\�(��kY/���J�28��`[D�X\쿀��"��X6��^���:��4��v�Q�6��j\B^��o�"����N �)!��ܣ5IC�5p��3��]{Nm���S����\[Xo�2!��7�����ʱ4�R�f�q��;93�a�.*t2�S��%,�%��pB6�k�S\�b��X��[Ht�����.p�����}�xv���*����K�Ӧ'��F-4�S�T�\7@�ܧ��G-����3l��D���t�Y%�0g̹�2���
����� ䷻ �I���w|��ʇBdZ˃y^q�r� �����n�H�T
�$>R�:M��{Iz�˗����D��6M�<���j�k����]��2��I)?وu��ˁ�g��-��[�}��`(�{mA�ȅ���D���X�Ӕ���%<�_�]�4�l����{��d���ë�:�>ֿJ܏x{�V�.�Ui�f�R��Ҏ���?�S2=�$M7-���U����x���>Mf��P��{4�9=v�F�{���uXu+�蚷�����"�^�t	쭪��_\k��VMl -o�#�@Y�v�r�Rb��@���k�Vz!T�^Ԫ)�.�x�Ү�;q;�`��-�uC	��L���+�Qo2:Y%ư��^�.$g���g�G�Mj�`l��i�(��op�vD�HeK=�?ȴ�v���aa����9*�˯��F:
d����4a��B5�ņYv�S�y�����1O@yꧧD�L��H��V�2X��M���i��,?T͈�-�`s�� �3Y0aG�3�
>���n�:`�w��0���;�Qï���2c�ı?�����\�'�^L�	��3�X�f�lឮN�xwނ�*�_ÇP�޴�!�{8��k��}��Dw���Y��]vC��зN�򂙫��g��h���L4��k��0���7��*Q�����:��i�fْ�mgY�\]1��*��ө_���ol��KJ3G+֨˽2�^����m?�߉��gB5;�z���{���H�A�F��r�
�[��D����	6��4��wGwa����f�hJթd=�`$-�AE�Ur
�s�2�Ժ7	I�,�>A贆�N���"�$�I����v�9�WŌ�L�" �f3�6[���Z���=���b�LX8zi�ĳ8N�~Z��)�䫼yE�Q@'	�/I����5mM���N�2L`�˕ݚ�����<��G[/u����������5*�e-rg��|0��"�h=W�*Yl��3��M�kqP��!;�΅�?�&����Yᗽ��1g�0�w({��]��J!ߗy�'�-$�!�h�Nڻ{6�<�L�6g�e�'$ 5�U�q��X�dW=P�$;�'Uޕ\�u�U��Ʌ��I~9T��h��a��P�)P��4	
S���t:�r��|��.Ъ3���Fx��ۅ::!XY�]��\9�<��dX���E�!��٤���F�ؤ[�b���A�� `��sF��6�<�/_����{:�wq3�6{H�xId ������4G��\�d�(��]���w��s�.�H��
��I�ܽS(��?8h�	 � ��2$%TJ�:�7�i� �z��T_���Pz~��n��?��SY=���]��H�K�"�}p����M�v�U9�9�k�d��F�S
�	,-�Mk��u>x����0��D�	Λ�9���x�5����� ��K�?����%����٢�u�n�~>� е���{�f���-vvD�ȳ�b�O��du�Y�X�h�Gu���w�,���7vA.��^ܥ��[����
���Ч���G�&���T��M��&4^M�c͌�<���7��K,Á�V�X���e:�):�MR�.�mD����ˌÙ��v�J�W]nO�kO�P�Q� DM�H~`��rZU
P>����]���7e�TA�)��p��Bǋ?��s�Z��^C��S�u��)�Cե{��$@FtB������#�g}9,��K��+�#�ӳ l�P�,����K]}��s���5��'�#f��+���^A<m��vC< d<Uo��<S��.f'{����������)���Æ�ꢓ`5��r��%q���������*��-��.j��*%֙�~�cm?Y����O!�Ï��r-��́>oi�Q��\~;~mO	a�p���CΒ�:ɒM�G%=]��I�Yv��d�_ �q��ي���HWn=��@��¥D��=m�@Ħ��jQ�D�ST
��X,i����qk}�͔�2z[�F�s�!�0��z�\�'Z/���V�����V���Qa�������b-�����"�%�U�EQ��E+�1Z�=�����n�����2��&�)�^�>#��.N]*Q�4D���6�߮!���/��
~�*�t�@�`�ZPFu ty(F3GI��W��9�8�?�6u��Mۧ)Q�L���BX�g?q$�}��mg P`��#Hb���Ů�qiJ剭"§�@�Z㖰^��&��A���	��T�Z�N�k'U��z��O�@� �phbI	z��u�9��N�qr4K�u˴|��x�.�4i�Ā�<�����<�{�˒\��	Q� �Z�����N��Z6c�<�25��[�{�uv��q)�Kz���9� t\>��}w�<Yd�5��yfw6�Y&�Fj�s�B�IfkǠ��@�_��*��	߇3qx;���q瑨8p���z��p�'��A�J�2T��K��p�%�)K[�(X6�Jne��
n�S�9������<ᒑ h�_)�_z!��\�|�Q�s�b��h� ���ݓ�-dUȴ-7��Q����c(2��&�|õ�U�8�ް ��$��+Tb��u����)-�: ?�W����,�{�k�М*j��E�%�ѱw�=c0��NjŠ�  �F~�G��B5�cn�o��h�,���ʇ��hI�P�R�j�m��@E]�4��^ h��u�e��4��p5�ڊ�B�a��������;1>��*t�~)]���z	��+�R����^���:j1��?�v���F�C�qp�
�S{{j�|[���V�����"�Y�Hӈ��}�O�`�3��~LL��n�%i�$�`��2:ULD��~�9��/<R��׃�Vy3E������� ,��u�yϹP�zF��=:(���%�j��5���њ��4Ց5Bڬ����}|�������b��R�
	�=���3F�Mz�ɼSR�0��n�ٹɋ�ᾤL��K�bY�f�r���}b�Y�{��t����Ϟ�q_�zjo��n���䟧��!�e
j|�����m���z��ݪ�(��{Gv���I��H��!xxDpy'#�|\$G�':�����O�����|)9"ә�A�;<�pA�M�0�A r�l�������!���ʺAmI芸7\����3��c���RM�o�V���n'�Pg�aUEإ���l_��te�s���p�4�S�
 ��E�0��p�M�^k����A}�`U�Z`g�O��R�1z��C�y�����FʔZC�sVo�Y�������xtc���ZZ=�̊L�Ҝ�UEkľ��2s���#�,&҈�m
��F�~+EF���K&}(|j]��B8�ڂq����)XnP���H�FJ�S#PM���ǖ6[n>l��&@���Ŷ8%zi J��v&�f���i���L� ��z׺��$�g�������N�ѐ��l%��
y�ԁ^i�~>�>7ָ4m�)��#��xIYe���L�6�*���Y�H%��׉�M�9��ܩs[ I���涥r�D�#�X�k��v�g�&#���|�W������9z����ϼ: wGB�MW�����x�r��,C�Wa�҃`� �н6�⋯�"�!�Imw�~����u�F�a7�c���9�꫈4`�'���6 ��6ӂ�l�Q�A��	��a�_��b ���}��B6���@�V����(h	0�� }�^�� �Zt}d%��7�ػ�ܰ��a:�^��1.��+�|k|��R߃��,g���e�0)�<8K��T;w1WA�0��'��K&�}ơ��\c�A��#��퀻�|
)�3��T��Z�i��U�(��J��s`�j�z`�ک�E2�m%�t˷���aSV���I�/ˌ�v�]bnw*��B񽤞����uIϟݤ:YȜśoK���8VPd�$�t|y��t���頲$�]�UL#�Ȁݡ�u箟��C��4�QO��*{�G9��7m�h4�B#y���|1>�p�&8�-��@���@+A�|�To��� zA;�'^Gc�[��$��M��E$5��R���8��?����1T��1d[�p�-4�?';�
7��i5��G���DC�~�贛�6�'$in�ǂ�ń.x�O��z[���s@�s ���61˛��Z����&��Ǭ��F��"
<�ک��i��`�;�~�V�����[��{%� �	c���4 �k�Ek$�`��Cp��ZrPD(��8n�>�U��(�&6R��aT��,�M_�݄}6�@V0PB�ї��&�m�Лͥ���>]�E4S�H�~�P�6��������<�}H�js�@�\c\����r-�<ׅ\���S�C �Qu���> Zl�r׃���&}c�i�X��u)T*�b�1����ID0����Q�!�_�����]fda��D�.瞸��#�?$�c$��߭y7^�-��1]�3w���MWN�#�3��;g����ن
Rj��~�`h�N�v%v5|�������H!xS*���ٛը������^+�S.��^	KS���1��i�G�d��rP#�3F\����Nn�^��eK�a��0�_aP�����\�N)v�v�̄�5�#�H�w=gw@͇�]�}#��])m\*����
���#b�	�=�g �R���;�s���ߴ�m�sQ�R�"2�N.�3���,��<��
]��նRy�<�#D�g+�>��%3`�%������ ]2˾1sr�l�aj��f�w�PkQ��yo���F���T_He2��Tj����]L�ʷ�>֗n��9��5o����f2�&3t��
i�|a��M>�Dz���!{F����g�3���F�t@���oS�V�����^a"�[f�
��*0�է|��썏��J1W��Xm��'Y#r��=���MT��]4F�m��G?ߚ>��\���3�\���mr��m����X� gu�j�����[�N�88�W]y+��׶�c�D�+� �2�/�R��/���o�P�no�<|p!��.,�8��R��g]<���k�#�s�r�����U&j�Hh��V�[t����ç����S��8#���:��A���<C&﫮*T�Dt4L,��ӕ�n�s
�>�E��=��xۃ����Ң� o:�}4;c�6͋�v��1�u~���͂��M��,?�A$ �j�CD]�K|��9>.�X���+HS8Nlt.P�Iʏ v�y���6�7V:��fMI$����[X���p=��dD�#��Z�`<��XA��q��S;x%�U#�K��g���m��y�л��;��m�1c8�i=�!�`oB��{���PmN�}X�jV��$�J�k}� �X)�oH��¾9H�z�3D~ձ��tq
��<�����N2�T-�� ��0G@�@6��<5��S��W!�4�QQ+�@UIs�H�vCa��U?���l<S+�D�rG�2T���66�PC����	�(zC^�,�ȸ��P-<�ٷ���@���f����z&���x�T�!&vU���2����/��]չ^
Z���*iop������|!��_�m�j2���C���G^��/O1�9>֎�Zu��pf7A��O��*��,�nu�'�Ѓ`�
�l�G��D5=&��H?)����)rn}�~zB�
�F��fJ��(�L���ݰ[��%����Ĥ�-��@�~�~�tЖa�� �TVW5tu�ֽҿ�!�2��3E4����s�RuW/���T\&���G9 �_���;Ȓ'l���v�1��%�]i��NM��Z��b��I�*��Jox�O�ly��9�lLZ^�L3�h�	�r�wuR���J��!��X�8W\�3w���k8���[�}�L��H��C����9M|�p%�	m�Q�uA��͂������Q]�!�fxMzm�x��.S��3���(��i=��?I�h@�%Y��hO�nO�ō*s�V�*�\@6D���j0��.��p%���ۈO��B>T���t��Y�$�\;tuТ���4�A+���K#[Z�p��fd�����<f���F)�Rd�7�����#W��O�Nt��	���QP�Pt-�0"���[�,Y#<���n�1!��#�[�ʍ��1z4ߔ4w�n��x�f#�������¥`?P0R�u����c'�"m�K􄴐k	�~M���M>r�aBHV�D8&P.�@�/k|v&U_u�@���d���� ��f���(�j��?�����/� л�ɋ�N��$۰m@[c�$'d�sZO���^N��*Մ?�j�ХMV?o⊔�l��q�\�$<���11~�v���f���*��.��u�/fr����6���`�]N]���L�ND��bo4\�Co�WS���Zp�O)Qzާ㯹�VAK6�sb/��%`�P���vy��܃�s�6��g�����#���]+�?��VR��`��2}2k�3��q����:i�|�n)���Z�6�mןT^�3oޙ}}�F�Z>y�O��`O�|f�c�<p�C�_�.\�<U�ʊ7>��2a�40�tX�
�7�-��(�}j	�{"t�r�/gv���]v]l��������x��~���mĝʵ�'��,C8��:d���
r��ge�S�^��7{ՄV}sV��a>��J)4��&���k���z�߮%�l��e{�R��z�z�����#F��䲠;Ӡ{v4��Q�1H�Ũ����K�$vcq�T�Ć!^��=�X�=�&�2׏R
�;(���,�ı*���Z�z\������R���y�!�W���#���:]�,���5f��y��v��|'�-�5Wo�{���)%6p'ݨ���4��I�]�MQ ˝�E|�{�[���bC}�y���)x�|GB����!��MVf�E�夋��Oj<(j����8� ���ܶ��kCyVV\V� ����{�Lt�֌+�mQ)��\�p;�|G��,�t��)�,�)�����I�>�&�$-8�].�!;T����Vt웸dѩ�Y˚�+G)����_)�~|�}�![(�:�k�P�/�x Pĳ)U#�9�U����,!�Ķ��|�+�f|Tf|����^��o�/u��hO�$�x>���冞�]�Ŋk1�UU�3x����=�>�T��bz�ԳR&Ad����w�XQ�M�͌U�����Cء�*Wvtu�xU�h��fL�5�5]�Fݭ�=��h�.kQ0B��>7��9�,�6wn�����U
5XSȦ���0�����!��ctR�X��mX��{��]�-ot��YA�+M��ahv�k�%Iҋ����b�Q��7
~ ����H9�Ѿ�~��;nI`����qAIe%� �r�d�#@�0��f9\�<��%�7U�4��*��y�8MŁ�X�k�7�m�3���t�Oī!K��zq��W0�&���1�`0���	m��ۧ���j�ҋ`�0u	�S��M��P(6��)?m��������Fo��"y��5ox?&��m\�,��qM��7��m�+��M���"���0��o����
�S�Zp���Xqe��m�߼���"�%���h��?8���(���E+���=��F��~#!�����{���e�T�b�ۆU�?�5Wq%�6T
����͝�N���BK�Z���~<��c�O�X8�)۶��1~Ӵ��'��TX]\���e��i���<�&���: aN��[�xG.Kwn�"�b��
�����g��u�O*X*��|�3�~���C���D�Γ4�i���V��eu�B�t���P���U$ٯp���-wGb�<Qzh��=�3�r�F@�3D�+�"�b���[tx���IR~	��{Cj�5�NǦ���iP˱Z�w�^���($rӍ���p��zMّ�,x`���H�^N��+	��Rv67a����;���3F����e ei�aC�Q:T@��ՋiR���o��
W�7��C�J��P��� f՗�Nx-M�=VT+ӌIP��B*C�t��)�	�C`ZzԱ��������hqN^�9���¶����~}�2���C�kP<5y���)*�n�۹�_T�[E�l9�Pz�ԤS$�8�A��y�~�Hx�^���(���{��d1~J�������'����SD���� ��M����-�<�C~��)�bi#�w��v�8?���y���@b�.p��6h��o̥<�P��h��c"�x
�!ݿf�?���<un����[��A�n9�T5���b��u�X��	��L7��M,���?�u��_+OD�G�(�d�ܡ�,px��B5��=/���N�tXW#<��XVl밒K�OA;<-�*���w�>9C�p~�7�$�����f�«��2[�} �Ͱd��sd�ee@�r��'*9�{w��)=9^�F�����ɖ�{n�+�4D�<MQ;�t@��t��	�F��ԈT�|������R��&0�nsvK���3�~��z���zYYQxw.�Wer;"B���P�-0���&��.8/B��c�5�Y9]D���@ǭ���#�u�EO���B��
v�w�N�v�G�~�+l%v�N�RB���\���#�O���߾����#m+��
�tE��+��V��B��zjC3Wξ����a�*�\�J�I�[�W��i%�?'�~k�C��|C�Xt�S�I���(���Y�"�+�z�m��˩ygԛ���e�1u��c��D�vmB���l4=�τ��X���?�u>�X���F���-� U٣׍�`E��w����b�53a���9cb�����	)NnlH��:�ĿT��
���Rk
���$�� ٺC$L�������r�C��l@wY�U�+��?�BtS}[/T�w��U�<Z�"Ûs��Ā��$�����_�|�K���Hx@��옇ɍU����6a;�W�"گ�CjJ����۩1pè޹+�~g��Z.���yBr{��[�K�_���d��:�W�VA-�ݓB��-p3r�U2d�>�W�����R��'uF�oL�_ae�����f�V�RN
:Z� �9F���7q����u���A�� ������!�f�W E5g�-�b�&Wo���hu[Y�0
�f�P:ǉ���c�
V�%�U�Uh'@��Ңݕ�er�P�8��{�,+�ԏuh����2�-b��_�#��/:ē�.��c1XrtX�J�-��A���)ˍ�ݨ3)�[~5��J���>>C*ɴU�W#!n3���"^���.�������>+=:��O>�n{�i��G��4r���+5�I8ꔠ䜎AЏ�,�+HD?$�}Z�v�4��6��$)�q��+�]��g�o�Df�n�U'0oV�g9�f���yU��䔋�D}�͛�C���z�=�dT��rr`EIl�~/���&p�k��F�����Ϡ��%�z0������i�q�0R��2ؚ��M�6�a��[~�T4e�_l�P��=_7�ʴO0��s,O�S����^L��m���c/^8`�� V=��m��N|�A6�)���4=���p�i�i@���W졾~8^0�I
�۴� ����5ǿ�ł��e�@�Tk[�^3���,a&���w;(������Q�w)LaǞ�pI]�-�ۡ�riL�Y�2(��n�&]���}YPy�P�IϤ��g��9���V����x��&!/3����_<$���_H�ѩ�'�����-m���FE���������� h�|�Bk���-"t��ܴ��#��-�N�(jx�q 	��[?��>]j�����F�S�n��wBm�ID~���D���������<c��+�Я�J֋�*�e�!',�� 3D~h��@�0[j��K�zB5�Ӝ��U��s�\�g�;�QU��8J~m�q0F߿�	n���XEA����e-��fV����������6~(���Z��}��n�Q��gX�vXH9�kѬNͻ8\.VF���h��m-�l��`���+遯�4=�µF��~�2Ü���4H<vZZ�AK ��1�S4��� $�}�^%���f�I!�$29����ש�f�/�|�	�d�]�u�_P�׺瘬9����+�׉��`��M��vϢ��7�x)�٪�VHq�|38�*���L ��W��l�5�Or��K{�w�3N b��2�)r�ZX�{Km�S�z`�i��}��78b{j�H�)W��I�2 ��{  G���:�G((�2��-��a_ӆz�,�{�o�a��LF׉���x.ϳ�w{�w	��8գ�X�����D7��_QU�ߔ��Yg��1&v�YM��m����.�	P���е=�U�����3_�Y�%�'Ϟ�j�`-|�G:l��vE��,2��:h9����ǧ2Y�%�~
>�V�LI�;X�|����̜5��=W�z�1#��}ȸ/�$�40�*�
i'��/�e@�M���^2�{\�I��`����G2:BWɇŽL�6�7n��k������$i~Q�d��9	R�7  �׸�p�Op�l�����9:]~C�Q���������[�ϴU�C�Z�	g&��iL�TUA%���q�]�J�CT�;Ww�o{��%�����=�B�7
$��ӻ�7���ȴZ>Y���щ��%%q���y�e$�����+�w���f�X�����j�_��Z�y3H�e/}.��'
8��P"Q��@����K�F�
gp��x2�_��Ę�y*��)r�I^�H�n;E��SѿO�_Y�������X�`ƕ��?,�����G�Q���0 �-�~A!6�N3��E�xU�o��[�<j�9���*�zPl�/���������J��9�f�*1��	qJ2w�T�,�9G��t��cP�	A� }� 4�'"�@_�Ϯ��2u�A-�+��9GHq�,H�-��k5xs�4��%�p��?�K���thk���%�[D!�`��k��p�g���wW��u3�h5|3��4|Qu!ztf!�%!:�׵��P��~"l��;b�H?�	��U�4)���p�算wI2ś��Is�Xs4�䩢a#�h�J?��rK�  (*�z�_9_"����:�m��,�+�0,�������M�$�G{�8�N�&p������E�^�ls��(C
��q�%ϰ�h�;y�dݬ9�,�oU�4phgʓt�6�_]�Q��hҸ��B���R\CQ��Gظj�/����?���	-���A�,E�1,%�g:��,@G�D����O�b.,�M*�(  �^�M:��E#5�%��rF�(��������\�U���Վ�7N���b.�ԤU�S����X~ X����W�`۔�`5�S�������`5G��a��]a��z��2&�?9VZN徐�g��Y|�{��},�K��h�u�d-��a����I֔�K��]��	��R4���`h�D$/y�θ�dN�5��h1\�飂�Ր-�	�AP%-���3���i{j�Hu}m�iW�/NA���W�}�!�#U�7��T�C/^��o��O�n��A8c���!��K�^���<�c���t��J�x��^]�����@E�l���(ul1b8es�b`�CN7�y�j��� j���ϔ��w����72T��m�`�!�����p����́�,s��zNk@e&C�c7��j������&=�!������,�7xm-��
{ 7��_��[~�?hu�����^f�gk,�!��p� ��R����K�T�.�z�F�-��)�����vtqrp-M�`�/�5�3&С܀s$�;7et��&�zֹ�sz���Cl���i�}�b��a��ơ~��b�����ړ`_�M�4���.��)���#�9?�9o^=�3���l���,o��Y:�'�9ֆ.,�XYt�O7�N�¹��[�	ɴGKx�iN��z�1�
�W�� �g�!����Ḩ1��[8�СXz�h�_Y�=��^g���m�pʌ���B�hl^���a����F]<��k��Kr����a��Tp���͢]A���d�s���kAܧ��fp$r��7�t{�?O�m�X��Rc2IC�s�� ��v�kYh�재uř���ʻb����y1�n?{_E�կ{f4�&�F��O�3G�ʸ����f�^��V&�DJV�q~�W{��z�n�R⏮\�Yx,�e�
��U��[(�I����"-$��&�<Mië����h�^�(:�)�����F�*Qv��H3��Q��8��Юv��m�Y�'W(}��.X�Ѿ(J�Z������%z�Ѡ@=^�q;!nT^Ґ�����n������dA�߷��m���\��q�i�[S�v`a��a�TvK;F,�qJ�*�f!9M��5ܜ����oH�*Y��@O���xᎸ�"?0��`L�Zr��:_��g]>p�}�#��oX�6Y"V�������!��͸�� 3u��L�<Z�\���/�芴�>x8�+.^˺��ܳ��I�%���SBu�*���.�r�$��Ƀ8x]�L:J��)�ƽ�M�fJ��'{X�iS;�H!�����H�}B3��8�p�7
x�:�'���D��,�^����w�7&�EܽkF��I[�b �ܶ���!�q���S �kֵ���ڭ�YJ������䏥]��ws>���d7�H���>ʮ�eH���X��h!���������I�2Ώ���>��Wˎ*yhX�j*7�)��pe\���_F@ L�[�V~4R���u�w-[�O�yf6�'�u�ϓ�.�x�A(W�&��-N�7��q�MN
V�z�����^�>�3�ÈTp#��Um�z�+'�9$_-�9�:}�c~؄}�	�nC
�<�����?�ڥ,�k�!v�t<��?�>1�h��`>�Zț�"'�7r�o;4�x�V�9�rh�":�#� ݿҶ�bJ�&���ɜ�UQ�8 ��8�"�5f��! ��'�B�pC�?9qX�v�r\ߣ�8~�@�"�YQ�J�$�a{�\�ܬ���i���+���Ĳ��[X�/0�U�  cVQ@�[\z[��M���E5K@�5]�񸔴�r��X��L�cI�<�a��*�6re��?�ʝ��Y��s�K��] �l�&ϚX�`6>��N���iC���	��%n��3� b�^T�+��yz���B3\�	�H��^Õh��Z�P�J	��GU�j��W�d�^��N�Z�c��X�� �8�rm��vp�I�D��4L�@�$gp�����t�`�&�^��7���Vފ��E�1�i0\X�R)��^�������x�=�_�Ђ;
�ǰE(&�K�X��� 2���e�Q�B4���]j`�jzHG�� ���UI�n
،���/�G7�0�����q5�5�Т�'M�(�\�O���⣗��닲����޺8�D�����7W�Et�	��t͈p�����E��>^���ҚG;f��Wu�8�W�ͬ�e�+��W{A��LPI�=0`�5ju$��}�[��/S�%�T�T����ԯH��9= ��/����:2������%m��_�$�� �I7�������� T��x�\>��/,�H�1<�8��S�i!����,y�lJz��g2(i9��Y2��0��L��n��V_�c�O+'���ϵp��~�����Eq{�h�s��S�ձ�Q'���.'`i�ϯnD�RJ?��SԺ�����~$G���d�~mf��}B��È�*��n�>g�q8�:=�/˝����V�����w�	�([~��1�	�k���@�bYnA`��e�Z֋8��ԇS���;Ȳ#�Ҵ؎�]6��ʍ��%ʉ�tV���TY��mCLvH���Hv�.���PՓ�"��`'�����$��F�G~m���*����Mi*�FY&�`����#a�Oy�r�t�o �Oo��z&�|ۡ/�9�<v��?���e�tr�.i(���v�a3QTR�h˺'k�^�� [����W`�ׄ &�jJ���1�ޠ^�;�u#����N���?�ꇙ,�Jp|@�WC�M�4*!5�(o�s�q^c�:ظ$�� q�� L<��q�Z²�F>�DA�d��|QBz}��x�;�)hBe�����?�NW�����0��Aa 7g�śVj��&��/��f�-�;v����5-0�����A �S.��Œd#�6j����d*���\�d�	)\��=!�5�1��3�t2ݍ?k�M@��I��#�AL+6��
Q�$^�(�0�z?�=��:�� �~��M����5Q\��y�:+Tɀ��4[d���ğ�hX���2���}����f��Zz���EX�V��|ԉ�4R��L��?���1[�W�����Y�Л���εZ��RȤȩ�0�Ā�A*g'3e��l<{�$rB����T�%� 3��躢1�ۛ���"����L.svο��a3�Kb���Ґ�����Z��a� )���#��ơ�4���^��X�dw�H��Ds�ۡ�.�X,#j������	۝ؠ���@W���0Y�(i C�/s�R�����d�#��@R8P�;Ty&�������@�'v�"5�����l|�ǀrB�)@��6�?k�K���Z��I�e�{�2!��Df��߁�oi�^����p����4�J�2p�xu��Y�ǧ�㺓�ץ��H*CN�Q<]iE|���N�{�4�4��h-D�߭Ǒ*ߵ�e���TPݻ���F�k��m�XU��V�l�p�P6�c"i�Q��iE�ӱZm��zH,�����B�9$Ŋ���C��۔D�l�2�sN1u�&7 EUNn�;E`�sp^ˣ�R��Nf�(�p����h� #���x?�؞��F�~����Q��k0w8l�}�� 41F��b���_�?+%����B�Ibb��Q�8۸/�ʣ!^ ��hE�Mz9:�(|�g�۴���&��]&����o�6d���vv%_���M96���~��;Y�:��}E,���,��k���&��fE���N��S:�D�X>�e�������:�x9���t����~͛$�r�n��o��7/���II�� �gA�<���s �����8?X�+���[q�AhI��j��$��(`!��vw"�� �W��P!)��t�=�vOԃ)J��y�_�/���q��X���U�m�?��m\tT�A��>V.�>�ƍ��&1�RFz���������i�#��g\�)���pb�vH�F6�5�=��v��#u�н��ٰ�5��N�u��Wc<�;���/q�6�������ӑM�Қ/�A�#,�-��u!\f�!�^�osPg�צhn�u�������P3��oO�z	ˑ>ƪW��^�i��t����y7g��P]#�]F-;�	հت#u(W�wJ���j���j�fO�"�1��� +��� ����5~�+�5䖸E�m���\���t�-��`�b"�(�J�<z~�����:��g����3o(���Z`!�n�N6b�Vx�"�<SZp�g*����n���6�V�窢�2��],L��΋-	%�6��0��p��ԧ����x%��5�K6�D����\?U�	P!R�M:��j�5B��k�l` I��s�`���z��0!|���mwغ�ea�fj���o�V���BՈ�0S ��dm�Ƹ�"�I}�˄(򇚬=�����F��wJ��l'��Ň�c��m+�j디��/�pd�d�1,��D�l	哊���^r���(��J�~g�,�h�`�K��S��7�[R?���!訙�N�%��o �y��Hk{RJ[b�����t1k���7 sr/l�Э<�+���3f�{Q���ɼW�6�>��K��Vh��da;�֞� R+b�tx�_��R}m����1����5;4[���1n ��v�-���iˇ$Q��:,婢>�!��vs79�ʂ�6r�&H�1�z�̱�ra���o֪�{|�쁚�k�����we��`ٕs/J\���\�x¾C�#}��-�I�X�d�������)��虑A?9�`	�^{.t͵a�
�:���c�J�1'�_��=�_ƙ��VkJ}d�������Y"r��c��&�C��(�"�?���-�l��+��&�3� �].�C��	�-bu~G��P�˛���;!�N�}���ǳlu�FN��}�Ħ���H��1�,��q5�YQ�k���:L�vN�0P��%��Rέ�t�u�T�ddJz����d���64��q�<�y�����24�g$'�?��Vk2��¸�g��*�kiNƾ��S<�yv	�����4,vk�3,�y�H37�Ns	
�7( <�O�@A�ea[A���j1){��� ��y;ݍ%%u�8�Xp��a��V�6_x������K�r΂P�u�Y?;�
%HNψ8ƨ8%���$�����s"��:��d�$r!L�>ݩ3 �4�����m�� ���Uou�:mB�̓����܌˽A����fX�;�L.寕��"�0tz�i1G��~�o$&6�|����C�}lol�G�`�a��g�u�j����8�*ƣ�y|O��'���;��G����Ϲ���>�Gk�W,u�B�}�	X�ZS�����`��ƕ��ϙk���kw���{���\"��؍��K�6�������:Y���4��ɛZ�	*}�#�07�w�syE���]$Jj5�bê�jn�b����b��ܓB`���t���P�ߎ����S!��͋ߛ�6�~�u���4�H���D�{y�b!���wj��Զ�_�xĭ����}��uV+n��rq�aUO{���*��RL�z4�Cx�ID�ro���O�Z|��{ۤ�F�0�*+ۻ��vD_� ȟL� �jN?�qK`����^@<I�?$c�L�dG�J]&jM~�����9�C���1�`�N���ƦQ�FH_�U%,U|�T!y���7�od��>Z8x��<����ˡ�����2q�}ݒ]�Cգq#����zLΫ�zR�7��f�r�(t*�򏊑���
s����a��|��a�@J$e¢�\Dۀ�|Fd�+��6����2�N	�?��#����ͪ���sҁ�@xO��Ϫ�<��	������1�{�����e�&����|_��?���$��3T*\��տ��i�t�YQ��׭Å�;)��j�Q���X��\s*���[��yx�� �h����mBd��%&)v�q�+'{��O�Fg�f�>�!�7L�o��.?V"~��`%�m[����l�,��*��3��b1a��ra�=j[E2����`6�'R�MoH�a��>4V���v��'~���b�p����!5�׈?��8����.��u�\R���]nwO����Ņ/�iXJD�>D~�����6�;������wӵ�xT��K ������a��U��j���O����E<�p�Hxjީ�c"�UfԤ�xp��p*�[���[4�9��ȴ�������i�ЅE dT������,�+��3��N�v�P��oZ��h�0*~ [��o��n�g���0N�� �9�y%���1�p���O�@�����A�螾Ude���?8����Q�),c��A�ST��?�X/�h��<�v�#��R_D�I{��'  ]k����2����T=�'#���@�і��;�#�H����Ǽ��� ��Z��U�����\��Iރ�/\S�8���D�U�����tՊL%���6�{�x����㩲�-d2(�(Ϣ���"����a.��Q�l(9TG��'Ǵ�@bOu�R�|��9ݲ�U�,�R�{��T܍�NT1�Q6��(x��͆O��3v�3�UТ��+����Cq�=�9���g~}�j\ε�ٮ��Da-�9U�Qӱe<~�=�<�S?S2G������z���:1�)�g*�w?�t\���Tu]����YNwN�����7M�|��ƙ5x�,�=z�����3 �&��j��+=X2�T!�V(ϗq�&�W�L�_�[��t��\nH�h��U��~��f�CHV�$M�dl�J�~9R��#�T��)�%�J��������pm�[vF)� W�$�����vF��������
�˨ޅ5HVHZ����l9�N}���T���ͽ���a��^�e6�Ѵ�?`R@�o.��&�W����	�,6i�T�t��W�]��3�v!�^|�M�?&��o5�x5�O8_���3ń_�.��l��or*ԦG�1
�W�eCk��Ѭ\�O�E������cϛ�B:mj�@SM��7�P���TgL��m�>Se�L��������1���-��tr+ˢ(�� S %gJ�K �rE
?_�Am	K��6N� ��'F����9J�xTD����=S":6!��n��%!D�H9��a��Lހh'���:onЦEXQ|@��P(K����&�d9�E����-Y%+4�}
�z�D/Kw�)�C!w��؀�\@�S&�ݠ��~IcR�C� ��(o,H��Ic�Ȯ4�S�����~�s�h�^2\a�
�7�
1�a�R}����x�Au}�0s�<���� ?�ǥI��ϮP."����Ͱ��~;���3���cL���T�K�?�m����H���d ��B�/#őƵ�)`�wƾ��-��4rv͜��|s�V�z������T�G�K�w ��P����`<��Jn"��?�z�Gbh!�|��O_@n�hV$��Ѫ��)�?�#��c���ө�?��^b�g�:`������N����(�y�~\@FF>A�X�(��M�_n����Y��{��Y�yo����V�AQc���;	���͈�Kcp�~�CPق㥭�F�0Zvs-[d��f�p�jv1l��QLK ��C/�~G����u.¶u�^Hi�W��O]M�H�� .{)�$6g/�AC����\��(��Ո����VO����cR�8J�ib��U� 
TY1�""�G�h�KZ�@?��jʐH��J������*���&=g�Q֜��Kj�礊�U����m����zL<D�G�*�E+/%�����%��Nl��M y�ȅD���C�dy{"��H��H�̡	m-�#�%�L��\GK0���ܡW�G�� ��u��L��C�!�1�[�����7|~�yd�"������������ײ�4#�:b_0�#�Bcd�qG���V�V���4�Z�G'��3�Ϻ53������Z��+#���1��a���i�X�
S�8}���|[%�䱳�F�+f=��'�{����2Go���w`��kl��>B+�N�u�l�~�3B���gTs,��J���k��_�M�ޞS7�eN���E4����ֶ���Ш��1�z�:4�A�rY��l&��b@�W՜�����+g�ǴLE����S��(���Lc��GӶ[^
b��q��R�����#�!�hk�8'4lT��ѰVim:�.�?pO&ѷ�p4. (��6܍�w������k< Hg�}z~��RK��c\���g9�	g�Fш|J�֦���& w�oA�\@�G=��	�Gfy���A `��5�E�1;��Xl㉐3�[��P����H�𷭟N��ޅ����p�8��B6y����s#�A�x����^�Zv2N0'T���ͫj'���<2=b��l�?��4]l�˄��(�`�0 E�*�]�Ѐ��ka�+!o�I"Ԍ�����+$����kK ƍX����ٗ*q��(�ﱵ��6���J�
�40�@$���I1���V�7�Ym��v��8m�4�[mt	�vy-��˭�2��4h7�e`,�7w&W\���ba����H��w�q�L�ե��U��`�]�@���~����5/�G��)�HeU���@��خ]�W�&�0���!$*���v��p`�K����,C�������ʜD@oE*�^��r���w|���N��>.��M��Є�������iz ������f�{�pv�Q�J_uI�j
߆"��2Ku�����f@B)��*��_\��w���S��B�{�[�������0�X�⋋�>�OtP=eP��ɚ�:7`�(�}(A�&�-��9�/=($D��P(&�����:&��c�<i%�F��g�Zr��ޅ�������i+�S�7��ե�4*ax:Ĥ�Yͭ�^k����v[v��b��`��Y��~��}�<N���?&��q��kp�⽃�6xG\6�T�d��M�Y�v�1){�.׽?�3B�Q�� �&<�������h�s3Z�խ�D��l��"��|Dڌ��q~�U�1��9$Y�&J��ʮ:E�,$0������*�墳���x�� �x��`�a�/�F�߃�[�7����m�^�⬉����W->-ϣ��ݼ}ra�5��7v��}@��Os��I��t�5�Ԍ�@H�	�G����_]���CU0"}x�(Q��(>�� �0`�$4�!YF�r���v�&�R����B���}N]�ZY�-��N��廠[9�T��Vɀ���\\�٩�n=e�KA���\�P�_�筡+J���M5���ƍG��y�IZ���!�Z�Tl㞶�/O�b|��"n�z��j�Y�倽��Ȇ^��_&����`.�+%��/��ݑ�d
�-�e�	)��QO)�Ne����x�NQ�,�ΫF���c�0�J]y��<<Q����n@ N������N|�rL%�i����-�v�!(ۍATv"\qBE� �f6��6-���� ��d�A1|���o��ȡ���Y�Q�V���a|�!j�M����.��y2R^��H�a���m���(/�?���8ˍ��Q��}�O��cr'�C��,zB��7L��D��{,�⬱j$B�����"H�:׶\gc��cmM� ��d�O���<�d�;�P�b�g?�����%�F��ub�y�wT'%�~���I�B6����䁇=sP�J�.U4[@+�𷎟�}a"^�}�W�����;�EIB���:�w����hO�4Ut��'1y|k��`�Zi�u�����H�Q�A��x�E�K�!�b���YX?>�S��z���Y��`��)_;3�E����IC�7-��c�i7��7R�'8�X�9D�M�`�2.W���f�2����k��qӖ���i�E]��2�C9Ag�`Ps�*߽�=�&8�o6��s�[NU!C6��9ci�qfmK%幜�wY,�x���%6T=ׄ����G�H�������Ln�[ɴ��*@�Fz:0_�[z�膅�H���s��B2_u��D��S�.�՘}�i��l��V�����2|M���#��A�Z�������O�w	) #��O��mJ�<^u��1��<b��0��M`Vx>l�B�7�&�m���C��QMT��l��+����&��L]�t�����!�������uy�����$Ȕ�<�-�L�Jm�W61-�xN�Z��hzy;���e��ē����<;n:5��n >�'��(C'���K4��(BІ�3�� ��p��S�ov����$�X_Jx� ���mշ�:@0��(j� 1Y�����NL�\g	)����B�@G�m�yTՑ�}:qvl��G��7��Å�+�=#������-�^\�jٙ�J%	j�p��'�q�m> 7Љ��qz�3iL���;�jkP��<�/f�JK���
�ly1��H��ŋ:�[;�j&�c"�ǡ�<^�ȕ��S	? �&2�A�Tκ�/����M;������O׬ŝs�
�����d�[�m�	�����)��԰���aؑ��*��\*/���+E �c�Ձ��ϥγqK�5�y��A�N����߀m��o2Vk��1��]ů���3�ye�+ŀ6=}�aېp]��č�Ϲ�&�*4�����چͿ�F�鉉n�G2���i��؉6���Gh8�c��\h���Us��
#�	��QjQ�%�+
��d�E�,x��}W� ��v$�Z�Y�0��(�HhI��Wi��9T�,�Z�[������*���p`sD!4����1��#~��^L�1IWԠh
mT�/��獼E^�A��-�ށ:J�����[#�9᠐32�
wق���H�K6�	�pj�d	r/w��|� #aˤ�	H��-2���eC��q���V:�Qgǡ�7��I��U�I.�㱖���Bқ��)Mv���v�HR��Zy�u@l�k�r!��;J� u��ן�b}���N>�� k�>h�"oo '�@��m-����?���ڰ^c�`NS�+��q��y�7O��Ԅq��z�lX~x��(�*k�4���愰f�������j��fFkod� ������b�ڑ�s�T��XM���+�ءᎿG�^
�_�]���Sư:�N����hJ�N
��O�?TƋ�6�+�/����fr��0: S� �8Z� ��5� �hF]`�fzV�w�� z���z{;rY��H}�g���:�n��ut#a��ϒA"��Z؆]�7'LwȸEb��k
��E���d.�=G����I�h��;�L	�J\�Ɔ4j+-� ���e�d��aXQI��#���V��eš��f��0��|�&Y��'���8�+�	�63�!�ww��:Q�%�)\��-��R�h��H⻨Cy .��(�����F�o?�~,��?��V�Gf�v��^���9�PX��S��5��x����7�#�w�� �~��F������`�\`��l�+�:�%�ݚݲ��|���� pw�k"���߫<�aZ�<��y�_���0�����7���iU/!Mln���`i��`��y?����	�շ�Ҙ_+�0Z��t=��ra��!̫Gb��h�rİ"�&r%A�3�{�$�ef�0����i��B��x`�:��q�&Nd[�D�tc)⻱-`d?�>1r���V��<�È��֯Kvڎ-�9��[��j�:>��k���-�l^�7�I�b�~������26S#���Brq0 h;BU�{�ܮ�4ď�����;P�/�(�����",��v�&[�_��d�&��ױ8Ͳ�Q~,'�C��E��ɡ��I���W�m��8.��d|D`{c��x�o�,��
�����>pW6UX0g����$x4�( �����Ż��!|1�ʐ��E�zc��� \�*�hG�j�uμ�m}���{<�	�_�ϸ�r� �5N��Z��u~���jŐA�#�����O7ؚ��n�����m�����O: ��L�-_�yIȳY�3�sf[M���hx`���i\H9��Eu��zB�
!�J��H�5�d)�g��>%�Ѧ���%��S��[)�;���XS������FOu�m�\��������;�|�ن�����&��B�|X@d1�cظ}j�޽.�k��x�qRI ��}�_���#g�Ֆ�=���k���A�����纐u�a�i�����%�ACB�.S��$[)��b��ާ≍�Yd�|k 5�Ps�����"���v�S &{8��*�� $�`4E�%�`��h@^��8�q� ���$(Bt�-�}�1%����Kxh�|�>0\G������J
M�QX.��>��\"t�����?i͍�b�A�k���C�b��v�J�s�h%V1_j�ow�e(K�-?�����C�ދf��X��^�1���c���q�5�mX��?���}�VgͿ����n��Ϲ�(\��&�'�x�KV�9&�/�q�A^��Z3���26"���N�V��P*��^�����BU�wϓ|9�����J�PVL�O,'>[t\
�1o
h!�r��p#�'c&6�Ź�cfJ�o�;�6G�1�fꮇ������?����1�jAꀽ�m#|}��� ^�����S��P#�?����0�Bjl����u�����<�f:����?Ͼ_����mP�G,��G#� �^��i`c�o#��c��M��i<��⃣�9;��lo�"8�	T��Xv����*>5�܏5y�����$���@$%t�D�5g*�^X�omܪ�����}m@��}����ެ�KO�iɇ�v	u��|:7]�$��yk���O����젪�}����?s�
��W4z��޺�רy<Ca��uN $]��r�p2Z��X�n��갘�i���LtخAԵˠ�G�`0p�Ϟ���m�6*�<��D��uE���aG�MVR�d�[�3�����y�Ɓnh�ۊ�~Oy�Ƿ�J�+�_y1K�ƿ^�R@=�Og���F�o�0�e��A4����R��W5�Mw�K�ī���u4z�N�ɫ=0b�W���3��ɾs[�B��69?�����M�n�'Z�:*=A�;�yYU'�=8�hh@��n����l��`H�z�@�T6r��u����B�4a|=�Hq���<����H���"S�o����I�Jvu��o�Hb����^�>�V�s:sf��� �(�t�b���@aj�ֲL;�ɞ�fb%B)��^cB��y��*�cR�/x<��|L�z���N^�ƺ��5��Ǒ�gX��"�^��8��{#n�Ez޹��"'�dg��,y-ڑQ��&��Y6(�\@�ʌ|ZQt�41ۊ�3L�k�G����h��*na�B��2xt|���vV�s�'�$�G�H�u��K#�TX�L�DcCSFϡ�؊6ׂ�d074i����|�'M��3_}b��D��Fϱ�F�KǱ�5/*���)%Bҫ�bU܏ڃ��Y<5}X��,��>��̜A""�D8�/#}IqQ7ub����O�y����o�t�Q�y1i�6��Y$���<sg9�{�ֹ�F=b�Z(�]����1f�����EI�$�{�A�g�萐�cŀ���K�$|��ړ<�UEo�00g�O�5)�Qª#P��	��9sq_ۇɈ
�����]&h���`�g��*�Z����頍�za�
4�s����g`y���^�F��9�@�A��HBj��y�L_簸"(��p)F�Y8�Yc.�3�����Z�Mm� ��BH��Yp#4wT-�x3�*P� �5��U��t����a��J�1b�b�D���NEŌ�gcq<'*�h	�r�o�֋�MW�g������D�e�>&�}��rMA;��9�*bFܪ�������F[Y�<cF ��1^�:)��B�"�(�B�����tM��$▾TJ��"Eͣ�ȭ*��� �������St�a�rXY�};w��>�������H7 �[@�K��Ψ���~�����6��C28���>�cS/��0Q�P��s�J���t�__A��L1��0Ps���$0�nFDD�6Z�qV:�2f��^L�K�5�����s}醙��@�3��hЯ"b��4�M3����m��3�{�<�p�IX)% V�2������^E��*�:��g0�͍�-]���6�@�ّ#O���{�y���X��g=sI���<��KWZ��
hY����xe�EIt2q�0}�nQ�?H^W���#�N�ޞ�<�DЄ����#�~?D�pę�2�Q�<A�?m[�S����k�3��Y�h�O�$C��W=��?�+�K����ذ�/���>~�Sh,g��	\|����S��|b�܃���ّ�Y�.5���n3�(�̪���lضb����K�۵$5��q�jұ�]�ԑr����=��sQ�Zh8�_@R���#������1�/���Fx�~�[ȃz1�m*��V]N"������lM#>���&O1~�I �ՄHʖ�2�~�%����$A:9����=ع��ή�{��=��Q�A��C圭{���Is$�^C#�G[FSVb1 L%\y��B�^vx�,�!a�cG()��8�u޸<��Դa � -\և��_+l܉߭�>��H~��ۣ��H�$�ՒsҵѰ�3� �02��k{����|�����0�
ϻ�{U
��n,�B%����mS�j��	;(�4�-~o$��GՎ��DC�"�b�pUu6�N��DK���Aݻ	��Н W���2l����w����l��^���6 m4_��4iK��+�>�`��6b����bDj	JCN�K������nPy	�w���:	��Н]�	����muȾլ�Gm�닎gJHh\,'���T���d�֖���S��[p�f�`ׁ�n��Mtr�}S6sdp"���蒤&]���.����G������] ��s8k�aYc0k6�.�x��w��Lf*c=%e�@椶���'�'Q�D�aR.��4����l�#Z�G�-r���|����!֒����3
\]lV��L�<Wo v�Y��N��}Jl�Ə��)���X��{�(�h'2aW�=ī<c�0r����=��̑g�%��l�b�-��D�<�<s��8�)<�K���m�Čw�2�f#�<����?bU8�Hv�� �{q���xO2<H�����a��:-��f���(��!-e�ḢSU�hU��5t?Y� ��!R.��Em��� ���&�ֈؼ,�����M����I��t��t�%��G��� �y�"�qQ�cjH��<{�>� ��x��s��-��.e~%/��f���޼"�c8-IK��5!=˖@��{1{�a�*�爵lB��wt�
2�&�Wˍ��I���B .P�&S�'�7����z��Y��sV1k�P��ۉ!e�6�����'��� ���n�O���yC�r�o���V���. 
�7��H�坑ȄK�^Z�����l
*��b��P��'W:�.1��=�*)����UbF6�kJg4�)Hk�ȥ�^���m�kHyF*頉Yϸk�$D��h�ۈ(�K�����T�-'�&B�-=�����|5o� �b��o�u�.��Ue��orَ%^�yLt$��X#���է�i�?L�dXhn�YaW����Qg��'L�<��T*%�$ت<o-T����w�Tu����M�G�������Y*]_u�^M74�����(E^i���~�m��[$S�x��_�p��"Z�P���YD��tժ �\�xJ��b����/���sw��iί��@#�}K�������<F�ܫ�)�L��ֵ�#�%�RjP@qY6����`#ñ���C7�H��=�����4�'β��������T9��T�΋^�N��Q�8 �3-��?]r�[Y�ps����b��v@� -��4@�ł�
��m���cQV&:�blQ�� ��6_k�w/x���Z	>���l�k�rͮk�jz�`�:�CF�R��mKMlr|(8�7OA���v
��P2yw�Q�4�%�$�Z�+23-����Ѐs�6Y(����m�ط.q3�|�Ķe�]*��5}͋q����Bqz��N����ݵ��n[�p��"�	I��na�ť�ט��gX�����9����@�B����b�f� 
{��⟻�!�`�� Y:xy/ϥ�����}��4.�-)n/~�-�a\�{�-e���q;C�ӹə�l{�PNdjDlpBC�D�r���[�[�Ǳש�@���$�;�8G��=���2
�v�@��	4���(o��,M��NM�I�a�ο���nq*�ǟ�P���G��7�0����{��ș�0bP�X�뗓���Y8��s��D���)皈,ZS)�:Yk�&o�;��1J~�e��n����@y�z16���00�+��<��%6���!#� ����A���;�F`�:�[V���!�g\�:����j���F�.���B1|��+��׹Uv�R���{��lC��������߉�'���W����́:ؒ{�Q�љx��G�{�Z�K��V4��li��Q)_57a9xspC����)w��!8(O�k�HZ�/H�檤����.wo8��o�|�i�#R���hH�;���Y�ꂖ���`M��D��ÐN�(.�Uɡ��ۣ>�+�Z�����{�����i�~�h�d˿6^���mj�,vť���ݐIi�t�	�M�E�4���,��{�ĭ�����_-�ApveB/��(�?�G�� �Q/�s�_�<p/y}���cWo� ��B{}����sͻ'څ�����;ybH3+����v4��MԘ⧞��6�S(E �fb`{�S��S^u	��Z8��3:����q{��3�[�W�+��2�s����o�����D��w��߉�{A	pc�p��tM�<V:q@	��)��⍘�O���d��vD�ϯ	��u�GA�%�ݬ�8��T�ߝ��m�Φ�`�q�8RY�+���0[7��y��o� ��)w����Ą�ڍ#N�4���ŠxwTTщ���3��k�����[���
�D`�I�G��Qḏ|	��� ����s=!d��Aszm����J�Ήv���^�Y��.�Ӑ���l8b�ե�n�1�=Ǘ�5f�Wg+��o&��lo�H�p���A]oൖ$[�e#��?��֓gƂ�zTvv�g
�y����R�"�~p���\��/�SH�C@?E/B���$nt��j���w��:v\������pY����,��P!��L�n1��P�sOg����=G>�uY5Q�m�!P�� �9�a]����
a��1˸~+�������@}�0��lk�j���i��r�o�W�4_���M���k3��/%�Z�>�4��p�X;�����p$�	�:��숂���|��������놙~��Z���-Y�c��jK�6Ep�C�'%"�ʵ�j��Ov��5
�7`�*p���A-��1sf*?[P���:��WS稿�_�
���4* ֯n���m��,�AZe�c��M�A|�}39���; ��e��L������2n0���Ŋ3ZgW�#�|�����LS޲Jk,dЉ1�ŏP�f��A�W�p���7�����f�ptsmW�7N+ݓܞ�3�`~��B�ӊ��0���vj������ٻ�2>�������D�H�F��ʛ#g���
7��DP���ny�~�5��I���!�Nl����ʉp�򽢍jq�#@�t��Ϗ�����r��־����1���xV䜽�ޮ���7A͖�����b��F���B/;at��R�!��d�DU�ՕǗ�t�iBX/���.�,OB��>�ɴ���hEX��Cǫ�����~��1֪'D�vߟ�xy6�$N]��KR1tk����.�b��9s�w�G�X*�3�d���~/���Zl�/)>n�r�J�t�p+j�ˏ{�L�t�O���w��&��hD�
��K[gj�T�c������YqG��==y��������l������=�l���l,��#j��ã�����g�龾J�Xi�ep�b9�����D��-5 uN~ۛb}�Px�^� Zv@^a��3�)L������>໅�ح��)X�iA6���gkL���a�a�䀨J$����Nl��uUME�^n��G��uE�F~�0�Tk����$T�^���_�Q��i�d�zj�y�rs���s��eO�����9�qY��O�Y3�H��՜�37�?�q�>}N�k�1�d��M�*^����6��Е5�fLCS�j5��)?�8 �k4�vuC�]��':LpnCs�ُ=�Ǵ-����;γ��h��3:��r�o*��U#F��k�k�Q��氱p��F�f���N2�O�!�o���^� bk$^���9K>TJXf��V�,���;.��M�hPl���w��SuIL1�E<l�Ǣ!tT0��(�Ն�M����~�C;
֦��"dB��vg�]B��eՈ�D�����q�<���� 7��e�t�Y6VZ���a�10Ff}U�?�'z���p��pˉ�Q���,~*^����C.��Lt�[ȑ�u����I��)��Ȭ�y#^�&��/�a�5�L]�����G��$b��؃Ģ3h��
�j��l
묺M�t��'�y@f�r�>��4qAgo):�Y:<�Y��� �������$dĕJ5S�c@\�&�T Sh�.�fK0��vwXO]o�K%��X2��Ib��+��QB:Ų���F����<j�N9�������ZU�zv�ϥ�"�(�������0���r"��	Zo[���`&�Kn�<��X�b6��3)҆��=W\Dodγ8�G<�%����Fpk@%�%c@_�h�*6����˧�eϟ�EkGjZ1��q"+�xA�j���Vڇu#�w@���۠$�-����z�g�F�p���� ����Dw!lB�w�$�d��E��t�y�r�/Wh5F��o�kOl�^� S{�z7��_�XYa�$W�7�P�̽Z���#��<¢�jW(
Ͽ�'����S���d���!�}����3����k��IM�܇�;�r
��LO�x��	'J:I�)�^H��!��h�4�&�ó����m�g��� {�O��@�op��K�?;�׵s4y���Ү�EUD.��{�5�˸'?$�ǭ���U��,�y�Ȟ?�7��1C�9�{V�t��Ӧ�h����[�:(\�_T�3�ybւ$}����d�N��nk�8e�OMO�<��F e0N@cz��=0��y�9	�]�(�fj��	o���I&]Q����y��J���W���G�~�{l����LH��7�i����7s�K��ukq4;Zõ�G���O����C�j�u�4ts��a��Y�jCET���!������Ŭ�Q�tQ�jp�+D��>��l�4bS�aW��Ss���j7z 
_|�K�#,��2."P~^�p��?�ʯ���gWFh�V���Ն[
g�K���t�Ko5��G;���8O{|g�bؚhNx��0�,/����9�j��V�X�im0\�{[[���݅G�;Yi�٩
�4���o��zw��e��X�	3Y���Oӎ�� QZ*��wtP���n	B��dS���M��ue��⩿�����-n7�j��E�	�) =O9�Ka������3������ܢ��s��YQ[��?��=I5y0d9޻��;d���E�c���(ER��Q�.*
gl9�3<��6;�@W�?�u���D���ujPMHp�(����j #N�O_�oGQ��[�c��*drI���1�O�)X�xAp
 Rv��&x�B�''֜ǎ����V*1E��jA�8$�����ِ�gh��Ծ�Lm�����)WC���L]F�	��0���'��נw��b��ā�כ*߼yT� ��<�Mo��2��Q
�}۬�:ٶC9����V�҇ֽg��oOڒ�u�H^�=v{���t��Y��A+�Ҕv�l�I���pa��&���	�k��M�_�>��(�:�q����W9��0}�'[�q�!j�-E��e(UFѬr!�6x�7����h��:�Mx���K[���[��"������(�ɿ�1A� Ʒ��	-+AC��S�!oV�{�`��]�h����(�8"�\���R�*��Q���PI�^(��E\0��&�&��P���M��P!�Mˮ��t�߮�z&7�G
C�W"ۘ���B��'[EHA��?��iI����r�PT�a����S3Z5F�E��] {�͘I�N���	G��T�m�ПW����^!qU�W�8�8����s���gv~��~=���O�1G��@�t��>T���r���~��0oY�����!�����䤋�4���;���du:�)�����X�9pDAh��OWΕ�a���5*8_����tp��4m�$)��B>d�02�sw1�;�S�
{c�+O&m���T�[����JB��*�澸��v�H��x-��%��&�� �PA�S�^���D�ea�8JNy$a7�&��\����)�j(?$g�[�N����*��Ş:�E������Æө���*2�S���Пa�'�|�JLE���=
���C�_���s��� z%蚿�͐6��$-���DЃj߻�~<����~{�}ą{mԍzd�K�����e�D�Xh���ǜ4�t�ŕ�{�\jT���!4����c���6��$b��o5Zm������N��-�&�h�~f�LQ��S0��)OO��x�5܇:���h�I��k8�T�IU���&8�7ڣ�r��%Hy��r!���~�ĵ�"Wա�#�JN���ӝOP�W�����VXfb�q�Le��]�3��R���Ss��R6�ࢇ޵a�"⥗��r8�E�^��m̯��#�;��̹�`2.�@���LF��೬	3]Ո|��*�Z�H�E�`���mI�'Q��dv�#,�5�����f����ރ��ki]�e��Z.�j��,�t�x�!i��2�'�;�ª{���aa^�f�?ʱ�ti0�>�glk�󔅴ʮ�N?�U����'��>��v�#�b�ᘤ��|�؂�����Hm,���u�I��D�3���	6.��f��HP)��eȃ�� n��N/�ɯ�s�/؋匃wB}�=Z��N��(���rPq�_�fMe��o�،~8�Gg�h�J�����6/S�D�C<�c%`GQ�p��d6l�_Ȓ��8g�XC�r~|'���7�+<�[e8�?�&L���C�mݝ������u�P��(��(�{D��G?u1#�i�Y�L�np��^:�M��]p[�6}�J�a����B��<7���Y�SSG9+������@8�����!�7�lG;ݝ�[��nЊ��90�7(vb�H��w\��O˅y'̄�#�Ÿͅ)����7�m��<�IM ��a�2ȥ� V��c�;�۾T`g�t��� CS��*f��	U�K���kf�z�G��#B1HX�L'Wc�����&�Y��{��2�E�Ys,�m��S_)1�#�P	_�)�l��Q���ե�U0&<����>�JH;���2ߡ��Xv�����1y1���N�n��O�)֧����/XEM���h(�/-b@�A2��7GJ�ưݕ��ּ���>��wm������	֜�3�dz&��T�G�f�o�0#��[�HA���TT�=�/Zb�%j��u�N��'�U����'C�^�*��짂��k_�
UU���[6>�t�2G�+���͆�{z�[Y�K{�a��g$�7�L�u@��6"$+��	N����@07%ȗh�z��AU�T�� 5مAkr���Z²A*��U�+f��0���آ�[���^6.��=���Cܨp�#����n�C�V)��_.�!U���N�ui�ɿ��S�s���5�d5?Ԭ�=�� �;��q�ޝ@��m�������)�!ǹ=��P�x����5'im���0�X,����O�ԏ#�1;OdF�����3,ل��� u�����F�V��1�hI�u(��k}��A�&,O��s'$��ck-�BB���U�)�u���*3�潪������x4���)ve;ó~��fgy�ע<?����e(p~@T:c����������!�o��5o8�Xf<�cP�����~}4�;��Ye;kX���d���A��ԋͻ��5ɵj�:��2. �F�=;@�z�� �*&��m��"-�T�)40�!Lv�D	+ I�à]A���(�-�~�������N�p�����RCx�p�\dJ�@A�C�[%�67���U�QS�7��̙���S��`�VR��+CC�5�ˏ`�8��?�$M�ו����4$l��.���F^=b�����M{�un����uA�=�p��¡����a��P� o�)�S�,�dd��<��H�l�ƌ�@������
�8�0)�cyT5�U�q���n�Qq!�r�3�-�F���3
�%g�9iK�R~����	�>?�w�5�	u��.Q�x^���֓X"�X����g�]l"�@���b�<<@fn������6�8�o�n?Y�x����)���i���uE�ڤ���H��˰{��M�aVG	P�Ir��c�	{���O����}�0�fL5j5��?2�+��1���8G�D�g��?8��`QY3qHϣ^�FW0%A�(���T|�O��d�7X�����M_��귅f��R�JlST��y<�	g�R�Ք���<�쏎פ)KU�[��g���Q7�����O�^��V��@��u�a�[��w,_��	�nd�(��1O�}wu%qn�1�N��h�x!�	�	>.8��&�;X���-��aĳ(]���2,�W�=���Uj�ۨI,�������ҷ긖����/�t��i�3kk�(Jf%)�Km�l/Ϝ��*����l�f����=C^Qq9b��55�%������Ł�m5�FZiE���@9����9��#5��b����g�Ͽ�'�Ty�>�H1\Msߍ��Xo����1o��G`_��y���ڢH��&"T2W=mi��Y<��&���<�T\u��|��� �6vj0�E�Iu��-:��.�8���3aԆ 0��L��#P�ٺ�O�� ;�}:w�+��Vd@L�=r��O�l��)���|�f?]�,/Z�e]0�*t�s	�g� \�h
�	"��v�$��M�?ؓ*ͅ)S���S�.�����.Ϙp᝙T���󾆩�j�qm�Ja�H8���h�@�jN����<��wL�w�yw��Hb?���m�}:����O��!��!��i�Θ4�P-�$�z���G_��<�UE�hX�W�؁�w�[V�q$2�e&qEGv:4<�$��1c�M���i~�D�|��yb������| D{G����R�I�"�Z�bg�u�d�kU�i�w�2��M�i��zEr�:��pr�_����Tq�U,tz_�f#�6��-��Fj�'����������l2�ˇ"�W:Հ�Q�ֱ��{j�$�f���%�K�3����9��[N�����/<6���'��QE�Q�벤����s{�����,69>�S�i(����(n@9� <�]9�[!������Ads��@0�!����
rw���^���I����5��Ȭ#}B[#�z��eo	] �R���l�!�Q[�A�W��|R��I;�pm��ՀʪI>����t�/�%^H�'���t�o��� ^B�]Ͼ�~�z7{�2R Z���{�X\	je�r�T�u�|��$��0�Κ�ٴ5�LY(Ay����íul�H�t-H^�賴��L�V?�JEʙk�>E[��<�G�B�32�Ӌ�t�Y�$
��W����qز�e��;�;�p#QJ��2w����6��K�>��h)Kg@������d��$��Ǯ��+q��*.:��덶t�G�XCH���|0���������dBE<J���5�uc�}�i�~���ߐ5��Y�,	d�X��c[l��ݮݠQ�1��)7���>�1]s^=C��s�tz錔r�7���%]�|���6|�#1�}�I�
�(��h}�	sb�op�f۴l�T,JC�}����;����)r6I��' ��7��{���n,�i��Y��!�C'��I�>�HTqh�0��!��.iA���Lۥ!���\�%C����o`2�]�l�]X"8n�lCG��H-�؅�u�l������f���
����Q���GT7ƿ�Y�[3�@(H��)�d��K+K_E�5�g�T짟D��u�3rv���&��1�`
�N�W���iX�-!N�v�o��&�ƍ'�x�ղH�W�R$��{L-3�	g�v��V�k�AI������~��j����H�Q��	���l��v
�/��I7�Y�'��s
�>�j����`���(Wܦ]�;u�lU!!N�3����/)4�E�`9v-�$0���?�W��X#h='Ӱ,tke��ΞO��d��O�I�+�;۩M����a���.� �-�X��
�`<�f8�9M���%�^�G�-n~�f=�jt��;��.�p�S9�C�����
�y�`K����g�I�D?��U��3گf-` ;1бX^T���?�Wɍ�8�
b�6���:�g9|c��@ũBUD�"Ť���yv[n'4�%������&���UN�DZ�E����%5����"'�f:�W���ց��F�h���2UWS�1�+����x������Z����,����{�>�Xo�Y�����#U.TC?��Y:\v�
uV�w(W�A��b|��<�IY�ڭ�|{;)�?e��\6hJr��!�L5Y��y���A](���5��L5�HN��J�a�oЌn�H+��b�������{�0���}\��� ��������"�x'����PT׈�Q�B�����2Ͻ�M<Ci���@�k��%�L��d8��g�Z;RpH_+�a��6�|��V%��&w��/ݚ�$��]�E�/z@[��Y��:M%�r�s]ަb����9���f�	�̨��f��1�l����Լ�ԧ*�8<�ֶ�B���;�4T�RFMO%�M%�x�d���#��~�����6��E&DM���1��
w��빗m��2�ք�a<4�_�M�|M���H+w��jtuj��9�Hn����:Z�I��������i��&a�q�
�\�����`n���e�@H;�8յ��H��&�d���ޔ�(��}=�q{��0��j������CJ�q��a�ck�!X v��`��.��>��A�Ȱ�L_F���ƈ&�w��_��7�Ś2�F0�\���w:���O��!�pq���t/�xCh�U7!O����I1���mm�ʨ�>��� �F������B��n�ZI���*dP��`�Ha�����h��;�6�l���1h�[���c�g��N���r�Y��K��	<G��Sm���Bb�R�����7L%fupG��@0���*qXF�P5t���y��i�Mh�= 폎Ld۝c�Wi�������lKb�$F���5����'�̖�?p�^+�`qi3_�Ӑ;�M�py������s�I�EG��e�8>�r"`mv i�3�R%u��Z��4i�H���\^�*��:d�{F�/���.�义�Ov�ҍ�ę2��Xs���k���F��I�q�l�;腏�N"������@�I'6W��]�US�E����.'eVu��c��$���0��q���[��J�ф�#���y{�Ix�	��(�n\N�j %�f��I���4[����\U�b	��[�p�C����?D�#�hb�O\���z̨��P�����dG���z�G�>=(�.)�&}�����ݣ�����$��'�L�5zV;���RM5ݧ[j��t��
�����T�DhV0G��.�R�'�v:��n��Ú:
�r�5�Y�}�J���=�"���_�qcQ/���2�W����|D��*�L�^m����$||�C�_���JV��~���̥�h�����/t��p)�?��Ht�ڞ2_��F~�/�Smze�[E�bC�v�d���ƐN��j8Nu���R�ֺ�h��E�3;������[.�n��Q
��|�e����r�@���ۇ��ԉ�YN�B�����d�W꠺��v�P�i��M	�C\�i9��6�h�
�`��^�.�m�Z\�׀��R�,τc�wy�Q<F5`�2l�è v̫�ɵ�P὞��Ŭ�z��7#�����X�
;���9�O����hh�Vl ���M074H:�Ե�_�lL�9�z��2�V���O7�����tܞ���̮֮f�^:��Ȯ��K��r�v"[@<H�I���}[����}	��a�I��@�Y�3?g챕d��j�ޮs+��߱@��W>"2�@�MB��ml�S4}~9�SMN���6O+��i��%䯰EO��֗=�����WLt�?n�QU��o���ӌ������ǖ�mu+����ٞ�R�c��D��nzgU���d- �q�߳V��?�b�ب�=���Y
o������I�J��`��A�%�<�c�X燐W3_�G���w��5�8wBEx��
iĹ�LkpZ}��/�1�ra5 }З���`�>���}�ON�r��Wj�q� ]W��H:@��j֋zP�qs�?����:8��|.�ĵ�p¾��G�T Ӓ������"7Φ<�\Y�5.�6���gCN�
�W]6[���	]/�^zA�@s���
U.�!dR��o�"���O~�l�8�$��ܵ�o�M-����O۝eg�Z=|.^��m��Q��]�n'@R�/L�j������];{�=`�3|e�bR��Gϗ���(TL"FZփ{�Z���P�� �ؠ��HT�҇4�����+������#��A�ȸ��>��kA��GnPX�S��G���9�gZ�lj^���sѫ�o�<�j��QVCߑٽ>���ʚk���o�6�+�M��q]����;e@��;ד��B���e������\�I!�_ըR�zѫrX�f^��]��
�ҲSuoZ)�Ssc ,s���Ua��<H�.�����a���t��L�Oa���wli~�O���]�Ӥ����S��2��4��F���]�F�t�7ݍ3����!��A@<�P��1^�������n��c��rk��y'�m���/DJ�GՁ	�Xø��5��Tz�\���e)#����ߣ�<�D�Ӗi�_�eN�W-3��Ͳ�����[e�c�V�3�h�Ȯ��zv3d�B�'�H�S��qZt�3[1�����8�G����H*уU��@�C��E���?!�;�b��g���)3�2�4[�e����]�W��09�MJ���*�x8��q�m��|�E"&�d�����AF���$���g�Z��
���Ȟ;���}�h�gR�������D�W7cw�T%6����`��KCr`bt7��#��{��Ƣ�\}�n�F[���c�f�"#��M�]Aw72�l+��NG����kG�����j��f���.�ͻ�%��Oo);�D��%&�.m	Ү��5�8"��!P��ZN~ON</�v�S��u0�-�k.�?�ғ��9��AX���=l^6��'D� ��K�%��L�Y���<a���c��hJ�ސe涑q�8����C(XD
�x$M�c��l���s*��a��1�����������k\�0y�3��$�`�}�_��F�ٖ��W^�
��\5���v�w�� �oT��
=���=���{(��x榹N}����  ��t#�j������E���Q���Z������5� 75��r�˒A���M��O[	� �Rq)�z��&���[ �~�����l�'���u��*l�)� nWډ����'PC̘*���(g���o���T
�Kp_=X(B�<;�+�n�ĩ|������c&��l�ک�3��Hd?�g���3	b�!Zx�6����̷�-��	��uN0_�碡�tS�q�Ģ�Ha������M��ւ���Vs>�u(� �l�	���y���4h�Y�9�3��椿?eF� ����krn��i@����	ip0Cc��V��E�5W8*$���<���+���J�G��9�IR+����k�4k�;��f�<e�
��:�8��sM���f�㦴���:�[u����ɞ��(��� X��~��מ�1�a:�|�'��]�D��7��'���Cm����w�[���w�RP��{�_z'�-F��Ԡ��P��
���7]��'�B3|#M�]m[{��G��:}��Wvk� ��<�N�(t��9����(��6A�aj;��3~�ͳ1b��ͼ�5���A߿Ih[�"���lrAZP��*�r����a��U�](�>M���+Q����ezJ󩡅�����}u*���{*5�+�F�+A*kG���=B�u���7���8.`%�C[I��*��%R�)P���p'�����!C�}>t#���%�f��͔����N�!�|1y�ҺŏC�\��<#T�Eh�Ok[k�.�9�,�����c�IE�Cؔ�Ôsp �'����^�;[�K���gO�>{�z�n?���I�=15+N��R�=�y�I�U0�Tmg�d߃�-�0c6%N1������3>���1�߀�c�$�T�s<��n�Ms����л��Jl�5��p�*�s��D�h&�Yİ�;�h�P�=�@��ü)������Ni����(�J�)ת��IHU�54�д=�����/���5@N�^�kٗ�o����I
��O�����N�3)&{Z]U����`=��.5��̷ڊ?���ntM?���.)��80a/<��ڠ��(o���/B]�'2t�ݓc�^��Rp���%�1�ԅ��l��iZ�g�'cǅ~���ϵ������$|�m��e`�Li�H�d�Xs��G���f�2��XU���g�)I��	��3�^�Kq�?�ecX��ɍQ�o7�ɮ����ָ �֌��o�U,��-Gr�y�ג��j��H~E�Λ�!\���+q G�-��m-��-e�@�N�i��e����0os8mЉ	���K&�a/��&�#&���Ḳ6U��`�n�
�*mpo��j��)�� Ҷ��Nս��������1�c@�1ٟ�͸�z,�)���k�<�b�R�l��]���)Q#� �:�L��H�=�%Q�F�����>
73܊fo2r�,7�̰GᜄQ�Q�O3d��1��E���k�����/�^�c'c����g�1�߯�_(��怷�M�O�h���V��̈́ͮ�ؿ�X}�Ŕ��τ����}7�ϑ�xt��uƽ�V�M){$Y�ș�b���3{jp���6���}u&Ny�?��qY]c��ϸjP,�W��Hw���.��9	i����]��ᕏ�����ѣ�e�Ӕ(���g�=R�i!�NdQ�F��B]̫��	ή�G/=��Eʕy碲���Y*հ�}:w���mNy��:�"؇�5-:�~A:������z���њ٬p�Yq�'wy__�Z:�Ls��rП��m>�WJ�),6�nL(�X-�����ܭ���Ms��n%��2sC$H�2	�C.�ALţ�ffK���=��L%��Dk�J)x; �ߞ4RDQ�=zb�H���w�%��n���m��՞��*�L�^�(�J�cھ��h8�Q��p���@����cxO�Ww�b{M� (}���j��^��r�S�N�Kc+T�ݏ���������b̡��|5;�2�U��=p��L��� D�ۏ��@����˽�y��9Ԭ�;1��'��m�7��\�L��AQ ��r^�9�x3��o`�I���7����+��;�uU�����9a��䨮�=jHP(qh���/H&٭��y*���v	(fH�W	¬Hp`:Yъ�s�(K%�?#�d^=���8Z�03��8Jy���Q7�e�h�6y�p����213�+�2-@U^Iӝ?�e�=N]i{U���æ�_T�!���p΀}]��}T}�}����o��=Q�1(�ޡ�*5xz��8t�6�3�J����%�-�,Ҕ�fE%|6��0�2�2����s�	h���]m��{�(Vԋ��~|ț��$E����+�/w�E���<���d�6��eJncj
S��.5�h84;t'6���rR7$����G�^�.U�.9�'���'���U�\_�E��@^KEk�C[:@���&C͢~�?��*��0Cݾ�g����܉x��Q@�0,��s��Fm�G
��&[!��n�_cE�����j�J��v�JfI u�^��v���]OY&���^%D���[&���I��p:�Ra��q}JX|c�J89�|U~�e{��6qRU�WU5��b~`���N���!-//;��K��Y��jJ<��$�������a�����0ly,d���D7m-�]�Ka}'y�ҞH��fV��Ĵ�H<��;�;�\�r���"���t����O���=�͕g�x�9��6\g�=����U]]%+ �}g<�)ѯ���<�b��|I��u����Y�UJzMOd��5�P�F~s�/�����������(ʌ!��{�������	�l�$�Y�^݆�#	���)3�{�m�}�V�-�H��ÃB����Q\-��O�]�{��d^�9
�D%�
�LB�S��TO���E�0M�6�Fy<���Yc)(M�v�Jd\���+��o�댵D�Ih����cΨ����y脘!f������&Ub����ye����Uq#��U�!I�nh,F���q� ��PiB'��[S��Ҳph�a�Lpڴ4�l�c5]m=�?8�f.2��9.(��ȁ#3fT]�bb&�����T|��3Ӯ��U˳�C�&�5��"~4�,�<OHv�y��@[z,�[[[��0�L���\=��mD�(��D�Sm��=�Ѳ>�]�QY>���;w��cW�<��5�N9/ms����<p��g��q�&5EZ0��!-��A�m��Q�zx\A���
 Yr܇��hn I���*`6��s�ߏ�����Y���k�շ&2u80��} ���2�,�~�V#$�kC��Ѩ�����܎%^f�Q�N������EN�@4���J@��O۪�� �>�r��������[��K�.���q��K�Q��u�&�v)M�.�< Xo�E=�4nu�$X���T��
��<v��I=�k�Q��(��H��!������(u\��%A�Yc��!�ct�E���^����s��1֣:&��[K}u��(�Hi���+t�2D��䏰>�߁1\�Y����p���{D�'_N�9éү1�ϗ�}�`fs��E5�G����1�f9�J5��#N�X�����6dO��FS2��l�߳!�!��:T,��C0I� =5垴
Ny-�%�����>�iP���TbB&�y�tU<��������1��x~���⾕�����U2�I{����ጚ�;�W#ʮ%n���c�pd���ڛ@)�Yd�[`Q5-~2�Q�����T����ꨡ��7ԅ�h���٦U�^mG���<-���>�?t�%��"�	TP��v0��s�#���O蚂o�Kf7��c��b�&�ǹE�(~qN	l��k��9�Ń�n#W�g&oA�H������:�w��t�w9fg(hq��r�>`�a� ��^Y9�vi\0�A�c}�"G%桧����=�@-0T�eR�7����J���8${[�h���{câs(���<Mil~��}��@�Bn���q{m9��zZJ)��l�=b?�%0ފl�dH��#&{\�@o =,Ty������,T�f�I(�У�*��V��*"���+7c�K�bi@?/�ڞ��=�NE� �H-,a3}_�v6�2�y�p�.,�.&����mI�����(����?;e~#�-�T|O~.�ჸ�%5G�tǽr����6��I�������,=��d�ú����{��̆u�]6�%�Y0#W�`5k3�I�"��s͜�[�C܏L�W]���Lm.\���<����KA)�Z�6�M��Zc�'��Oי�g�~��
���;?�3�P�o�
�C�䂦'�h�ڟƩ����rٯ�f{����N_rT�A��]����3X ���l��U��)tx�8������@E�Ch�����Jl���V�9/;��Ҭ��pA���{� 3�� ��כ�_lj�v�3װ|�z�9�0m~�(7!��a�~Z}���d�Z��p<-�iZ�@���@D�`�:�x}����]?_ �1��[s����E� ^"#Ԇ�E�oݖq�g8���̩<q1�J5����w���b��h$S��.��G��vk�+���~���OnD'�P�G�U�D��w���4X"O��5!�k����Q$Cϴ1�{��_̑xr�f��:5]Q�M>��>�Q|���*Uv��(��-���ﴛ���@�~�Mǰ�C�i��A�ʻ����%35��!9�{������eR'Z��nL��Ë��m޼s��ƛ���T�(˧��o��6"���U�؛m*��ܸ��v��'�)~�1/l��#5��nS�����1{e��4طx��Q �zz��6^�H�<�#P2��>�ؼ��Ģ~��)�B2=H���)Y��ET`NBƩԺ�a�'�1������cT���l#�*j`����$�d���c�I�۸�)�C�L���`�im�j�"t�U�Ǡ��_��IVX�,,�͒��੨���:�k��2���" z� �nW���	���)�@�T�@U���կK��%.K�������$�	s�'(���Ъ��)��4K=<�ʇFy
�#dv�No��옎(hi��dS}0j[CU��$0�Z{�%��g'�r![dkN�l*����'�1��k~�ן#8#'�-��k�!���Y��im�)j�
�"��/nj�ᩯ
z��5����W;�+�H$&��0�j(�n
�7���3�E �r��zl������K�ݺ��T>�O������7�<�'9��&�
e��� �!�߼�b��\�#���+�S�����!���u�,�O��Gv�%�&l��[�����y�,C��p���쥚�V��]�!�Mm��A��p���+���{�g��NȤ*�����ۀ��/��oT�7��oN�1�~��(��|h�h�*R(@?��@���`��͝W`Q>7WI��h"���[��]9�e�20�c�����S�����xx��6���	��q{υ,�����tL����̞�a\YZ-�][���߬�6�����P����3Q��Ve)ŅV���
b�v^j��|}�.��y/I��Ji{��һ6�?LԜfY}�f�5��c�;	W�6a�t�xj��oAbW=#F1:�ϛ��x&��%-�h�}��&h�7�C�z�[��0�Q��	�~n���p\s��7���y�F�Z��um$�=�&�{�	>�{��VyC��)4
��A^5d����k7�v4�ZYp���O��K�	X�ip�����{�H`/;�r�@����\/8����k��A@�	���s����Q�A6<�B���=f��J�� ��KѦ"q]J��`�����Q%O����|���N�5�;�3e��c�EX�&����o�ӆ�@c�L.�C߽�7RP�0�X%���:��䀪Mw�T�~�ܸ�r��cN18w�$-~ԂH[��Zb���*i��R�p���V�0ʍ�s�6�!&%�X7bT��J������i�Te���ee���;o���5�s�)�J��Dܒ�z_I�dc���;���.���ʛ+�%��j�(�lC y^��v�\Y�9U7q�^�-H�b�Oe5ӂ��=�t�����I�K�Lj�)�%���Iz�F.�(^l g�����]}�Y�

�p�E1sF�}o`�?	�K��ۭ7Z�L�LGB�D~�k.��	zf#��%��@���X)���4B	Va���6D9o�Yx��Q�iВ�U@�\l�FȤ�/����f|�&���Ҹ2�l���vf؅�<��1�%����P��$�ME(Dg	�0��z���J��~;	�������v�qpf��'� ;0�1�D�F�{�F�d�ndO�F�5�Tu���o��pQQ��Dqݟ���ӆ��ɛ˞RPZ��vØm)��'m�m�u�3b�{��C9�$T ~�L'��z��4*����P�]�X���a��,ֱ�Z�^}�E��݈�gw����]g���q�H��C�mZ�{P�������h�f��7�y�h��AN��"�߭P��OH�R�_۸�rzLbe���ϏC�k��E3FT���K�3����܏�'�x7����%_�R�
��P?����}T���F^p�!�	����_d߶��Y�����������=¸r��|�I5��If�=Q���I���� N�A�3j�\qT�PTdC�Vq͕�&���-��ڸ���}��}+(�n�UC�\������b� 4X���hF�����V?p�G��"�{�)mcA�Ei�qļ5�yI�n0��}�����v��aC�3�x��,��i��S�O�R�QğK�n���q���R��F
p�m�Z3����>`�R,�&S|����,"���8u��]�^�pqR�>A$`i A1t|�f��q����n�3��d�GN1U���Ğxa�]	�v��}�u5̸�=����HE�zui��x�8�*�wB�ϯ7dj~�@E�N�_E�}��C�j=�����XzZ<�z�/��-`G�!� �@�ݚꂊ��=EDv�F{f����tW*�!5~�J�NI5��@R�����_p� ��M|�Z�y�4�a�8�[�{��t�73�|p���Y��Ɩܖ�Ī� :����ġu�t��ޓr�'�N��ytRW����oK�^U���|��L;�(�V��1z`8��x$�'a���ٜ}���f�~S����\18�=[��Sku��8z1�nC>�f��}+�Z�}̐WU0�Gf=�Y��I�t>)�=WL�<���!%��T�dߖ�D�Y������E� O�͗�,�x}�^0*�C�|g�����/����A;��j��,İ���Xӭ{�=�˔)���- �������#�W�%��T�#�Yni/�1�0��n���-�p���d,��F)�h�ҧJ�sHd[�!��T���\P!s���ys���N�ϧ ��0RQ}�n�H���?�$���wm��v��}�m�s��yڇ��c�*�QO�&���竷BV�^��A�]�z�q���B�]d�,U)b�Wu�EUާ�|���g�̅�LlM7+12ѧ�u����غ�S������~�e#����G�q�Ǯ؀
���<��I�Z�=&��VZ�]��-MaT����P�A%yB�F��X;�V@a �S��O��w�N��C����Y�#֢:B��
�o�x����Y�E��c��fr����38%��Ζͦ����� �#T�<��`��2�3��]�g��T2�U\`Z�	P�j�mj2Bp;}HJi%�{�o�ӹ;����(���KTP\�b�<���̨h_U������vQ��)Ί��{\v�-ot/�t⏋Osm��ё_d���ռsve�B{aʘtL � !�ݺ8�P7�2F�aI��9x��d��9����7�15�������RmJ�*f)�_F��Z��֙�{����ǵ�v�5q�͐�bW=���b�y��l�����{���_D�0)�0����g<�d8L<�1z�����w���
�;/�qY��֮�Tʬ!�G�x�,<���Ou	i�!_[~ް�,V���R�ܢ�]��D�:"���*�����dx~��$LoJŨ��_\��B�-0�B倠8Qc��M<|Q�Ga�n'��t���s����@������{F/�k�K�ɫHAng?a�z��?d,t@���uԪNJ��"�R
j�Ү*��bQv`��70t����w��lc�=�/�Gxޅ9�p��If��Z;ŷ�]W�ɯ�1�:W�A�Gi�E����F�6����?�����a,B8�C���r2�[GՏ.O��@<�V�$[U�{����x�X��S{��a����4�P��(�������ALS�`�ή_(�]���v���2�����h���2��\$E�>��s��b��>�4Ee�k�Lۢ�0<$�v�v��j�mz��M-������s�1�M�Оm5m.	�}O�1��-��=;�3\�#V/A.�j�,QJ��[.F�����t"vB��
�C*��t^�OGL���Uf'�Z/1�Afá�}{�P��3<6P��aO�C�i}GwtY1,����DAy�d=3/;��c�$6�)�6?�
R�Fx��q�y����{�eegB@��)@�V�-g�O��h��*���Dp�w|C�g���M;ƔU[���~V(�uDC�u0 sO��9H`��Βy�L�'����!�"7���U�A@D��!�,旍������]�ƈT�%�!�	�,�B�R��90l�wbB�^E���{�����?ͪj�"c�YN��Q�H0�)� rz:��e6���#xt\�qY5��W���U�T9��G�s�[���	%S��W�	��#,��ʰ7#�`�ϮK��l�u��8��H�YǷI�c�ޓ3R������M�d�{B��� pq�=5���$ ���'
�B��N�B}��h��Y���]���1?����-���}�����R��>�!�%?3*��X_�?7)(��ta �!�c�u���ݕ;�nV��E�&��~��)!�dh��f�W�7c?AV,���G����|�#����Q?�0Z���Z���DhДj
��h�;Iǐcv����_`���֋H��U������9xA��H�߲�*��C����:#�V�7D��L0H��圑8����*�K٧��ׂ��u
��"%��U*כa;5���c� hhe�r�*���w�w��A��m�Å@�GX���X��Nl"����;���4��쨅?��@�N�aK�)T��лO���`����<?(c���QE|�@(A?�}�~��pn�x�#��ri�ҫ�2,y�<��U����`X��U�:ƛB�LlR�:�ޚ���)Jh�I{7����&��{?�^n|@\�?+tg�̲Go%�bP a�q����
/2kI>L��9{�N��lʽ�!:� rM��\N؛�\b*�ٛ�+�rC G' ��5�|/#y���+�Fc��Ư�w�3^�(��YjM�jt�%[�Y
Y6A"�b0`���M>~Y���nU��4N�M���8� �Ժ+�Qɍȩ��sD�`ѝc~�Oh��Rd�3,�>_��2V���A%�Q��Aq��Q�j�\ڞ-+vubц"������>b�,Q����`���mU�����z���(tTA�vtc%��~d �ai�+*������~�ӹ/����!�7�)(���8���%�,S1閾����?�[t��b����]��b��f�iX@�*��5��ժ^��^w���(���LõB ��K����>=�� )��M�� 6ڳ'�.��d[z�ǃ�WC*���;XQ�I�86�U��M��2dG:�#�Ge�/���9Q5��a�ՄLFF�'�'L/�q��HU��>�Af��'b|(���W:m����w �R�a$ʢ�rC(�
w3Gs��<-_�d�[���_9r�=N��̥(jh����!��|�`邐l]�K�����w�R��D��Ud��Ir�Lc�%���Ǯ�)��Ͼ�y<>����L@1�\ۜ��?�C�EŨߟ2���M3�H���lX[}^�ۀjͫ�����=X_֜ԽﮮL$��P�3��I��ǴY��4`�8lc	g��3$'�,�W�K!�/j�@5m�EĬ����T���è�
y�a�9s��{WY��y�@�x� ���Z���0�`5]�l��\@��I�����9�S����Q=>q�`��7S�k�rڴ/n`�3S�o����$d;�(�*\������ۢ��ť�g@��s)i�=��{��%\�AS�$���x
q���+�X7f·�U#���	���hN�iɴ�������;V˫h���nV��'�6(�}0�Vә>�Q������r,ò��SSzHs-��r6"��.�G� �ޚe=���#t!=��7V�mB���[d��獯�B����{����u�C�簍Z����L�ѫ��;
�b?\2�!��ـ�����ڪ@�`��AL��:J�5�cmp���Æ#���ȑ*��h׊����s�ժ���؍t6&-�?DO?,k����pk �h�N�K$�Ƨo(�7#�$:���_��l�I��'�_բ|�Zրn��������WP�hů��̜F �`7ҫ� Ac4���!�m���#�9�`n� ���
�&��x��U������s��e�wz��f����DNR
� � ��D��ל��{� l�!�Mݥ��#f+��>
�V���������L��ƹ>!9?\j�,)J2���j�{94��i��w�ns��O0n�=�S�ԄF?�W��!NadY	-�4���i9e	̞�ig��!}é�$�V-�*y�C��j�dh���h���z+
����/���iN=K���T��bI��d�r�7��� G(��d��"ڧ�����*���6G��瘎Z*��(�-��$Fhh򈊆�2��)4Y�67�c�4 ̿��i�=vs"���yj ���Fs��O��R�Z�/g����@�a���i<���m�����Q�o�/;"=�GY_��*���J��d��H"�mI�"�JR.���L��j��͵p�,1�(�QeeG=�z���)g2d��?a�m�ƕS�ۤ�)u��_���^&E����1�SϨ2xs��ɣ��8|(�JK=��9y��tI��'�_�+{)��Q� �&�����m..�	�'��eE����h��zO)+-�V>*�_
ߴb\I�Sh'm����Ц���ҥ�{�i!m����d\���
�?�Ԩ2����^��?/�;D�Sx�w�y��ڗ+N�ko�x��O=��_���G(FA��0�כ�g[VIľ�Yc<&�5rm�IsaNVT�sb+�zY߲ ��������h,�Κn���)�^䠹��;�#u����WN	�&�x�%�3L[����AQ����*<����\:Y#�(���
2"}��%��L������9g4}DU��W���#��X
[ ��,��}}����\�"z�߉�6��qV!�7��}6�5��~ ?�6-����+���t�G��8�p��d��ɽ�Z��\QT�k1(��F��w��v�o?���a:�h�{�|��f�m����V'K�tk%T�:k����pq  �ٚ��>Խ���i8}���Pǂ�Q���8�C��/ܰ4��~R�ߝm���K��a��g̌#��r�Kɢ{9K@'|����b#�ޮ�}i[�^c0��#O�s�9@}�cg�%_����q�npzm�6�X�/�H����ai��"�m��n;�j��֪�دiCz�plV׾
R]�*J�)��5���J�6��Af���D�t��z��S�<�T�o�#o���9�Q�#$<c�u*^n�T�8�<;��/���A���_`���I�J��g��7�㨻3f��i���(S����_���tgQf͓�Nݏv
��x����Z]�v���T}�~����-
`o�z�N{$T%zr�C�n.�����W��&�G�1����O:1�U�ä��~;U@tL�����6[�	�u(*x�e��%��ߒ�ljh�i4l> L�ŷq{�JSm(�����!\\������zG�b�
dyO�Pe�M7h�6!�V�$a�N.��2Dw{�]Ӳ��QĹ=>���%��(�7d�I�pFu=�G:��:��f-D��mW2{[F]k_�'��u�+�&����իW#���S�{:����r׷퀸8��oBl����؝�H�z�>}��w�iC	��(��F`��8�*�TL���x&5�Dp�Ѷ�[��҇��s[�K�r&�t���T����-콵'0;��Cfd�M�}U�z���{��>�B2ޙ<2�|-��WKd����W⻊N�� 4�WK�G&#�z�w�Z�F ���0XOmc��;��d�;�@|�WΚ�5WG���H�U*|�;X�[���.�'n-zw���XAꕝ�R�خ���(�Cvn�AԒ�>3u9 ������7hU?#̺�z�b�0����=�7&|�/ש��A;ߞ6���0�$��d���ۅ8��ɹQ�pk
����2I�� "����H~�˲ۻ7�?7�+��#�$�@.�����*A��0�M�r�Ǝ��x�Q���>G�
�+�W a�ڎ�A��� G`�X��LH��$`����80+e{q��Y�����]�Q������w}�M��̘j�!�U�@`�֐ԫ���*¶���|@P8do�u�N0���r�~/>|��Su���tk�Q�h@�����0KW���:n����9�G�z.�e^�-�O�y(�ֺϠ�VXݒ4۷pB�.�Ԥ��c��F˼��iT�W���iK��	]��z
1k��и�Y��v��kQ���O�դ�D�v�51`�Z1�[�"F�U@��$H��_���z ��ݠ�A;�4�L�;I���l��0�O"�P	L��e��� ��P?����V����"L�<d7&-�-��ΰΡ���/X`�5K��#��+��a|�.��0_���Ho$⎄��٥k�3� 	ї�ֱ���?�*��mbm/�0����������KO��BU�W�i�	{�"�$-c�&N�0)�y)r�O���<����㒥����(jRq�{l�'�8�ɓ W���%2��8	1s���~����"��<b�^(�ۇ[[L%r$��D�f��&��eڻ��?��Π�����n;�Cx"c>�o���$����OH�R�ހ=5�k�1[޼�
:M7�Z�m��v��C�q��כ���5��y����.��Ԋ�KXH�I<X'�Q?�f$bIo��er�m�26����}lQ�Ѷ
P%}�H�3坅[�⿼�7���2pĴrWG��w��h�@0�-%B�7Ia�VJ����7ܘ�R��H�/M;��aD!� ��3�qm�ڢ��t�88��(�l�Ji��5�8^����x=93;�ۏrY`_�S�;bd�f�S�s��<¤Τf�7��Ky�tXc�S���b�N�+�<}A@nh��{Ef�Z9-��#���QQ����!�����r�
�s������[lVaX�DV-=
��C��J�V��������c��D:� F�@�L�:�c�����񥍒F
V��M��	[����L'��&[s�djP( ��^^:����2��%f=3�2�L^O�\��4��:����+c�hT�U�jV�:�����'2�F��$�8�Yn����HK�0�#N.nSH�����U�I\��ݿ�����@�3�M�|�W=�OE�ÞQ/ "�w
&3��J̨ͦ�����7:�x�D��2�s����s���:2����;�2x���f@͍N)�3ə8c|�?��c݂��u�SDƽ[k�UfK�����9�"V��HP����'����fxė�E����>�S�r�'�Jp��g�0����3WS6�W��7�
�F��q@�M^VHB	u����7h�Wx�.��O�#αc�ʟ2���Bk�_��4�"�߹_�7-К����q��"�DR�R��Ā���i���J�@m��[�����P5+A��	�?H�`W���m�ۙ?}�|�ui������&�����SOJ｀i�8�S�#HW��1 K�Ng���.����4㊉�Y?�����e9���S\�_�Cr�S~C�&��B�inpeɃD"Ƭm����1[���,̆����We7BOX�VI�	WG��S(j!���k�3.�$�"�:xkZ��o!h�s5f��ib
�5�r�N�:���&�F6Q�rb]�;6�SΠ�S���ŧ�;�����������H&�r�Ê{��f�,�n������x9D�T�^\"�@�>�]��BePמ����C�Rx���ϗ:�<@.�%�?�p����H1�� ��@$Œ��`V3�*�HKo&#t3��n��SHF�q������̴y�aY�$�7��̻ RF��:څ�?��8�Ð.&��~#I�"�PKh;F�OX��h.T搼	��ܣ�qY��ܟ����,DK>?����^�*}�ҕ���(˶�kvo��s!�}E�O{��8&�4n9���{8�]�)�F��{Vl˔�F~��!9RIp��E@�1���ސa�[P��.��t1W[���sZy��c�)�hׂB�m����`-�b�f��$�����$nJ��������U���(�2'f����~Tx� �b	� 	uOPJ<���&�B�����u
8L���( �|8!�L� ����dQ��#�R��
X~����4J��wBgP�˛p$ֆC*��^�JGt�(��N0v��k��V8����� ��j����U�R��{U���{�-��r����R{PD���(��~zB���0���4�ҁ�H�W�[I��.<�I��n�&�}|��`�OU��t���$4�=�`���݆ȈE�i�d�sK���v���-Bc��T��7_��r������-�vZh���H\�%G>��*�s4d�{ִ�!���,��2��c.�OY�U�bĳ@�9��xy�W�GO͆��
j�ˑXφx�@z瀸��N�� ��S?;<�s�4��k���3�f7۽��h�1���g����A�M��)��]¿:KuWTأn�P��?���(���ǎ�@�򬠗�B��nI��)�_S�f�
xh�Uݡ����|6���EqN�)x/h8��"5�Ш/oU`ȸ��u� �#O��oW�E(�;��j͑٢�w�tF����
��Z#i�cN����n���L1��SU0�J{2b�N�F�ڵ��4Yߦَyx������������L�9�bC����3�Y���p��Z�Ƶ\��EM`�׆��?E�W�UtL\�:U#z%m
�G��=�<����8*����̨QM�Qߦ�' ���ބ�>����l�@eu���؛?6�X7-��=�O��o���(Y��f��h�)=�"I ���(�T2�����myǍ#t����-�3��t[��6�¨E�nĪ�RY�n(�v��Ӭ���P襰z��-��s�l��#�z�L�H�1��kz��I����o���6t�4�.��H���E�� ]��iч�}/�#��sgG=��Imb��,���[d?�U�"�8�BO����R"�}�c�L�N�4��?o#Jb��d�#Ϙ�|��ѐ&� � ~�61�[,''��m��H6wV���V�{V��@����#ܫd�()����-5�)'x���,� �����H�[B6��ߖ"p�z0:Q��i�k�\_���j�|Am\�Ht��T1V�O��h��o�����A� �g��)��	����@N��ӋB�n_j[�+��O���4�ݭU?��"}�<�0�@F<�dCb�H�1U_ɇS;�X��ʺ�C*H�rWS8,�%�4���E��^�^���}��!<��lq��:b�(�+Ti�t��e���|67vN����騡*�*}3����9c�l{�M����?�� ��4��d��0�j�kV���Ήb�q�)����<@��"/���5
g(bQ1����{����B^�
�������Xt�vD����O-ëvhq��ܱSiS��O��k�����zz�q8��gRn�H-N�i��E�{u�D�{s�� Mr�0����*Y"�E�V�x�3��d�I��"^�Hk]����;�ܢ��$�j�p���:#��	VO䉬`
�C��#*l��ю���/���:��̊i�R�>��^g����7-����R3��]Ӂ�ř�E'�~��ם<�V�P&�g���P<{��2�.���C�H�<���\c�|����7�j���D���Tx4�@�3�H�
�I�iP\�Va�9����-&�����t��Vz٬���Y��_��r�Q���/��G����c�uԀ����q�,~M�C�,uFj��5̡�&���"j;39E�/�jL�D�����Ы�6���L��J�*�H:��8bZ�뮳7c�RDi�;:�>�uTC���
����k����ĩ�cw��mi�.Tu�}�}�{���RtZ�z?��e���gE�ܿ��������!��G��ƅ}��c�d� }|sm��-�W�n)�(�&x�����mav?T{��.-T���+ �h�:=琩��H�p�,b(��(*���t���?�\M�t��?b�$��	�Ǐˢ�Y��(������?yD8�5q*������B�lm���bϿq�P ����ج����G!e�J�C#�.x!+JpD�"�j�UT���Z=Ղg�2���K�%d�y��x_�U]K���}��c&�l@Pt������k�� �8Hy�]�1��j8bβQ����"�0��$�dsl�m��*n�{z����PsSO٬� ����+�w}@;8��!C��D������.�ɛ|�?r������f�sr�ed��'�F&�wf�Um�3�J
B�5��H�%�;~A"?��?�r=z�Jm.�|�,�;tjҚ�[�<�9PG���`�� A�'	Ũ����?a �wR\���<�pl�w��4�o�Bd�"����xi���`(	\����n���f��Oߐ��v����)`�L�W��P��������t{��%�躣�|I\�ƭ�;�=�*��Bb��ȩC��uq?$�p�=Ag}P�uu��g%�0 7����H��m4��t�Vs��s^|��SVZN�S�`8[�o���@6�`1!?�p�ܞa�X]���>g�e�j�?{2bc�*��ζ�BE>�d�^bƇ�1KR�ůZ[#xL��0�
�q�*�<ɋX_̠sK^i��C�P<�ـ�F�=���˹�SK�_�
�M��4� 8����~���H�E��Rv��p��� k飿�䜰�̠�k?"���)Fl
��ݺ���,2��57��|���6�N��L9p�����d��҅�q T�8��ɘ�XrC����?u5�$3�ݽ3��~L�*��?�����r�Lo�p,��Q�X��XxB�����io�u7Cs"�;9���y(���ۆ�G9!��p|��QIhs���M�qm:D�B��Sͼ5�%u�fW�Al��Kƽ� @��aKKK�!�T���l��e�ΦT`� 3{�ͮ��U����� l~�f%����s��k�30�WN@?��Ց��Oe���}Yۘz���gШ��O�s~�W-z�KH��p(� �W����֓��M��V	�)]}-$�ۄ��(ImEYyK��|K�����D�IQ`b�nE< ^��;۩����h����3]ª���j�{�!6�������ۼ��m+q�&�&�{������� ��5��q<��Y7�o�/7����9��I4
���_�fW�'0����IeM��"�:h����k������V?�˟�۲��!��-@ގ_�"J�K�FT {:?T6���Bu�/�M�ܪ�<���jP+�Y�z�Y�ڿAӕ&خ�if�����Rϔ��i䬊����U��%YP߽����n��2����t�^"$��Q5��&d�(e��6�I<��,�|ކ�p7�ʙ��k�(��-���N{1���.�a��������R�e&���(�ٟ��'����J,���y��~�R�
y��F͚j�-ߎsk�ѪQjYp�<�s���Ｌ��3�s)���(@(�C�W݃�P#~�4��Z�f(��!kէz�R1Z��K%HP7��*x��>�_��nO��DXVrv�+^S��B��q�-�7I{`�����q0Y|,��p���@\vNtq�.�h��,�	���h�����Adh��Ō¨��g�R]��?���^�p�/��.DC�M-4�D�moq�hAb��N0h�'B��+�ҷ���A�%ݣ^��Q��CB���x�E����~�����?��ya����2�n�D�}m���%�l�������q4��F����}F�o�}>&��*�p�>xw~\��4���2L�a(�P(�%s�����np߾�I)�N��bRc\Hf``�N �qt�R�������a�g!M�%���u��C�T��?���Pr�~��q�.�K�P��Y{���Yת'u팅�����E����h�������g���{v"�p�߄6?�U��s.��"<!��x2�٤���J>�c���;Z�[-Q�Si�$=�o�yT��J�<��������
e�=z�y�82�C�&F�z�$ӵ�0P��T�c��
b�\�G���\��I�� �V�-������ɾ*��Ŋ��p��D���ܾ������8q��ž	�~r�6f�w���y�}�n࠻w�:�8��n���'7�n�r�z2@�GS�UՕ�V{66�.X�S�y܍s�%ɸ�Nۦ�j��G&�G9Qc/��Q;�ϰ�~m�`Œ�s�C�Lj�8d��a��mZ���p�/O]��ejҴH��`��nFض������T^�����d�98����	����+S:��r8��s�?\�����ڑu��r�H�%�ԮaCV��"��{Y����$x
fU��❥m<��覃�o�=[�^��@14���}�dԵ`�Ύ`tG*{G�ϙ�U���4L��wnN�- �˞���<�Fs7Xб>��nxi��\d��x�^+ky�fV�5I�ޢ�g�^"�_g�����S�f��Z9rOL�g���p���'st��m\se�p`�>Ez8���"n^6{-�3١��BT�&
at�0b�6��;j&��Xd�A��iV�\�m��DzJ�o�;R@Լ���}�m����QH�+w�jqb�O���R/�fV�p�,3����)�U�CBT��o�	F�m*`P�ґ6
��q�<w"�;�{0Us��e�#,�����?u�hn����rmW�A�:Oɶ�Y:g�'�=ʥ��<<�kRӣð:�9�D�9'�2����%~���u.z�:��E��u�C��_��f�G�T��2m<c�j{���XNJ�+�14���R��'�ֵ��hE�,������Ҋ7K�����2r�v���[�!�@C�頞���fQ�5�>���.�:����g�U��d2�0�%��" �`�����
a��E���+��� >��/g$���X옿l�SD��CH���E���j�{�}����h������E~�lj1��L����qE����Ť�E�>�ȣB�{�MÁH���np�P��Bx��=/Q��Ŝ�*��9�j�{j��=�}"	NO5�E��17cCJ�'�X�}�J:�EM��k楪�izx�]�Ok�D8K�7�n-d�d��x�RFQY�����5����d�&΢h�5������F�����J�x�a �u�q����v�������C �;���(X����J�j�jr	J�"ϩ>���J~5J���R��&�QQ����E7/�_���~؏��H�|��4PQ
���[�	�F�uG���,�Ƃ�2qDJ�#�3������W��ป���[���K�X���{�>%%�!v���v�h�Zs�(�\�y�EN�F���v�����Sc�([ǡ$�/]Lҗ��g�G�X�<QVܶ���.<�yl��xQ5�:��7ꄯd=myP�C
vDh^�/�{�
�;ݟ���W�ݓ��O�$ �_�Adt��8逅_��q����] ̊T�����5�-�,_�ضM�n8�����"��ٖ�aZj֎�e�(�F����eKq�,�+��TkX��h�� :��> ��_vVrT��'�=_���vJ�����5�mr[8o�8(z�+S�v$f���ѽ�O�.㎘t+N绉Ba-"�b����]%:����>$���vAr(���z��>�7��Yc�_�zĽZV�����Uٞ��&�oʓt8���r���F�ew�/	K������V6S �l������e���t�)��C��;<���0�<k	�g��V,�#Y#@��u+ � �H u?���/��u�_r��	%16y�J�z�f���g�
��k�	{���Ц(m�ȩ���#;�F¸π�N`^�\�N�	� J*EuM� h���5;F��p<M@�[�J�E�p��L�0cӧ yh��<��ʵ�~���҂�`��!�����x�ʸk:��6T�f:u!���z�Ɣ%��V�V�\�G+p �6�H�f��q���%�*�^�?V��u�[A��/҄��_�d��V3>S���P)�,��}�Yu�TS`��E��\��e@��#�^�W��o�$�ގpn�;���/����U�0��΀�K�g+��By�X��]se�Ǔ�G��Pd��'���7�M�I����`z�L?NzN'�����~Ԋt�`#qL�T���z%��0b���yJ��I�p�f�� 8�D����=}������f�zȘNҹOH�!F�]<����;N��)嫭��/�Jn�3���&u������#ȷ���ۺc�- ����mċ�e� ��б����շ�n����Fd�m>�Aבd~�w�/p�]��8(��[�cN���{Ho�/�|�ikg����bLUs��I�n�(�21�w�aG�/��#���"�QdD},٘P�Y��*;�?�{�U�8_jgi��O�Y���0jaN=�����׼�/'E	�|��2*��̀��:��B��?�k�czo"�o#�n�O�����i3�js�,��D��bP�z�߷���㐩����ဎ��~�'�|1^Bf�V�IVr���v�����SD�f���7�+�-k�"Lt!3h��-qнLd����!��kZS��j:t�DM���0�Cd[<�j�q�ۖ���K*�3}����y���A2쟵Q���1�C� Y���|*�5:Hp�P!��r)7r���S��#ػ{a	�ɍqyL�B<�s�OS�'�5כnS0.\�U���{�d������n�Ss<��a�A1��k�F5�f�B4P�ı��_(��ϳ�8J�v�i��5�V@���m���S@���f	+J[gb�	�7\0����[�����������l���%��*��zt���G�Oa��=PN��8[~�NB5���YQ$�Wi�P�T^;�4 ?Mv�����]�]��Ҝtጋ݀6���tƛɅ>��4�U��0"6V$����6���W�8C�#|fsNU���������?�*<I�{�w�A���.�㠘`޺��l3�1���:��c���O69�.��>�)����{`<�g�1O�S���*Bl�T{����w\#U�vqǊ(	AI��S�q��V����ܸ	���h�}�U0�mM�$(/��,B����e�9 ��(W�ތ>÷ݟ�4#24��b!�E�IR�b*��7�:)/�-,W"��-��L�/�� *䳳5^����S��V�E;f�Ӣr�Ī���CI:�mS�+���_��*'2w�����`QJ]%��'�8
�S������¢��SO�xÇۻ9��97���^�s��X�S�N�m=\.%qS��b����h/��{ d��v���51��cF�*ȇ�
��Pm?8��k_���f�6X�x��L/������<��	�{B??�����l��@Ӂɵ�	X��U�����3!~H�Q]�M|�#�����k��4KtN���1p�N��j�k{�0�?��f#�#G�����U2=>��,�������(jx��8@�b�� g�1����JD�x8C�[���I�;�� �L�l	���z�#^B��_�?�>���}�y^F~��(r�iԝ��Qt��$.�p����T�c�*���fQ��OGc�)�FǇ��-���w�r��n��;��?u2��kY��i�i�X0� ���h�4�é�`-Ź/8�K�M���u���Qh<�F�kP�/w�p^�1�b2HN��*�@�Os�-��P���>�g����[Ƥ@���pfm3q1!v��!_���6�3�M����kmM]8���W�dm���NGo��7
%��94C��ǻMA�P<-=���XY�~���������N�9�����v��*�Ϊ�����D���=���p���{�2�:.�NYYUS0=c#��]ذd�CFI[�rBm�l�pU *P�bV��S6��� �yϮ=��Q�2���ʚ�J~��~�O�r��B����{]z��۲�4�^�����r�$�A@����U�w�����f���Xɇ�JK[����$���t�i��n��--N��y�`*�#jdf��z�*ظdh$~gCfGj�h:�(,ja%��Nju@,���0�^_�:]�6��U�Q���0O��Ѽ|��Uh�\�L�+(���]�-5�sp^�2]�J{��8\!&\�ދ[9�,�w~����8�E���@c���e�!�j1�${��.;���N}��Z2a���1vɉ�%�;��y/mRG��RXo�sQ���#w��Sp�i�wpz.���/�j/ͼ�m@���h�[M��va�����I���GQ��Br��;�=+���]T����K�������.�9�_f�`�p8"�Q7{&-���z���E�7ƈ6JV�I��t(%��	!��.U�F�_ޫ����q�ľ4�[����e
����M�Vm���j��h��,�*.8����G�9O3e��n��<XŬfU���ꁜ5c��RR�h�#Q`Tm����1[8Cqd�����m��`�p�| p!KO�Q�� N>S���ۈ����k*���>�m�l{�Db�@kNV�)�v_��i�'|_�5�y��}�; L�~�u���ʉ��b��
�0��e?��W�K��R05�0���ӫo;I�Z�(	2��I}�B�x�k+K�w�3UGf-��d��>@�{���Y�h�&y$�n��簈A"K2B�Ą2=>L&�<n��}����˧�\*�m�B���#�S��I��M�f���>¶j�0~o~#4Ǒ2�#��+��	�3�0@e�	0�|�����ԶT}�5�%��Ǽ�d]Lu�d�=�(o���%���Z���ݱì���>;���+�
?����>7ѿ4�+f,�E ��1K�𰺀�  TMbU�G�f�΂�7��!ºx�.�����#��-mK��F�S-�^+c�!�/߇��Vy�nA�5���q�w^�~�㘺>�TO�#y��l��،��=�{A����wnᚋ�xWP��f�i��v�$�ؔ'��TQD�nA�� �$�&��!�@��󅳝����o>ʗ�g�%����*��4ғ�p�;s���b��].Fh"��݄����; �*�e�