��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�A�R�|�%�+��}Tʸ	"5lr��~�2�����
�rn��8\���zMxSΪ�a��|2���7+��@zG��5Ynq��-���;�;��S�l�����呮ϭy�&U�}���D3S���BY��c/͵���d�o�f�>�X�.�.<�t3X3'v��=b����Q��HvW��r��P/��̽>�K��YY�ݏ7s��V��F�I���M*m��\� s@�rqӦ�oK�[uĥA4-ʈ��~<��R��qK�DK�4鹱�Z�)����%��-�r��?�Oݠ0�c�0j�C'sޏl�R�mG>��u7��撜!bƶ�EG�@��]%��
� (���Ą_S���sPJ#ȓ�l�ܷFS�JyA����1[���z�c���[E�'`��Ѐ9v�U5�f�?������Ky �)�X$��8�����;��Ձ����_ph�#��.1�~Ό�d�ɯ`mj p��`>��gM_��'�R+�Ƭ�ᗟv�����`�!��a+�'9��m�c����+ש�		�n=����Ϥ�
n#m��hr9����r����(�p��C�� d��}`�W�S���y��+&ɲE��֬�ar��c`RM��F=O\u�tѦ�"x�K��T/�����U�w�.F��Y�?H��5���vخ�'q����/��G�3���BY��˩��tq2�X>NP}�Y1[v�ݟ'��lH5gF��o���?m��i�L��7&����-?Lf��\�e�O�՚1����N���J�o`�x��Wݤ���;��v~ިo*�&�;R4��)�s$|9�{Z>���cĖ��	f��S���K�#,]��t�1`�7�����t;��������<d��c!p�2ݏ��B}kT�&�+Ge:jY��3�7]�BQ�K�isŢÿp_u}��l����GY8�XH%Ħ�D�e$&����8�.�}�TtӮP���f�D�*|�8/�����b-5a�@�X�� %�� �t	lӪ%H<��r���'_�Qb��s#�t��D��@�s��������LT?~IUw�s�r��Ӈ&�m/Fv��]��Y�e|s,��siI�e|-��f�O$��2�'�U�K�Q�&�#�+�e[J�阨:*���7���j�����$�9k��籶x��B�\�S$.��=S;:N�p
�JKH��z��iPt�{��
�uyB�" |�&/��W�6�6(]���I�]��PE��]O�g���*_�����\3����Y�U ��#aؔ� ��}��#N�; �L�:��/����asg� p�%4�8,�/�H�'�:�����p�_�S3���Fs�3'&��d��z��,?�<���7Z)�io��؉�����b�%YV��Ǉx�!J=��:u���	�-�,S�㧒¥N��4xt\�7�@��C��*��{sL���n����������0�C2B-u9�}hdş���3`��v����p�Ӫs���+ P�{���@�� ~�7�m9�'���A�Bk�p�
͆���N��#��?iZf� r�9�
,�g�7f!
6��n/Y��N�8E��nK��B�n�$S^��gz;�mڧZw^+,���|�{��c��D��E[X$j;c
�I�&=�+���� �c�n�O��A��#5�W&*0�A�00�S75�H�������WdMG��f��Ixq�l��:!��`/�`�.b���Z��P�߶���Y�
!�m���}Ĉ�e��Ҙ]	W��*m;����\j�?�$�1^����^a��6��$/�Ӗ��{Wס�o�*X�b�����㳄<�gj]��%�MQn�!���[uR,G]�$r��R�V�L��E��0��4M����"t�;����W�Z�\�`���µ�A8���Ī8Z}�)+)"�S�� A�eN�7��bH^	ޛ��D[X�=�@�Y�V�(���Lܟ���tO��\A���k���;�{��+�A�gۮ �sK_��d�Ɍ�� ��2��U�W��3Д6�C2��_aj�D���`���P��_g.��#��R��h,h�+��0l#^Tٹ�% ,I�ϒ>_�^��Q�ƺxZ�Å��	�t�Ρ^`go��zBCf�k���ݜ_U�$�E?�E[xƗFd҃���ԥ/�%�mH�;v	Kz�$�c�l��!S���9�_���f�WX���B�1d���\�y
9�5�����F ���x�<Ҩ|���RԘG6w�Bi���i��g.cO�I���PD����#Y#�n%�c�
�τ�D��-�;����_0����$$^�:<�,�G���L�����0;l�p�&��r�b���1�%o�Zf$!P����dߒ����~'sy��-]a�<����\�o��[�;�TE��e�tA����h�nM�	8�;�b+WݒP�iFb����)J���đ[g������y�H�pք�G�MI���+�sB4����t�o�d�'U+�WZ�a0"V0�;{Ԯ����v�M��'�Xې��?خ�]��B=�M_�gG��.	oy�s| .W�]�1��M�Q
 �(~3��Y�x���e�Z�S�����'91u��Pn��b��v#�v�U�RƑ�뉰�'�����ۉ�����Nn��0�i$�Ń�H� H��
f���`���_����;�����Iy���9'���}Ye���T(����
{"}L1f8��+.f
�GfX�|��Y��MK����z�ݻ��_0lK�o���N�9A^ږ��s
���c����A���EZ����Xل�3���%&� ,�^�P�#�A�r��w�A��W;��9hX��Q6�0#a$��+ܾ+���S��Ňm�d��wo:��Q���ļ�XmIy�3v	�gmq�(=}���箵�4����]�i�o�u#4��F�cO�aC?U��B1�� ����N�2YG-�|S�'Pz��+�ͣڑXV'� ^vQ$>S�̱���د�ǧoֶ[|�!]���
T �<$m�����9$����\�xc�e���ۣ��&]\�U8H��lD�����CŌv�`>��v�#�XX�	9Z�3�P��9�J��dTu��ѐɺ�	r
ûTX\�����V�w���$��f���4���Oэ ���3n�oNx���y��y�QzÎ����C��jz;���D��TU���R�L��=C�?�0Gq���ʩ0	5:�w��Ŏ�k&��>/#
��k��H�ê�AK[�N�Q�~v^B��ď5�+��'�9����k��K�.��;���ů	�jY�R"�s6��x[N������k0�{{���q��i�k
r��A�{�ག��ySU�*q�����W:�e�9=�Hjt��Dk��a	oB��
�f��7�6|�Z�f�%J��뾴Ԫ�����J!���g.���a?aҍ<[5�1%������7���y,��V�� -�!/�#�j���: �u��1���C5�Rm�Kz�����`�2��<�:�YL���'++��_�T��_��^!hk$2A):N<�=���y[Z���;���#��K?�)>�X3j�ʯΏx�&��Mf,�g�^|.��W���.��Y�Yd�pC����w���k�o,*���-p��8�)H�f�kR!�L�f?���
�R���<��i�v�xpZjz�sh���X��oW^eh�U���B^|W1�4�D?�c���H�mM�Y���jκq�e'�������$n#�$|`R�z���m�#��K�������41KX
��:�`�x�/���xHL��ɏ|{��׋�;��?�7� �[�B`�g���Tj<�A�#<D��GP�VNU|v���Csb���WP�`�	e�\T\���%���6���43�w�PQ���U�>�nAx<U��+(y����OʙR+�A�ޕ�@H8o�i܇,�8�, �����9*�n��`���I&��a���	�����6���,��|�@Y�1a��+�����L�>�2����a�;�Xf��[B%^�NE�)"ໃ��\T���Y�?�Z�����u6ڹd
�<���<k������6��\���z6��S,S�AQ��[�(5���?
�bШ�!��Lޮ��m5S�4dQ�f�b�Z҃ߵ��&�b��-�8�u�� ��?/��%��ꐇ� �Zq%rb�u}k+�OH�2���!i\���:��ĹKr%�Ҏ+ܻJ��Q���h��{|D)�W���M5��)���^sf��+d�&A��O����;���O5ǫ��T]{i��-w	dC�M��Z���(�R�L�Q���׸�W��.��:@.Mi�d �8��+s�H��I̢���K�'@�ƶD��i��Hr�Z�����`�`_�!�'�6t|&���}�ʆÄȪ�U�H�ƀ�Bn���0�G1H����Ug��ܮ����T6;�{��g��Wā��4z��<�P]cB̦X�a!E��T�� ��]�TI�ɕb��$��<n(A7�b�j��q�����C�R��=�}��
�B����mnIس��=
��U*S����i������GU��[d�9ΏK�4��a��x��סd��~��)Q�2[�Q8x0��zq�<�IY�i.r��ǧ����4&�;5-.���F�o�b��Հ�_�-̇qV	H��w�`V��s�y��1����t
�5)��v��[�0��nN`��Va��uG/!��p��͡�jM��3
	g	1c����%z 8/m�g�/�&nZ+�b:�3���>SZ�����1ǃ?�'1>rv.=862��8�&��7 ��#�-�� �����m�fէ��i�z_d�5)�yΙ��6(�C�:B�;w�G�jY�(�q�-A!�'%tҩ��:WP+��'����R�5��%���}�'D�>ƀ����u��z��bM��ZW!�bI0{�����䖀Z% SCu0=%B�i
�Uu�_p��� @>�p{�(nm.](k�{���r6}G�f�'ث��H�&A�{wj�ܢlz�%9V�_�g�� $��PܕKT�ڽ�kF���,�[=���ʔV����f����!��o@����8�\���lHӇ/�ܟ��E�>h�r���/�ۍ�L|��Y�
���#
��$=�τ��}���o����Z�D��sG� ���i��O�$d۫4��۴sx4Ӊ*S� ��ҍV���4�DŚ\� �-�ݚ�(�p�n
ce��Jz昼�U��
x�"�;�c��%��x���?s�cI���F�Œ�`�����DŇC����������f��ˉ�� ��LX�}���RE2'����Z�\r��6��[��ݍWUA?5��9}\f�V��hA4bӅɣ��o���g��3!����ޓ>*�J�;\�,mp[��;*u�#N[���ZO�Z��<X�R85a����6oP�B��ߢWyْ��d�^� P���2^g���� R�$����W���ht��~���YB@����ӯ=�8�2�b�ܪdÀ&�ˉ��6��h�C4~>U9��~T���Ԏ}�x��$Y62�n��L=ߥH;�XǬu������x0���qY���3Ab�@���heȰׂ�絾�O��L����V�� �`�\�\�S���|�����rѾ졿l���27Y[���cB�^>�������|�b��h�9^h\�6Oj�*�6���`$r����A�t(վ�t���f2��f,��V��ϔ|㭝:�DB����9�_��ؑ����2DU}ךA�o:�J5Pn�	hΤ%=��ӧ�췤�8|����BU��f�+���	��q�32#M�w&U�r��G�oY�8�f3��g����!_��"i猲z�UH��E��F�52o��C,���)�~��Ou?�"�>g�O}	W� /��ҝs!jhBXt(eR�|^?�M�Ã��C$z�"?G�q���̹���������L0���5o���pyq)�0��e�P�㞤�G��&�!���k��6����zSO��1�]m��=%���Ĳ�ok���5�����"�BgG�h;aKa�r-1���(C�Q�w���X́�k�c�p�O�aq�M�����&���z�%m村�9���\\.$��ʺ�0�ntx���6�p�Π o�X�ni�y|��gc]D�t��a�s��j��Hu��0AE覦s	iʒ� �+�	�S��
|��o���,���DȖ��}�Ќ!�ߧ�V"��d�	��c�s2�)y�]KTU�� <�d��E��@��fQ�l�=��2ܹ��$�m�U��K��x��	������}dM�6��s������ʐ�����0�օ��- ��+g6K!%���d���p�����% ��J�k�����(�����N[I[����*�tF+qO�D�g_Z X�jC��}H1��ԏ�Rb��_XJ��.�!����7��]��V�?�Ԣw��ln��]�g�X�t�����1��X꺑<8��0���/�4�n�fY�B�ђ�%�"��ܫ�;�S�dh�pe��bo:�"�O�������(�bُ�wȡ��\�	�~<�갺���=�	j�F��⢯{��$a#o ݻ�(]#�'�a�K����;����6���`�٨2(�� lM]eA��yq%uUh�X�f�"v�Ny�M�3A���| J+��~�f��{�Q�X�`�>Ɍ��l��W�uؤ���M�9
��,��'�za��5u���]VV��o0�����&\y��p�/*Kc�	9���[u~�9�o���{^�"���7 L/C�����������q��èo�lΘ�ø���n��ޑ���PFK;�Es��1��M�Ja�79�6O��2�b�g4S�Z����l�;�����y�8������:Q��ىSt!��/��^E�� ���"HaH��N����>/��YћZ���l
@pX����ɭ�[��",
rDd"j�F��	�Bt���[C��7�7N��`Ƽ>��\$w�J4��g��y��$)��֕�}:]���_f|���Kr��v���up������7�V+�\��a���	�%��7C���#`ѡ
h���|�J�A�G}�^��� 1���WXO꼨:����\��J��upy�ل�L3��{�^�}ݳ��Z��>��Nz���9#�? �ȏ��voI�6���Y
�ԍ�q�F3Yך;x��|�"�*F�aٵ�mH�n����lI��e�`�] ��y�&̰u1�:���s%ڦ�-#� j��h�"�#u��l*��� �T츩7�x;>�b�A��y<��r/kK%4��'�Nܽ��Ĳ��F�b[��P<�f�Z&xl����9;�j�:R��j�o[����jҍ먟�!͘�DS�%l����Ɛ�5���U�7��\_��5�K�_�5^	�$�'A&'���KXK��:;h���&m���E��KD�!�$Q��J���6[�SI��O�&�Ӊ�������W[����y���m�}�{$\>�$�:\�NS
.��x���Q[�@���?ɛ�Q b�]d�@������ΙT��.Ҥ)t�͊��0�Ǧޣ��z��h�Axk3J�u�X�+�Q�Q����`y��%��Ʊ�:o�w�t�������~���F���� -���)%��� �e��k����'U�ET�æ���=��.�/���mW d��O��A,�����⑧�kF�)l���MM�9���k���C2���$,���j���$���fNI$��kB����ae���P��m�z��i�����>��0"����/�y"���p���+����uQ+X���?�Z�DW�:�xa[�}[U}N��k��
��1x}kg抈���TLvx2s�B���T���G���3����q闗8��0=�D���h�3<�g�`��H΍�Ƭ�}�o
<������,3���?���B������0��*�� �!e���s�ʨ��Б��1W�g6����2�!�Nz�u��3��-u�<�m 7�&�9#����Q����w]y��PJqF���*h�4�|c�?B��pI�)L;����ë� ȇ18���Y��U�]���n�)�6�5�[���K��S�i��i ���3](�[��]�x��@�R�8`�\�O.�Z�	-��P�ϭ5~d|�¶fE���d���Z<�(QkF'8���i�[(�9����~�Ӭ6z��h��ɉ���R��*�Ud���@����_�+O
���I��"=�yh��e9�ɴ�Ła�!t~�u�U
��{�ìƜ�>dj��6�Q�6zz�����������VV����r���L5Q����H+�]UD�a�	��T@i�����~Ď��߼|i�A��z���� JŐc��!��jL�XK�'�4Xr�t�R�)�E�z�"l�$هPd���$`��i$���-���,6�'��2~a���O=5��;-bc�Ȋļ!ԓ�T��1'<+��B���\s�S��z^z�"�ž�L�p�O	E���\�TB�(���O�[>՞���f�i�i�T_���O�ޡ�QsU�4�6��p��i]g�Ӳ%v�Z{�H�< �!�?��c�@O�8��UF��Rt)��mi��f�@N.�kA�ʸO<K�Y��&ж���~L�,ܠP�<��^��ط9e��"�%��m*�*��A����L<~f�&Ȟ��#_?'�R�9��r���S��N�E�+d�Y�Z��C��n��^���>�R�g9��R�u⺃��R�-u�2�h�cXE��*ʸjS�����2'� �,;��J���0PKV�k���%ۗ�jbp�a���?ќE�2T���S�!�"���3]ĺbU�V(�\z�?��"~��6�����oy��+Q��)�伛�
��E'�Yh�]�M��A	�B�.�z1�z,-�X�Ê������Ճd7{�wwF�L��fV��sx=�^�lfD�׽G@;(��"p�ogF�J�Լg�<�t`��>w�2<t$kf��h�#dк�,�B��뒙Q�E�3�$Z�������7b��Q���59�@~s��w�SVI�Yo��-�+��p��j�%:����[�o�r��::W�M�|��MۊnP����C�L��	���Խ�����;t;)���*��HQ���
#������p�P#���"���,�����\�ծ�x��g�H�d8�B97)�*L(}��eތ�2A^�V�N����x�P�]bSWib�"No��5��衜�	M	��h����5�QЖ�'G�Jf%�`âr��	D�D4�i���৹#�U��<��`ˋU+��gI�╝�=���f֢�`�`r!e���� @c��s.~����j���Ne��t:=l����SxT�F�uw�|�H���ջ��?�&Ʌ�C�	ӯ?�v��0���\�G�}�-f����y��9������j��Ua�0�NRRw��ab�c���VJ���l/a���^z��}�`/Y�j%�>?$0��2��)?���p(�������;J�I���#o� �_�A�ȾF`aB��߱>	5�=�r��Ҙ���n��b���ZiH�ᗖ&�	��1����EH��]�w�
�X��j�U��(*��N�7�`���qc�5O��>�̯L(Sz�,�	<y��x���� rֲ�;(+3�Ii���:"�������F��"Z+Ĕ�9�e^:tNH1���?b��٤�����h9��6|�65]��OM�K����o�?<��j�Ŀ��hQ�Ԑ�]�`c���4�_�����9ͫ-�k���������|����Ү?�=pE
��H�lxW�9��Ɨi�,e�Qz���Ȫ�'F�*���G.�4C�(�o�B�_B�f�*gu��?��>��DERG��1� �`x�O���[���V��D�W9�l�f�C�� L(�s�rts�-�-��>�*���O8�QT�0V�ȫ�Ԛ�`ϙ���k���˧+����)�7� �XY�w�$�� A,ZT%��QPM'��������/Q����V��Uk�I��������Nv��AO���$LqX�S1���4�n�D}����9�T-�p7JuAT	�i��^&�vk�*�;��m�I&��:��ww����ނ_!8B ���׽5�]�|
�M��"��C=ښ���"���\�ָ"J+�0���@I�}��7�PͶG&��WM��������b�F�4��;�U�I��e��G;h����_K8e%����J;ad��X.������x�Sj X�ܲ��_�-��fN߻�.q���wE��A�z���r��.Su�����Hۑ�(�<�ZY���U�?�l�ظ([Jl�t�QK���L5���_����P��R����q)�a5�'G��%������5kG��n��8уg�$Ԅ��@0Y��s�1�|��&�D)H6���A�^~V�j�v�8/�w���:�!�A���-a�i9)* A����4`�y��L�e A6����'jc�����&�|��r�a���i[vjE�8Г����Mf�=�4�g��^�!E�+��1	O�W�NR�,>F��zȤ�-X�%�v;��6 @��(���.��\����w� d�U8���zJ\�x�,G%+݂�cD��r��LK_ag��:�%�4�ܡ6g������p㧤Fv�]��
32Z����|>�U҅�{�ƼIT�w,%�wzP�3,������kl�aY��ؤgS�v��"��"�vԃ/]�,�5��U�����^d�'�Τ���@�"7N=�#���A*X�`�j�-/U6��W����8�%LK՘g��]in�|�D	�煻��G�NMqb�I޴���G��5�2�Ԛޗ�o:ow؎j�Q���D����W\D�A>d�IY���Q�.ܿ�G��M��5�E�����bM'U`c���̨ߦuP�5�<E�v9s���&���IY����t���x[��G߈�wYQ�����w�x����/w�Ī�-^���*�"1������
�]=���F<�VI\q0�A��g��+L�B�7��~���o��ۡ7�p��l�<�ˎ$�|&⹪��@z�-C��hō����zE�>��4�W��Z�&��إ�\�'i���X@� �7p�;����3<�V�h��D��/���m��?C�����6n�:�*JH�H韺��L�9&Ӥ�H�u�̨+-�Y4�%�_|���]��<U��:����B,ղH����וr#	��ݎ��]|A�F��,���WQ����� 1J�Lh�h�5�x�&7�f�]^E�++wW��<�!��%��)��w̅$�29\��֤�V(C���Sa�N�9D�����Ԑ����d�H���B͞l�b>8��z�8|+��z�ܡ�� �*]�I� N���A�e���S�8&ײ&�B�>��'��R%M˖��a�/�ӳN�A��x��˳�S�ᙗ�L�;>R���]L�I�+�gn,�Х��5��sxZaÄg}G�TC_���F�p���FC���'�+�8�)��c8q�?�f�l�#����n��+. ��
�>�&HM-Z2���#dA$�K�}W	�/ХnƔ֒b����K������?}y1+��	��[���I�&0�����r+4��p9�����g�'��^AOw��it	�N�>�Y�㎥�q!L��D൙݆zg�Y�gj�P�}�`�jr�p$Ed7g�ec������S4 �{5�x����u��%:�� e���&\���6�x־i5�:k����Ϩ�y������j �67b��Ш�b��&P�uNI��"Ք�o>'�e��o۝�ЎubU��ƾ3��A#�TnQ�����J��Py^kh�j(�N�Tu��%]�4aN��V�n��2v��J���r��nev�2q �4Q�p��B�w�֫��*����i1�`g`�F�� b� ��-9XTM�?><��]�᫋X��2[��2��F�3�Xjz)���n�2���U����~d�;�4�ۯKƭ�QX��Ws���>�q�d~"�����2��=Ńތi8�)�ȓxz�����%���e�9����Ŵ�/���y��T�M/�����Rˁ�/�*�M�=�,i�+�
�9�P����O�`l��>,����>��������E߯~��Z$Tt�����,ig�o�w��>2,���/�V��+8T[L��)P1F�+��e3�:m��_D'!�g�v����k�E��y��C�ѡ��	�Cp?k�%�Uԣ8���v9���G�?�_;D�z5A���aT��C�B������3��}�W������GN���\��w#q-@���!�ϣ_���ߟ�>�P ��Ѻ��FԂw��,�c*���7����[6��o����9�{�����#B�:T8/���K	��+��f@td�&����[û�?b�c5�A>���U� @�I5��R��g5��h="�v4��yd-U����J�*�`#g`e��sED'��&����?#*4��x�ҩ�od���\�AvM�,���YEٮŧ�`�hn��C(1ߤS%���J�CU2�,���`L:E:7\�������'�x��@7o���*�@.�g�D���YA&	��TT�5����F������X�F<26�0�gр�J���.�m��?�PSK�mw�� ��h9��֫���mD���>�Z���EU-�y�;m���nv��&�e���l�U#���y[��c�<�6�?��Z�%����멐
$�C���\tݠ���z��^ǋ�4 ��Y�p<�g�Xa���.*�|��%A\�!Z$<��+�����޻�s��@+Uf�0!7fE���I�$M����h�Iƛ��Ó��<p�#{�xR��\Q��w&�ɢD)���HD,��7F��E�$s[�`�Y�f�x��.�G��&�Ւ�JyB$n�s� #6�$�@�_w��#���:�#��M]->��/A���J/�n0��5����Ƴ4�Nm�)�6`��`�:�J�W�t��Mr���;���F��j�f�SH�=w8%�nb�����G�����e���^���QP�p�դ�Sk�B%�y�ր���i�cm��UӠm�O8�w���h��i0�+�m�L�в.j7^����0�t=Z����,��?� L	�	���٠H��n9����i��]����5:��M�b�[=�9c�,��Ksˌ���I��J=���4�nd(�M�3�Q8ϔ����.�2'K���ۍ��B��֨��`h̯���JC�ф�b:�.y�:�&L��Q�
��.r�A���=�\ۘt��@λB�1�=���vE����&�� W���:<Qtl�o�1"��y� Vm���N?KN�z$ڱK#������XJo�w����V��~ ��u�@�&]R�C�m$ Ќ&i��(p���2��k)��n5��ւm:���$mGlSKѺ�	����f�/���:�c,�E��a�Bd^چc��p��*����w6���P����J⿳�,�|����2����ܽ�/[|"�ҩz�?N�����@\�/�R�+�o�#��Sxe�������K4-�蟐��r�FG� �n����������Tۤo�<�\+�
��z�yÆzg�$�����qG�.C����f-�&�F����h�:g	���ONb'Z��!Mek���fM���<2
c(�n�l&ɶ��fɣ�h$�/9�V�n�m�7ٷ5x��8wMxօ[sWxC�Sh=s�����r/��NY�X��Brv��_���%��h���J�m�.�G��3px�k��-�Ȩ#[gl^��sA`z��;p%,�	Ţ[����0]�<�y���9�_}9钆�����`%\`g��?���)�h>읣2�pb���ϩ�Kl�Ag�2	�1�//"w����J�{?@�H�c�y��ʤ�K�اW�5<�
���%��n9���Pݬ�RQ&�6�Ǘg��B1�>�Fs�W6���m}����N_$����F����j7ϲ7�{��	����R�ПupB�ri��tU�2��}H>�ti'>=FG������	����
�!ۥ�_:'0�pъݘY�duYHӋ8ۀ&�A\�Ѩ`E�
Gk�f?���,L�&�����1VH��K���)�VƢ�g����'���u���|�0Ř��SڟI�D��gQ��ҳ�K_��q]��ݘ��P]�w_���X����gO�pw�]��> ���~B)�>�1�4���z�W���Ǡ���������od��Z��;��}��Cm�d�o��+"�8u�m����ʍ�!g�-so(�$&��=��A�r�����Ҁŗ���gJ�Mi^��"�.��/��d��1��Geо+Q�s`xtZ��T^�q˔�43��T*'�¸D�Y0�MpR�ȡ�,_)�]M"�$�)O��6��3o�������wW�Z�K�
�A�>��)�͚�*�U�Gx�QQ�KΥLA{e�m�p��E" ����ܙ�{$�Y~]|����f�ϭ�R=��o{xN Ygr>&~K:�40���|�d0%�,��c�F4+$�R`*�����Ov�V�>{0�q�^�#b��:O#��0���`N�(Ǭ�:�Do?i6~��w��G�ީ��Hz@�C�R�Q�d�a�|Uy�R�Z�;o|<�,��)�Ĥ�Vk�>wU�W�U��l���2\��]�;�&���)��p���BK%}՞~j["��
F�����^������s���᠞�h�����:��*ov�z@����ݞDF]��ת���0t-}��q�RW�2����|�	�|M��h(u�$��ǥ5��mNs"�(Z�&��nv��O	��$��}X���Ք�����I��T��M�d?A�W���q?�K���~O���}�{P]�Z�{n)5�#���C�ިBy�U�lOk��F��V����;�&އ��=�{�R�+ {51�1C�������K�~��r��h�v <ٖG�*�MJ_ҁ�qRI�_��qP$h�)r3�Y�'�K���#���R_n��T�eqB>Ee!��v�\v�iH���9Q�&�iZ%�����؋zN��#k�i��M�����?T��q@��� ��⧙>�|�3?D���������b^Q����V�q�'U*̢>u�.b���<�
j;@/�$��PW��8-�uU�('@(��᫽��~?��xz����q/z�`���0P�X>ܮBP�
�SN|o�S�\��B�8�:7Ze���O����{9�U��\���]X3�U'��៰4�+�|�����!�E9s�'���N7�H=zF�Rq����o�����t�Nѐ~����j�U�����n�GVi�_�*Y�|���~�t$��i��{���0M	�-_�ٱC��- ��ݮ+I�LS�~2���a�>��"d\J	�A8�Z�?ދ>�:����g�5͙����K_�<@�i����9��]W\�t�7o�����w�12�K�)�	��Sy���P��b�s�>B�������O?�n+ϋ�U�7�ZSBN ��OByN�Tu�z��6�%3f�L;M�O5�+���i��@t9���c�/���Ӭ�O�.k��v;6M@�h�[eJ����T6�f}C�o4,Ī!G��*��>���6�
��Դͨ�ȹ�p�h���K��#ѧ��;{�
��1�>�J)��0U7��	ċ`�O��� ��U�wkCv���9a��9H�8Aa�5Tu�kJߊp�%L̊����]�8�\���%cMsJI��u^@�{�����"�f��#�XR����_�7Y�
�_���÷j����,����м4`�Y���P|UK(}[֠�&��m�2��J`z8��3��P	���P�%c	4��Nz�^��Ƃ�E�
�Bsf�����yh���=Ɓ��.F�aj*eLU��i]���yW�qx��������'�e�p��+gp�)���oD�Q�-�ל�3>4xʌ
6�͹���=��WS��� !�r�S9�\�D5��:��Tf<��ߜ\��Y�Z	�$
�ڼ�_�:�DAٞc!�hG�&2�jn�8Š{,N=�ҝ��p_y�f�sAi%�[e=�����ڰJ���/584~c�^r���;���Fz.��tQ���]b>i>C8"�[*�|�Z�'5���!X����tzn�L�%(��B1q���靳�;#�V��J=S�>���WA���n.���ny0q8�t1@��-�|)�7�O��H�.��e�1C)Ou�X�ܨ=-mY���)G���D�5���w�hc�1}-[Ɍ;����;��y�_�J��W���_3��2�Æ�r��n�K�Pv}nv�/l���wZxmM�ʠ$�wy�듯�DL���� ��`�A���Ж)�z���mb2�za�Mbl�ED��.�2.hD��L�i�%zEfa*��$���]�9/���v3zG ]VY@�����M���i���2�-H�ꯔ�D�6UG�ݯ�e�,�4h��&e�TΝ�O�i]��U�؜����1r*ZƎ;f1b�1� �~���_[������<KK��}��c׬M��on�_6r� ߲ wB^��� ��$PM��f���$`ıK"z������#��||���px������2-�_�G;�N��)��6�%w�4u� �� �^el��ތU?"���6]zDFQ �����4�

�3 K���/�gFs�����[��mdf1ԪeLF�>�oP��A����xmS���h��F�������	�7֊ �����R��;�G�������A�s�;,��l��J���GTT�U��DƎ�䄈���wģ��_�p\Iܮ�4�� ^N��ś��>�id�E>n*���F
�X Ne�p�vK�m�Qa�`�|�@�SKw��h9���^ʘ�9R�O��'��@�B�yT{���iւ�?�+�1�r�- ;�c~[�@�H_Ze��mF��w���U��Z�:q����ׇg�WTξ4`&d`����: af���O��ma��S��#�<��8��{W�)Ed�ڄ?�0�1�*�d`ݏ7��:4C��~?��?�]?y���%��@Rx*_�����8˪c ���9���؝�a����Wg� �5��P�>��d��k���U�гd>_���x�[�K !�6csK](��М��1��FxM��@:���O��E��p�� � itB�k^�)N�/|6j��ÐEe`f����F�.��Ӏ$�_�b����P��L��!��  B/f~BR�k`4u1ej�J���~����?C���!2����<���qt���!�C#� ��掃����!��X8&��Y7u1ÿD�<@��Z���Ti\:���<pK��<W+��M�d���
�8~�Sު�Y�Y�����!�O̷��eXz���9�o'S]��q���J��s�ɢ,�ӕ�L����z�j�d�fp�)�{�2�� ,��m7Қ��i@s6��Q4'�Ǒ3*k��1Cb~5� W����A�l�tE����C
6x�g���X'o��݊�`|%��!��	���6a�H���=k��G����
� ���jˁg��TI/�Pj։��y�ϤbD�va��p�g&nT�}�Y,t��S����m���c����36��<��z����r��N�LP�Զs�" ���1H��X�9R��:8Ҡ=%��Fr��k{��I�q�����)F%�=��.��&u�җ�D��S�٪!�+��A4���y��������e�C
��^�!s����:�S�v����S�,������^+ ��z|^̹Ae�_ɛ��TD�n��Xо��=��m���V��?f��I�.#�`{�������XEˉL�4�C�`W�o��
�2B޶��dp.݅6�P�(F�&9�	O!�9��+h�["�����t:�&tw��Y�z^�������*�.i^���y �dn�&���k �zM�=��*�����JU�c�i��H�<���������yI!��ŽA�e�S ������΅q����KD�Vq�u#I���Z��ĘMH}��4��2W�P���_ &.�b<��z���.NC��s	
�pı���dV�y�E0�,��������M�64���P�Q���⮋?m��Q[]�J�Ҡh��%���P��s&�SCy��C��U����ȗ�\mb���1�\��S��!�8������G1��d�O�'��w�[�:&s\����r��1� :e~j���*��
F��� ���+�9�×�;�R�Ai(P�*p�7f��12ZW��k��답ZOp$	���(��y�&=M`���I��ش�"`Ӌ�(+g��I|~��TMx3\���&o\7�{Z���mh7�1�/��4O=�O`���NBB>;�5��Z44	B^=oQW�y��/[㕙�0ё�Hf��x���?���mՆ�{�����Te�4�+�Iv;���S!��9	//��](M���[D�ʈ~T����f[ng��~�a.�Veҵq�ΈZ�w�_��VsiC)q��W#��d�sTP�����5�����;���?)O��K�v�p��'���󨷵����r��>�����4pyȺn��S#���2�LY񨏌�7�t�ӻe�ƾ�����m���K��sq0�F�ݥ6���C��_�A���B�����[�&����C�堂ck�����k��1�
N�x�v.lA���?v���p.�b�7����]���6 l���-|ۍAH�-������/ߎL�'\+�G�ً�
w�y\\��Kc�������Gl��u��� �?����h�	�5�I�������<�[R0�^�d�*%<2��8�8����`�q�2v��������%L�ˑ��i����
�j����~A�`z?.Ց��""AI����]?�w���1}w�P7���:`$�@�,F	i���q�C�������p�lC�r��"R���ߔ�3�V����>e��I��W�.o��!U�>�q�������m6~��������M�%���O;�^�_K�0�$����p@�t��G���ΎH���>;0"q�k��^���]�Q�a�=�����/�b� ;�>fc������Ԅ�{kW�X92��q� �[1C�M?�S�|��r�|0 �0�� =���\v��������- ��>�AOr���h���YU�L������Y$?j��Y�;���;��S%-b���!j���9�⽸b��C;��8�I"D$[AsK&�{�戂˼���G�iA_51q�)Uj]u3��pa��C�P�(�,�P��0u71{P�HN|��V\��Q�a�b��������S\Ս�|�F�O׺5c6J���חʵ�q�v#!n������H��� �� V��3�d��:���8�b����$��SeװĞ����E$��������ǚ�g�ՠ6���ۏ9p{MaJp��r�ҁ�g��G��q5^�+�2����J/ٔ���h�rA4LY�8��Ѵ�m���4���>�@�3(��)��������o\~�=4@���]�3`U���}��	˖\���7y��EW�:G���83;q�`��>����^^T�ԭY	d/�Z�b5�i�L_��a#�	�x¼m�ԛ��3�i���P��TN�'�B���ՠ�'�X9
e�"��E�wF&��E�H�9G!�}������y��%�>�}3��<d~%4�7`��Y04���8�PNH��r5�G��7���]�<��X ��-/�咎�@��;������o9
"���rH�3ځ?x[W�^���ߪ�c�]�l�J��)���mR}'}��A v@����NB�<jk{��~����o�Ƿyp� ���A�a4��TT���;n 
����&f�X�}{雁c�H6�����D�a.���`�(t�5쵿�G��-�JS�\��^��R���v�_N�P�7��O|
'|���wYŀ�j�J�*��+��uCe�����1�W�q�2*���Jy�0�0�䏛d4����%y�m����,���i��g��{N7�4Jܞ�uFIӓ�c~����E ���F�������P�7t�]�b,mN ԁ���M2��?(	l������5���1�g���1j�1���|M|~�Z��DQ����i��4�xN�JA�a{��3�AD]�Atp/t9ˊ�7Fce��u�Y�?x��_i
�Cz�����S��˳�4dq�d�X�8��e%F8��R��1��ҕlC<T�����ZC�w���m`rn�QJY����֒S�|Q�f:�~$-矜�'t�]h@���²��#���[h�������7��7���g׺����5��BjW L��^5D.:{��^�d1gIu�c�_�`r��,����*���(��{��G��N�"Ą٬R���DU���S��H��;t��0'%<"����h���{ �RB�ձ�s�c*�O^��]�`6��?�SI%.��`��1}�[���Z�u���ߎ�P6�� ���rS>7�P�\�����KB3��FQ�X��O��$oT�)�ŸJ��(1Ҡ��&��vb���R�/�+qOI���j�B�m���oЮy}mX����H�t΢TlgR��1;t�yi�퇣�2�2#B���Mv���\�T����b>�%
F�V��.a31(�̐�_�+�s	JU�C��k��d��U����<�լ�.|�|�(��B���k묤��3�4������o�H�+C\J���>k�|3��L�_��zl�$l��Y���昣��2���r��.���ڶC�'�#�c���F�u"��ٸ��+�S�D�=�$��݇ªhE?�(���IJ�@E2a�S���\6����~Olb���¶�L�,|�؁�	F�T���#����5��|Q�h?W)���yK	n�!�lf`ZЈ�9�=bp�n�e	�f[�+�1p��^�#-_�^��!_�s��?̙��q�D��k���d[�i��i_+z���%���{X{��얊W�=Y8l.ޡ���խ{׮ada]1�]
�����(��Mm� �������ƉYWL]V	�2�jd}��%�7l���I��#7���;[z*��Z-E���@wѯe�l,�T^�#/�^o�d�a�G�]S_''������=٫
�]��qu�n��
��ڲ8�Z0�R���^i�b��Ivo������K�R���1��ʟ��Q8��r~�w!W��B�"�l`�����33Am�Z�Yx�{t�$��GcL_*!|������ln�ٜ]�8 ��U��# �D�k��io�W��U��\�.�Er�4>5ˇ���B���������,�eU|�1�+%e�@i��l��XQ����㚖�t��vmv�u���̀����4R;$!9����r�!ҽ����r{�
��y���ךB���\���q3����b��?������[ݖ�i�gQ��_8�����j�m�N����_��Lɹ�F�e��6Ғ����m�up�$��!߯���L������ʖ¤'�o�[kΣ�
��X���B5o��#��;�5�P����M�2o���k@�𷠹��얖��f)��oTj�^WHQB8�
\�4�Z�-_���q��.����m'^޾�%N0ovb�ppWg[�q1�5H?p=ͨ�U-k��_?q@�$P����8�򋳾�����O�A�PlG�fI^���Y-P~+�ީƗ@.��uJ�z�Q�����H:�f2�fZ�%t,�!��I�*��8��3}��,]�[#(~9ԃ�%�o����[�nVh�q�?Бov[NU�-��0�	
��+���tD91�E��U���hfY�r��c�Ӱ�W)�S ���P;�~+=��yS�Bs<�!MK2lP>kT�cR~)�����Е���n&!c� �ȔS�i��A�e�&�ދ#��`��'+���-}S`����0'��>��H�C�MY'�$�}
��I�nT���RE�b"�"D���?վ^Ԛ]��~��E��|�������۹V�_\l/[]_ !`ݠ�E^|/�=�_,M�Y�d��H�'�`��X�ATY�/��@[��AO�}�K�|� ��,+-�)6sZp̃('k�9�(�l\)
�����1�NT�*Qpf�;!��$�0HӉb�^��[Ջ���+#Wd��H�e"��=Km��b��n0ۓ�ȁ�c�,9m�J_κ̧SR�ª)����)�/�/�����_��(K��C�p����{?a�|T����O���	&�̃^��:ӱ�+�e_�9w�2$�Ryl�E�_�ļ�D9�Ʋ���A.CH����]�c= ��|�;�&/
1FCu=)0�J'����x�޸�m�i���ep(��c�M����5�nX�U�;��jq ��)>}�N�2��Q��� �S��k����Շ�rρ��p�XZ)c!��$��� ��G_����� ~g}�œ!�.���4��*��f��]@O�V�`VR�)�9$��R��W��Ѯ敝4�7j|Y����ՆB�X�φ�p�o�I ���eWR������L7D1���~wu��2Z��6����%�~I=�a�3�y���,��r*���_��K!�%�_�`���Q�ߒ�h�N�6���5d����	��A�.y���q���VBĚ&Bw����w\�����Y�P���(�>���#�>����^b8C,m�0"��q1���"�2�%���1������Fek����D��@�Pc�MnC̬�,�r�j��.�=m�1)N��E���9jM��]H/"z�ȖHج�1��Ys~V�����?�hOm�*�`�w���߃�.D����Y��f�c����#�pQ�O��uQ�т�[|2&n2t'6�8�(|�!���U�u�/��4�����d�|�G��L>F����E��_>���g�>kR�T�e�����hf���Y��S=��i�S����.+���$J�}�I�
��vk��8�'��~��[in���:�y�6�VL!iA�`�0,󭤎�;����m��,����	ՋM �����)��<�ͬ���iK��Z�Q�}��1��$�����Z4�$8��N$��!��[�ɈE��(�ǹ�+��"�}<�0��u�f�G���
>,ECqa4 pۢ�U~�3��)<�=\t��!�6������=�� �#H���b���l�D�sW!iFhy�o�W	��FC:�r�L'�h�Qj��#��#aU$��l��r21�`��ǯ�q��j*�m��>��.u0B���]��=՝ڟ#���V��_Y4�1!\�է|���="T�Q��^�86���9��}�ז�����L\�+�`��g�-���H����s�C=�
9M�į�_y��Oi��l1m�q�,�J�e|���M���+Xϛ������e_P�<�$�kʧ��S��_�6��ɔ��>r����4����{�W	$ڍR��WOTѦ�8i@I��-Г�g*W<�u[=�����q2{$Ku�s��oGʻ 8�%QiA�(��1����[��R.H_f�������Z#+��P�jK���Μ骃7�?ZLc�a�55$��W}W���[��̚��0}�Og���eC*��kt2{~Z0��A��fIOB��|;�����7:�ԞL��klGY���hՀ���^AUO]1�Hm��<KË��&�����|�Cj���\�C�;�Z1�ڣ�9`~�l$�UpߦmxT���>��R�Ve��-�Gt�£���������92���9��Z��µt/ħ��(`�Ƌ�����f�a��6[?(��Ԧ�������[Xa�@�m_��%�����z�px�-�+�sw�[�p�IQ�NZ����oǃ�=��20�4�bS���!es��0YJm�e�_6,�Q�ɇ�����C�8W1�o�5�����%�\�Y�Z�0�b�G�Oe%s�� ��=<�E53"����k%��m��uR�II4�v��y҆�^�}z�{�O�e��)�d|,�	�(�[u�E��ۯ��=�~��Zn͝f�r�4�H�qvFy�Y*b��(U�(��\rq�	���{����us�!4��,�!�:��S:�`8����k�TR�U~HQf�W�^7��2���}%�lX�GLKT�͡���]hx�#[�lxiJ�9�*�u��E0x��;��YJ<W&K��R�_h�*y�#��P_�O$n����[?����� {�>��2z\��h��$pzu��O���g�(-IY�A�N
��=Zha{�>6ۈ��g	��4e"#:Eq�(��E�3�����h�dlLZ����.U�`dk�1C�{��9_g��T���O��uG��?������YC1���$>h���_)��������,.dlNm:��H���b_=�p(�h쓈�nw�F�Y�U�͆GS�]s]�W��\h��͎�DV�F��ܶ�t�k�e3���R|FX�W�|o��rV���@�q�ڮY� w���q�7t��Y�>*x��.���--��`	^cp��U}Y1��� :y%.�:�4�ٙ���y����>�oF��-���s1ulJy�Q�v
��и�J���r�=�DM�	���jbX���Y�Oc:}���u�(��_
�څ}�b_�]!�H=]�y�����Ώy�%�-Z
a;r��R�/'�P�Q8�]惮 �6����My��t�O��	�ΰo��EU{��^�~�	sҭzF>��1b0�jz�
�O��|;�%�$k� U�N�Va�Q��ȩ�A��ӎ���o?��5�8b���]? ��`K*�H�6�� �65�b�7o<��*#YҢ��#�c��k����_�[�����k ��b�<W�?�}���9s��F����mYsf�G�4h/~F�`�2oi�����x����$��>�~���(�Nj��~��#���Òی�2�_3������Ř��Y�H���.̄���r[#F��5��
1�+i.�uTP���I�^0^(qO�ó��D����br�OT|�JR}HL����wQsK�BS^l�ȾP|����7x���ss�ԝ�+��PW��"�>���iu�D!~=h���^�`�#�g1ts0}������ù����v�l�����,��V�4�)uG�ҧ��m�c���#������J����~�����2�D��|���_����TpD�ŋQӭ�A#ƻp�R"u��Tf�����U@��i��yz���	v�ޖC 2z���RnD��祾�����;w�x���ޙ��Zʒzb�A�P��P����UA��Fk뎵�e홖��(&�W��=>\8��z|{|\��2��M�<$� ��,�h�YO����+��7/�Χ�e��ֆC�]h�ـ�f<��_g�LFh��J]��yP��-�Ery�͛-�:�J��_�I��-#�c��������&�tҽ��S�9��H�!'&ܼ?&;��h��k3�{"��8��PPl�������)�]�^C�P��� �R;��@�%GEaUqţ��z�0k(ȋ��ҍH0Zj�v�����L��n7��ѷO��$��nqU��n��0|�nV=�?4��CB(��6�-EyQ6�����"R%��J�ئ��6��3H���׸r�^��9��z���hc go�R�H�[����G����[ݘ�@���q�%^�o
lAaZRň=(x�y��2����|^�.��j�)���5*�����$[�+PN�k���G��p��jN�]s&�?�|>���7���{v��m%/��r[7�% 7�.�?�oE�mK��]�Q㼷����F�s��?�F�L/�Um���e��JVP�Z��tc0`4_�?S�h&�S|Nj0!�;�H�eUOܶrR�7q�̀%��Lk�E�Ut�-�.d8��;�ք�3J�Lg[<��*�ry@�{n��@��T1WJ�N+������?���ۃ��ߨ��Er�Y�'}�rc\�K�Q��\r��QA0�S*{k2� 3\k�pR�ҹu@n�̰0X��v�-��W���鑐��q>+@N�>�5>+�Ԋ�ʶ�9�W�^A���8?����l�f���Uh�V1%�w��Fp�%�f��ŃM���<��|W���~i���n_4E�ǡr(L0�PM@L��JN���� ��M+�.��~�;��-h��Fm:�EHH����(�|.���xl��΂����,?T9��՘���+B�pP	��Tk�Z[�i[1�o nt!�]��S����]!�8fc�'�*r�����d37������d�K�dNZ���N���d�!^b���N����A??�0�x�jU9���.QɆ����ۜi]��o�0Ĕ6�������y��>]؀����T�+�6�R1q��~�tPQ��1[�	�n �t�{ԶǭoHi�����9	ޯ��)I�}iƮް�瓓I�)���{�T�qs�pC�d*�s]�F��ɯD{C�
��0�����{n��Y�*�6�X{6�����$W�����U���('Y|�my���(������Ă�a���ȸ��߸�#(�eW��9�~ TC���%�ϸ�u�)�ƕ�'�0ĕ����ϠVO��jW���������k�W�^�T�k���@AN.���>�D�I�����z�8���Hn�?$�ʩ_8ABj��XhH�b#����y��8[��nX��*�jq���dk�5�*R��Z��v&��L�(��@�!�%�<�[�Ll4"�kt9!��!�t������r������?}w��&ڷj�R�3oh��%EY	�S��3})�}�r[�_/F*��a$ʺ�����e��"��3�%�B@���ba�FU��j#�X���|嚜������іEX���Rtv��%�k=T[D	����<��VͶ��^����%|ܲ�Sތ�r� ������tF�S�
�	��9X{�2����н���J���=fɯ��q��o�7<#D�8�3|����Ӓ�E�G!�Y�O%A��̙S>	��,䢋��T�IJ�B�˨�����!X���I\sO��n
���t�'˛�nX,�_lF�|��ʪ��*Ǉ1q^[�Yv5��x���Q9g�n��&������=������_m#���3i&����/jB=g���/ LG��ğ���j$���^�V��[t`�l6|� ��MG~s/��9B|�������������.�a8�|�}�P��D�X�i�z�f:ED �ɚq�u���T���1�j� .u$�֎�a\ k��~�t�Eɛ
*�/�H����3.<��hL]aX�[P�����2<o��)�;\�ml�Ҽ,��Y)kSv�3=3��SC�8�lHX��it ���u��rd.����]��-�cJ��
f/(�s�+�-@˲��D*�uG�k�ӛM�EQ�Kj�W��eN��aK�m�G���`]����!5���&3#Y~x�r2_�us��>R�̀�/#�ź5kˆq�skCZTx���i�����T�9iȨrI^�^��쪳���2�"r� %��nC]�;�:v�����[�M	�Je #�uh�w�^�Z)��<-7����o�~j��_�u���M���<��z�TQ��Ѓ+#�0�0
Ļ���c�k%%��Q��@���-��4���nh=_t����ts���4�D�z�s�ݿ�o�A @�Bn�|j ���D��pnTGV܆h8vH ����6�ƃr�@�ԳF�p׊<�X�'�C7��N<���z�uȜ�1�>!b.lo��M�Y�b�HUP�9*4��1v��w��()d��3��q�1��"��G��`��:��žr�����P�ڱ����J=�E!���|&�\�	#Ur��_U0�t&�z�����<r�(��9	o�R�C���g8/���e?�."��1<���@o�-��><;��*/����C�S�/��~󢳊�"V�LI�s�g�1 �?��+
���y�,b��0i�N|@8�D�;Ś����8A��*�T	[�Y��~��r���?�]�D� ����"�R'3�ץg�w�Ö�7��c�g�A��o�M������.il<����e��1z��m�.���0�VG�feP��֛fn5S7.Xi��3�U������Ks��qL�`�P��LƇ�]�|�<	�.7F%��ZC��4Y������	+��6[b�<5ˉD �� ��������p�m�֗�j�⠖�V��T)���z-���%��-���	 ��P��`ƭ"L�D���Aƻ8e�6����`�|��z��¯��w~��½&/�ƅ�%�EQ�V���7����/��L5�Z3�GL��*�w;J�L'a�d����e�j!��ss��������Q���Q�'	_Yޱ�Ye�׏�!��]�z�Ew�v�� א�r���;�^J��eB�`�ڙ�<�Koe���\Kٯ��e������#��><"���g-� ͺ$cҧ�e�ֺ��c�8+J�H��{v�N��#�F��;�"r"=�O�ܤ����v\A�Ҟ�$��E�$ea#���M��C�����b#��ѵ�a���QD'|vs)}�Ϧ�1(���"@$$�Bo�Պl�\ǔ4��'O�8����'9�9��K5�z�[�f.n�{j�-g�{��b��r�}��gԞ��|�g�ɍ�Q(����}L)a�b�BEz�
�_�X!yZ�X�Th�e�*Z�C�@��V8��O�E:#K7M�\ʇ��Z��묳��ڂG7^3���'j���>U8��1Γ������̠\�е�j	�"�AȕG���Fi�r>|4���3�Cx��
}��g���V2�2��}�}y�M7)��0,���L�6�a5t��!U��n�n�p+B�Z���Qc�USu�{4R���ťK׊i�q��T��XsD]a%���LHR̍R�0$�4���q�~���%H3T6I���i"�ʥ2{��[Zdid���D��G��3���"���VW������Wg�fl�r���~:����Ym�p�4���^�pʿ��b[�΀�U�NB��Do�RwW'�r׍��ז�_G-�ea��`��z��Ұ#�@(�Z�V2{n���[ulŝtA��O �ݵ@���&�I;�����Ӱc�fa�n��m3	��fS �j��*�E�����ѿ�j�s���I�Hi���xDh����L�W<cV�u�[}�Jmۛ�s�{��~��4��dJơ��g���_��[����+9���d7��+������b�����{"�؞��H��lN���4Q�Tz����\�}��u[�J�pT�qv���D>�{1���e�N_����|fd J����5$��ET�(�"t�U�Z��&��C�!�I�4�@8��S�|d��ĹA^jx_�h/�9��S�Q���������A���S�������`*�3��^��a��9X[��f0If��,��m�a����D��P�Vb��cD%"N.��~kx��yݯ�K�D�h��L6KO��N~�|]�V޽�$��{hs��d����P����z˰<:�f�#��~w�dV����(���Q����G������%xc(9�9ӥ�'5-C��9ES��,��b\pO��!T��|�*h�0�ڟ��0���cs̴et��Y'`���IO%��k�cc[��*�䃐���Nq�/�|�$j�I����h��Ғ�%�����j��$D�pm6�\D����k=a`�Ąٛ�� >�K���w��������+�y 6�:�J=փi���K�`F�b(ʧ���f�T���y��-[F(��8�7؟�����M�d�Nh�5c��F��T�`�幚4ÏW����4<]��������	�&.�V�".�4��2ކ=B.�Jl�x�1��-�~;��@�8�異\�����r��{<��A��ו����¨И��Pu]��g��TE��fG���v�J�����0�����j` �-��g��E{�lN+�h�U���S*��t��8-G.����JˋL�i�ј$.GX'Y���q6�X�-["��Md0�c�c4���xE���D3(��}oR���clP0�e�ż�7ݠy����Yc���z	|+�"~��W��'xD3L�mT�y.�vp,��W�V��ms������pnG��W$kn�@�e��S��9C!r�ڻ�m+]�V{`�2�5LX�G��P�xy]��;U�ofL�r��&=�aC�"Hk|sXS9`�/-T��W�Mٍ��ƭz�~�U�q��)�Nt��99����6��G�.G��!n��d��(jr%m2�̪d��z��_ҿ=J��	F�����#@ٕ�����
u��2K��A��'���c�g|��ٞ��koC�3�T�!@uT��H�OZ����t���Uk��@��nt������Ϯxo2�g2�5_t��8h^ų�tCPe�V�=\�_��C�D�w<%����':�W����d�qvU�FH,0�tOǈr}p��0�]���L��������T��P�EQ�L*>���${6X��|����RN�����ĽmPA2�6@�!��G�՝��V��"}�ӷNo�j��Q��%ڲ���� �>0��_�n����c'��B��J5�{���d�����~SI:!��7uuɜ���x!�nfT-��+3M����.���f�ۡ�a#?Y?���$�i����7/���*�+�������h��My/Mch��t��O��I[DOT�,�)��f:
}1]�97O�"�LxY�x���F�X.�ޯE�%�{�V�_$"x) "�,���V����u(mxm���X�'Ŭ�e��md�_���\�r�F��U��(8.�����n��4�6Ҏ�2v:�'2�W��:�����q��TG���)�����eH�Y9�I'�D���Y���'B�2{����Nϩ�2#"źݹ�鹉l?��N��^(&O�)�֝�=�$��ƕ����b��u�t(��v 4�h�i�|ݫ�_����_��:���$:��jE�f����c[m.�`�I&@�+HF��5iO�������� ٮgTw��nW������� �<�zXl6#	�l�)��g�&$���q��<�-Pb�A|e
��1�)��"�9gn��1�_�$�}>�">��f�N����Y�o�i��@�)��w��(4l+D_C�5�o�*p�lQAjM�p�OAp�-�S��>���W;���tt�����T�A���lE)�#[p*��g�q���A*�aV�ж/h��� 	����y�!+,A�3*n󖂑���H��׊Q��"h Y�Ƞ#�9z��A<��6|�S���H5*�Uu���3+O�����#�JY����9�`�a�$(�vֵ�I�n�� ��r���eWL���׻�p[L>���Y��J`���|�c��t�R&p�-��)O��dO|�	��5�6�#����C����(�:1):�r��c�l��<�Ne���!�<`%�J���ZKԔp�?���`u�IC�t�`v��F��3��ixE"P��	O�6��[���JYٕS���;�b����Q5ut�[ ���~���ONR7u	����vn�us{����<���n%�$�����δ�������b94��ļ~Q���N�>;~dN�oHV����s,=2��3�Z7�^�u
ޖG����bzb�Fh��K1������@B�g�U��8)Ȳ�ᤩ�
!D�1Fy�O;g�p���+{qy��;���!W���҆�mB����=��&�p���٣m��݈�D�Ϥ�s�<"81=z���u�lp�5cqaA��K�F�*�=��:00@���e�� �:�0eR.�Tb W:I˃�#^K��؅�Ty�Vs�3^�@�яC��e�!C�Ǥq��Dӓp�3��� �}'���7�e���ږ�#f���qJ2'#��{b����j�a���zyi��ӝſE.-}���V��U؄((<��cB������l�|�V�E���D:eE�!l�͸�|��k�{�&t�x~��(�'mJ屢M�$���JpY����x�����������r��<v��h���b+�J_�����5Oi��/��3`񵱯a2�$x/�ה���bҰ�b����O)��D�s7\dE����=�Gc���S4��6�����rsI�veG�\�ݤr����� M$.p) �8�����h�Y��O+!�o\�ot��{ L��k�}K/_�w0�w�ޢb��۽r�M��?����o5Z۴�fV���2nA��n��	���(^��eMs�S���MLll�spYѪ�l=[�v}(�j���\������4�A��w�"�G?����a�eLz%�Q@�ڻ�Gk7-k�X�d�
C'�� � Đ��+˩�k��L��z�Ԑ����\tY�f�x�'�w�]]�	8-2[����o
~��w�;�A�i�ԋ�OE� ;1p,J����`N�z3�ؓ5`;�V�ּ0x�e.����N>]w��yO�;m^��	��;���nH��q����~�9m%�=F��,�I�^�벥)d�N��&PMZ���;�(c��ʱe���ND�����F_wD�0؆��s"��}xg4�h�`έ�-u�ۏ��
���Y��&�F]�3-�^իg��q�~�-����q�ׄ	R:�	/��M���Y��n9�b�?5������	>_��J��d�4.n{s2��)��x�L&�կ���f�ɧ�N�}��]"���f�����^��#ީ�W/�L��έ����O�Hh���F��<-�غ}/zyG��x�@�v�d%�5��DN�4�c�Qsg�^-��I_J��Ht�<��)��J��@��l;Bր�����R�G7�0�Q輻��B�X�<"��F.M���?ZQ�����H� <1�T���J������X�([�d��ϊy0M�ނYA�R'sL��Tl��S'k�mr] <}���rG�kZ��6����$EV��+��Յ�a׸e4i����)��)���{	���%��U�r���|��z���	$y1=έa��o��+��R����! 
�lUw���w�wA�;B&B��$�Dbe<.�������8O��>4���#����(��M��b�:�(TW�<}o�~k����=OSd:e�W!���Q��,��K�>��S��f�����{������l��K�^b����Us/�ӌ������|�ec���au�W�r�tg�*��x�;�PB���E��^HX�1�-OX犦<�n����|�5Thm��Q�4�E��y����EU��^�ѷ�ճ�l�)���+���ߩ�ӝfF xT�QeF��!���x��aAYU¾$Hc�M���m���4��i�V��
ʈ^��V�r�i���/�l��&Ι��:�罇�l��:�����}xl.�ٜ����(��L���9�
��w`�F�9嚞?��U��C�$T������X
�hI�t����=��H��������;�M�z��*}L�x�sP�_�h	J��U�?rad6�;B{=?G ��
��c��	Xʐ�mE
��r�_-CY�)i��S:����i-��T�9c���3wD�z���ŔJ$J�'D�p��|l�o���kp~�Q�&((�s#�b�e����+Ȍ:[d'ڐR��G��tjD�(�ؒȫm/JF�y�JRzS��ֻo�����Ż���A�W���6s�|�:��Ҙ�׀t�,U,V��Z����T�Rj.<��G�S�F��؊�̞i��#j��]�]?�6�H�Qv��/��x!��y�V,Q<����{n���W_qyN3{�¾�s&��/k��b�R�����L�h���K�1��� �0A��5�/���L~�<�G��	��D���\�U���TuG�wSy=�A.�[����R8N_=��ύt���O�������v^���%��L[�	࣯T��|��DjCZxb/p�R���zs�����]T��7.�J��|y�9�,��3��i���&��i�ƛ����(���kj�̞m�>��ŷ����8�]i�U8��ҫǺ�TL~$��ġ�);�g"���KK$l`c�Hm��|�m}�=A�>5�f	{`\����/#l�Gy���/̤A@t?�B䟕�"jQ���2��b3��	�A�}��{)1Z*�;�Cҩ���(kw�?N� VM�k����i���_1/�m�>�7�(ʨZ�: �b�[�1��\�����ӻ�l�~�9_ߊO�	���	��������M�3BS~��0jT��L�����*7�x��;���c���(�cK%s�qF!jg���ۏ���d�����	���	�R�|�fU���8���Btr�R�TD��5np7?���mj2�Ve�G#�����7��\;�՝�rQ)��q�5���}z�{T�B�sQ�hN�M֑��}�t�t��"d���Ĝ�4L�k
�pV
�V��|l�h�.�"���tY��rH'�U	C� =�(�@xw.8���X�:��s!��2�R)���e�j�s�����{��IH�IG�킛�t�@�� ck�Qǁ�
MMMf
+��Ն���9X�P����<��������H��F�JD�CPʔ�jX��5�vhZb�8Ā��~!T찗"�仹��v��(�ʆW1���c��L��?~^����ହG��P�������;��x���xE�� �{9R��	B\p��p��(����vݲG��`�`���g%Z������#iN�e 
%E�\D��6��0�Q���ܑV�~�������YY�q�'{.��(j�PY�J��y�� �9�*�0 ���eRD��v[!�tlt8)���ϣ'q���]Ѭ�N(G��x���B�``�����+���K�D�����\�!<�ڞ��.)k�6�2�n�I)MUԷ+!�^�c��StKa�c������z'y�cv�q��A.����!�Epd7�e=��k+_t�ΐ ����vَ
��8��&��*���Ԃ\.���O�8�"R%-i�m@�z�R��=c������M/A�}|ӎ�����|ۘ(�;��s�
lH��@�����8�c�@ ����Yz�71��Bj�V��7�>`�0	��H�Ǟ,k��T,l�*�Ą~(TXS֩�X��,���X�+#�����`.����X T����R��1u*�W$!;���c\m0�~E�Yu�g*@bz���y9�R�QQ�I���o+7-��<S}&Պ�Y��ߦc�	~��[��h�4�	l��flf��O�u�`xؿ�K�ܵs&VB�b.��'������P��1����|�Z�N���[�2���s�~4��5�պ%6y��{��kZ@;ؕ�>2Տ!_]��_�����0�����2uU@�����y��v~�C���tuڀ}����Km�SYݴ#�T.uH�6����@F2`�4!���|+������:=��`Rlч�^���pI�Ċ�XTb�.���1e�.e[LFm��p�D�s�sMUF�,�u�K�~N�1x6_�_�Nj� ><�8�\RM�Y�K�V�}I{h}.0f	ŏ��? D.PJX��)�}v�u�H%����E�5�/
(���H�v�S�	�dS�	r�I(��0���Ee��.�f�e��n���E#\��[�?j��$�۞͈mȗ�@�0{����4�$ �jؔxi��4�j���0-�`�.�：��Q�)�3S�w/�Ľˎ,����t~�T=�f1�A�v���AٴZ�Wp�c�w�	dH�6gyk�B��PT�ʷ����ٹ>���x������9 ��~�
�0C���)������v����ͭ�����VT�<�s�\u��c��E*e����6W����XA�U��K�(K;�q��9��u�ޠ{_�	o��LH�rS;p[��Z�5K䃖��%S�Cn���:��<t] 6<˫~�/�����(A�33���`p�b�SGP�"��[?��*	����-�;���m� Y3�V��㌨N�P��0�d��o^�����dŝ���@#��\���j�����{�d�{��丐.�Ɔyw�RNԝV��&���R\q,�i�7�H%p�ET���h���!��i��V���f`��=��fE�J�[��$m65_�#M�J>Zv������P��W�A�"��ۋOu�=p:+D��ӹ�^�����Z?=�"�y�Y"�ȍ����,�+��-��"gJAAC�u�3 ��'�� f�;�?�]_��w����r��e�w��W�ж	ܭ��KG����*���`�!�f�����ap�,k`_��p�|!��ch�<�b�L���?Љ�|���§ ��܅�\�O)����k�5.��K�>���rI���&��AW%��z���ZqTkF��5$����2�]1{�p:u��u]��i��E;o��AV�?��p����
�d�K��4̤0��������c��;� �P�. ����X�[� E�V�i^G/ed,��r���5f�YF���,+�CV��m�.����X!��[�9�Yr�}ھ�Hs���j\~i�๱CW�3��c�ně
����.j�2�s�K|_|K����Y�Ҫ��B�)��b�C����_R�C[Ԁ��r��%�G�sJ�mf����F1���JRp�Vp��RBk�a}�6��L�&k���Hm�M�F��׊D��t��=l��%<�nb� � X	�4��L��ť�pï�a�4__]O�	��՞�0� s�򞕜�8Apn2����3K�<T�=�S��B�t�}F���m	��o����\1�^�@^��0��2���#�ÃA�<�AQpcZ��ωG�C�@��>�u= r���Y�!L�f=�2�ᕿ�a�Ґ�(��p@������i|������4�ao�Dln���ϊ��B/]xL{A����tW\8�=���g�{��p�˴jlv��%Ԅ�Z�2�2��	Y�8r�ϼ���Zuh��I�����]P���Dpn#)j:�٢�5Z�/��G���T����js�R�7,ew���:�e�Z�Z��<��Jq8�j`��ޙ,҇�NP׮7nr?f;�M^��/�%}�ݍ������X(+`��6��4�˅��`+�&jj��C��I⏾,2h<��a��f���D.+7�g m,�t�gN���쀤V3�l���}����B֠�"ӊ!LG�լ��1 �\.���]����-��v�դ�=_a�U�`EH"�ؼ)�v�_*�R������$���p��zfkÊ��ko�'�L&�46/�<�>�y��M'n����zx��n�E	N���*B�{���?�-������� ����EE�A�@��zcoL� ��c�J]^~��<ԡ�b��7�2�+gj?f|p����,�.��W��(�b��_�T.X�ј9�X-%����f�co T,\��,;n���3����=�H�C��;?��N�$8x�ΖrXQ�����"m��M�Y`G�h�����f47��.��q� 7���d�.�ޤ���+;�M �!�<"�zV�k6pԯ���w�Q��ܥ jc	��]�o�n�4T�)����N�6��D�Ag<"UC�9r(}
��K��F-&z�����YZ�b�c{�.��{���q^�V�8%9�A/_�H-<�<"ή�X4��Mm6����㍼�-/O���L��6�g	h��Mz{ҤD�)�<JL���c��p�z!�j������E�I�$��P��`Dp2����	�ӏsU��=3���I�%;�u�LI_�b��`�	g5id�MAY���[��Ĝ�rGR3�c�*?��f��5��Q��(u��d,��gL�2C{��M� ��9���f���QL`�x�j��q��1|�Lp����H�Q�b�s��}�Q��{�۲������;OΣv�,f���b�^��״�q�.hJ{A��#R���@0�[i��id�g�M�}�Gm�d����BHt}�l"C����sݒpl��ǒ�Gi�N�+HJ7�i�{��lR8,�{�3~��Z�ͪ==eO7���_�
��dw�&p�u`�Sl��/��<$���Zn-�`+�n߃J9�펱��m��yw�Y��pVUV���>�I޴�NV`�N�3�n�g�d�������4��%�\[f��mٸ��-�? ��m���Y1�邴�P��z�E8��L��'�JH�8��9N�s���qം������*p{�� n�U��������Od�:�}�J�]F��[�G�J�L*T�W��{V��\��b�-oV�b�S J0
iK$�Ǩ�{W�c�~�
�9��*�h�E���m:�D%�,�p�e�;`�d� ����AӉ[��:u(��;*���	%�U����]iX�#���o�F���]>��N�}UXD�sq$�+�y���
��*��?s�!OW����n�Q�ͣH>�,υ7M��ۙ�D�~�g�mY9f}ՄV���S&��8Vޯ�r��ʹ�(�iQ)�����ӋVb���/�5�hr�\P��$;5tL�z�i�p����l,D�t�40��)�K薓�`U{���GA< ���C�(��t|��[.�B�b��l0M_~�Y�>8|Y�3'��vW�'���'�Uqt��X���seƍ�	a��W��<Q9��`�GTc��c,�����/=���SQ�D;�A�O�؏"�T�,�R�@�|a�l]�j��|~i��k���@z1���}�,�]VXP��b�J��w.��պW�[����-����l�w)ռ��T�*n��t?j�s�j⣾2��m��>���P�m9>˅-�0��ݐ�FLJkc�Mz�DW4[�\���B�ۂ��/����)��{qz��t���b�f_�$��������\��d�q��~+�A����eӊWT<ÍՠE���k��ï���w�'���[Q�mUi�����זAh�����#G��ցڽ���/I��0@&h8t{&$1�&D�{���Y�R��Ц��T�c��f���m��l)%?m��B�g&���p����F�(�{��q#�ɮ��כ
��G�p �֊�j �WG�j�ۆ�{S�������sr���/���ӿ���^gg��7��Z�����Ы���嘠2�?�!!Xw��<q?�y��+�'�K��z�򜶽EӤ�MK���A��n������P+Q}4gW1�Fb�?L��lS{��)�٧��� >5���gg�I`��5��jo�4O�d9��Ƌ�#�t���;�k��|=��C�3|У��t�yş�Y�!��s)�a������<�Q~O�����f�z�ru���V�~c�)���ñ-g&�������;C��$���@q��Pܛ��U��x���6��{�R�@�Vg�Z��X���F���x�4]rW"�E�"�4�[\͑��B޺�s4�&��E�,�و�Ϯ� X^�X���p�睇���8��ȇ�AJ�j2�ێw(K��L��`�$XG&(��Ƀ~)��4���K�9���ZQt���#��!�[M�F���/TZ %�f0K�A���,N⃣�����St��4S�Td�G��پ�5�[mr��C`�*7뼲8�l�{j�����>8XP���-���Ѷ��3ȧR�7�ܿn�z��������3�ȵn�H�(�yJ������_��#C߿tB�?�B��Ⱦnq��B_��o����w�����g���?x��_�4XG}�%1�|/�x��M~i<������l��P���E7IL�-'3q��{"E��?.�������(�����ѓ���Yխ/���U����S4�rS�^�v�!�y��+&��w�)����O&���~�'��������@�Ƕ�$�C�űq�����&P�80=�'�ۂg�_N[����R�H2��R�7S{ �#�@���֫,`>����,̒�7WʔD���-��MVdA�����-�3P ���~�Q6�"1�Ǽ� g7 [��`-	q�!�*�wk���D�SŚ��].ÊgDtw�#B�y��+ړ����Hј�C��8V�$ye�jVE��iH�	��B�(ј��ѧ��ҜdK?u���ǅl�5��Bk��/�Jޣ�v�ď��[��ω ȵ�`桖:��sPj�	.��y��$�`Hޫ���>&�`i_)D��yq��P�oB��{��Itę��N^�e7��:=�Ҩ�������� N�Ug�0ݾ���֤�Y�$�6ciԦ$D�;�jM룼AGRg�q�Ǿ&��s4[��?!L��N��Nt�8K�%`�P q�Ƭ3E]<��Ǩ�	��a1�㛪ּ`}a�L~Te�3�5��r*��>DA�UԳ-�w�d���:Y�� �?�w�8t��<g���P·����+�=^�5�,Zxo�������gr��	[�BZ�<�#��g"p�Ɔf������-�&;�	��C��a`�E5��H�,�fXʦ��	U�g�J2HH9�J��2J�:�M��ͦG���%���o�����#��@f-��N8�TFߗ �i G�/)�fn�Y��GybIlLw���M��:�兕Z������Xj�B&�Ob�=w�UcD��̑N���������]�����@�����"64ټՕ@F����q�M�y�_Q3�\��� 6�f5�K	y���u@u��`)��dI��̶s�f!��)+b�X��&�2A���}�������iݾ<R#�}܊M]�_��VŇ��9�r�xfx呟�+2����MEjG�74�dKp�U�����	�+j��+�� �|���ѡ��2�(��}\�A�j��oF�0����j���R���d�T�yv>Q0p��[S>h�N�~�E j_�)y��'���RyH��/�w�k���J#�b�3v6,P�r�'8��\5y�l���ٓe��B-#��c��s9QϬA���x�"yQ�����+�_�P��r(q�M��nw	�;
��Z�-����b��]E�^�lj�#��0��w9���w �,�����L�_�5�ᐵ�"' ��ԡ�V�4'[X"N��kqCdF��Al�=����#�}U��ss��^�C����qШ4C��ߥs���/����;Bi{����b�N��p�� rP87n�Y��`*�1�_k
� O����fol{"�����y'_@d��t���)��~l��Q�]h�� �\.��Z۾op	8�ag�[�eZ���l��M�a$JD3�S/�6G*<�F޸Ɠemq�B�d�K.\A���<K��7����exPH�y�<qE��B�RR
��@R$�SU\^�v���_�Z/ٛN���w%Z0%�<���!�E���C���ܜP��'J�Q�r���e���,��U�m^��W�'D@/�y֢\�w׽Ö���t�㪶s-:��{��(��B���"��*z�%<'�t_uR4/��6�Td7���)@���
���b�^�Ffd��@z���X�a˪��+��`�VZ�ݧ�Z/6��xn�͖��PU.�ׯ,�h�4���ӧ�Ol���m�8�l��n������	��]��x�I���˶������E�>��K�D��<4��0͠�d=��FO(���G3�	+�u[�*�z?��f��U����c�'�g��KG<&
�R�0PF��(M�j��yS�͛�sP����GOV�Y�\�誰͖�����D2��"�p�,qDE::� �>�堊�l��"#�II�?"��]TH�����rU]aP
����]���ݴ�H�&:��E[��m�`�<����&s����_��4����C<���{`����x��q���o����K��%�43[�ǑX��ھ�<�%���]�u��ʹ��. s�R)H̗���/!��}�	`A��b��/��6���e�����F�;̟����ka(G1���ِ�s�j���e��位+[���	ٗ~�g�Vo��\C��i�oRwq��*z��*��sɸ���
$�~�WD���Ae� �y��Jխ�*�'�7vq*�XZCf�]�~�[!�x�+ۃqǳ���Bfr80t�1�������c�������y�c���P_4����	�	��k{Dgh3-o��A w'-����[ˊq�7%���
匯�׈&����$�H���"��t��k� �˜�FP���B�饹 ��x�=��b����' u�����;�E��#W�UU{|3�23���N[qB��0\�U1q=?�����C���$>y���T0㞴�d�V�I5k�4��[�1}5����;�aS�N�z��E<�W�}[b�%#��b��I�X(��D�=e��G��{�t$�����X�Uц��s:1�R߇����p���Wc�Ӑ2rd�2�=��v�7$��h.���VCt�l�L�V2����O׷����j�IIniF;��v�F��J�n�m��Ԧ�`�WH��̴��+�kꣿ��#�<�H�#9Ō�C�B�-6�:8�]��z�`IK)��Y�=�k�9<�?�eN���8��zN��HxQT�������������ʜ��+J�B97����Z���^����5(�4w�XqGC"��d[I�-�%�evX�l��_�Y-n-��d8EWE��C���k�e�i�֗�{v�c+�]]t�Q���@+�����{&9�G�>�:���P6]��ف�4�Z��)J�=|佩��Q��!T��(K&�d��cFeJ�ָ��~&N=�p�	�6ͩ�cY&�*�4��]��]�&5�ãu��V����.�$�aFr2⣩Dm/��^�� �\d�"L `5��ʑT��x�ܸ*o���iGSs���� �`�JZ&��hN�W!%��y���#T���I�!:�̂����Eq�|j�r���~g� �:	(;��/ci��}��f��:F��`���i�?	��-�)���A��4�wl�HO}9@af�L��"�!���|�-L��v�=L�X�����2�h���w�H�բ�WX�U�ؔ|�c�6w�7's���k��*�s�]���<n�qM�#h��[h�N`�
����c�O�&e��@��6���u�Oi��� b�P.p�"f��>�>v ����q��K��|(��.���Sy�2n���*����ɚŪC�^������ݞ j`HV�d�|#v�_��t#^�J�ar���RB�3�pG��_�:p��skB�K"�3#��i�L�*�����%ʌ�~e�:?��Y�*�^�nſ����%1�����?H�N�ʑ3\�QL���d���O�$'k��[3ü���ވ���e�����O�es�=T�uGK�`�M�ww�������}G��PV$K%'+�h6���kᨃ�)�׭�«�@���b/����Gnr�Y�B/���(�q�;]m�"����5[��l� ��d|ş�pO�i�أ&ƕ�i��x>�*�Z�Y�POm� �A;�w�=�@4���{XjfB]Ɗ�x���e'͵�T�l���%"¨��H*��.�X�.�0�A8;�hDV J��t�31n�׺"!-Tk�AN!��z����%PE������F����g�{G4H��=������2��$�a):�P��ۿ��������4u忁��Y���5�&�%&��S�T����pASp�����e_�����{%}��\!������NE8r�lE�����DZN���
|�F_�ڴx�(u��`v}��� =z$��'���n�\+��� ��釜~�������`k�X����^S5�b�'8|^�ey=V��E��@��F��ۓtY��ĕ�7"ب�ŧ~��U�1TZ��^{ǲ�� O�Q+5m	,��%�+��G5^!�*�d�j�=��P��2�[����"?3Dy'��ܥ�T�������䏍�KI���CyV�U	,P�7��ݐ���B��:o��恞�^�ȉ@�Ϣ�`U0^��Qڵ������+v�.+�I�/y�:x!cd �m l�C>�K�f��+^��i�fSܾ�B�0L��͵	�?7y����b���jN͓����P$"qBҊN�H�%�}
�o�o� �5G͝�x���ܺ#)�FH�c̨~d�� #F�:*^�'��mi�{�������[h��{\跕�ì[y�d���j�7h' �D�u��Bߋ� ��h%}�ʈp�}^mlL%p}}oW1?�w�Q'���C�v1�˓fy�'X�g˂�}"���J�`,��w· 7��^ߎ�G�CZ�6�
ʝ����Hlw]#˻IAdi�U����eX5��~���Fu?��}/f�^4��/��8�]�F`�?�s}2� m�!(�s覂�|`=kcX,�;�1� tć�q+{�h��)"�.�9��f�K��&j�3��U��%n��Z��Y�����c	�]�����Yt��rф����#MTܴE�VG�����Ƶ�*s����7�/��~�[����z���t�Sk��W,�qG?9��LB{�C�������NУ�b#�B�f��ljoX�LL��_]����j����~����&˙��@�=�*��و� �.�j�����.9�I����o�R�Ճ�Z]�B9E*���9�[\�7$ @��WP�k]�o��a��t-~:�G�(n�V�.������Z�� A�6�(�T��C�e)���iE��8^ �ze��-��F����r�g��>3;���ҹ�.R�X����o�4r�b�%�rض���:�����s�W�M�0�T}�����s.s� |.K�*��#x8�4���������/�ߡ[U)ů hYA�]~}ft���2���MgJ"c�B�B���c���q��FƙW�;�����;�0t��c�浜0�O��e{��z?�x|�&j�rG�-'��1��P�m��Yv�O�6]?&�Oh�,}Y����H.'��3A�qN n����ܪ������M��m��P+޴�di*�)��R*S���ǏNpi��[
r��O�aX���Yצ�E���|���uq<�ªvi�l�f���Kktϖ4V.Q�ȩ�#��f���7�~XZ�������$��E�;*wP��ywm@�����N��(p�f��a�9�#�i�,�y9���XUu.&5�6�O�j��s`�F��ޣr*r1 l���!2�
�� ψ�5��Em�AH�����^�]$YƘ�z�Y<��y����u�*#&y-t��ٚ��"����ƾ}@,�G��6��m�i��i�$�fi1�>ΓL�URQ:䛈����
)r@�&p?:�=pBJ�D�S���xtXV���;.��e�N�q�%�ig ß8\�g�*�'<����Oϻ7�w�n-�d�a�����<z��~ sE���bĊ^�����(!��6���**͝���+�v�WÃ�v��)�_�5�G�(-���H��Y�* >3j�"d��c�>ꡃ=��()��
�p5�pô�U��+�d��ƻ;�<hq�	��w��T���[�16��2��P(�:�4�4�^�[K��q���<�I%���Nxpe:�Op��F�#&�;6O6
�w�mHw����<Yv_<퀝5	P�o�L�c�	�l�@��Z�~�%B����nA��V�DK��}+��o�	�d%�@q5�s�%��pE'��̱��ͳ��I�s����w�E��5�#�����I�D��_����ԆR����I}�9��x/Ì����6~����l��E�,��7��h��=g����CÚ����O�9cl���o�b5.^�r
R�_j���XŢd����Oٚ��=�ڠ�c���Y��l�[,���0�ɫ�;�Q�0p�U���#i,w�S='Я��|�?���������޳O��&�_X���B�R�2���D���\���+B�5g+u�|�)8�rCp�Ĳ��n<�K����/,�����l%欂\�Pbv$�j�D�"��۳�O�'7���l*d�bMs�y DLɓωA�kzg�
�6u�n�T��L��<���a��L.ꘑe�iҤy������Nw~�lh����a���u�im#�
	 �s��E�B{���8��.� "��&/]%�-����)
�#�۽�ٵ�;b�mBڬ�h���U��y X�y���7��LV2_M�^J��zi�ү����a��:Vr��r���iڔHg#�ɂ�C�h��)��[��L���X?
��������{4�O��]1���Fy��'�*��'vuq�v�/��[&��)]�O�9�#�88ş��3��Ng�����.	�c�~"f�*G{�6������zz��e@ŀ�`������ ���p��)�_c`���I�8��&�������d�k>����(2�zs�����K��VOo�ZF��/�ּ73���|�^կ��I!��K3��ns�̉�"�hW���)�j��<d���Į�k���u������-ɳ���P�E-N�GC� �ʜ�D�ᭁ�A۟L ��xA��e@{L�;�)NG�V��P��_kZ(`b�A�Ჰ���~l����؛Y�͜$.���3�/[M����	O��gp��)�����B���3�LQ�0�>ek���RyUl�E��)���Vru�5�݃����I�Rd#��+�s�p�9�#���3���w��.S��`�n���l$/�YA�/�y?)-wD�rm�~�������N�T�ֆ�9���%R8Ecr���̍5β�	�_�4��:�����	�ar[�eK���L� F ۡ4  �5�l��Be¦��g����ڄ򈾘�ǲ���U���E�l)S��`�\ԩ`]w�Cגu7���;����@������!���k��-S6Ơn�B�z�%R�_~c�c�[De���}��E^���6�6a��1n��5���s��Βj}����L��y$�/8�Iul�q�o5-i��!C�N9��,�7�Q�u�8�.0z9�����4�P��R����cO�#D�[)������K����b1�ּ�9��'
��
����&�U< R�G�14����o�Ps���}�PpT�2!�Z��:H��r@tL��Wb�*����0����Q��m�!��z���b��c�׶͙3|T0�X��ȯ�ƭ���d����5���;��`��.�7VaϤ#�A�piW��-�Ч}��1|H\�eY]���U�4Z��h�;����g�$����1�z5MgĆ�gkM'�[8
����J: �
���F�dܗ�Vf� �1;�s���=��,6�uZ�	�d
�6#�Ex��V��G{g�� �����c�k$�M���/b%���c���3,����rG�G�DvR��8��uc�ݧ��F������x�v�"�b�x����|�O����G��9�1�sU�Z�\#ɇ��w��tY�Y�|�m�c	�݄4Vyg;���ٴ��䡴z��(3
��P�*�����"ƽ�[b`�D���ԝ��p3�v�o��N��Rl���f��2#U-R�22�	�G�W���6݉�zh�"��t�������ST���˱�sm: �'?-U����"ui�*���Wb�/��M�/]��6A��۔Gx�O<Y�P���%�� ���'E��Eg�&��V�������0m�Ʊ.P���!)N��{���9��H�E��]�3	�,���3h��1{�U�ODk��U���y�z��4>�q�涂^7$���
�_��Ê5^zZ=���9��z�,��#4�ʎ�D˦1 �s�30�{6W�3��%�@����z8�sW�w'������R,��yֆ�Q	������5HM!I�O��BЂ���(T�@	�����<��Ճ6ʷW�G�e��D����N��uZ��HL�~\G��-�m^�R_Z�-d>���?L���IRZ��WEW��lєR
>,�6$���])J���*r�<�^�6�9쯮��q��Xp�(��2���N'%[�����^�O��+�~�;������c��?�\��[%�R=�p��ʞ˾,: _X�vF�" i:9�]ܮ���+����w�=q���Np�o�h�lO�)\�r!ܺ5���&3=���o/����k%#\(�N^�a5a�K�F���b$S��UD��4�Sb��ٽ�YF4�>"Pom�W\�?�(
�GK%�)�w�c�2p�3�[�r���0˪���_w�c��s�q�1�2;��3~��(��J�XRS�e�z�����ǫ]�c��9.�Ѣ��J��B��h�Q�79g�$�)%ϋ���)��`�߽��ö�g����Kn�<_�M�m�Z���;��L��������ҒT�n��b�\zJ���0�.�7�j����g@8����[եO�����ĸ��8��N�`�:%�ȩD;*Sݑ�d�bv�"��C8T)D�_[M߯�yv<q%�H��o�3�P}�̈́Ȗ.�T�)��/�{�<�l둽D��o���������P���ĭ7�b�	��\��l>fnC|68��[�Y� J��fM�?
��#�V�F�r�'�w���dZ$ֿ��\�=�q����J��@]��N1�"G�/��I�Vh��&._���)~ (�LI��8���/�d�n4$'>+�*ɧ����p�q�a��C����<��W�ޕ@L~]��v���,N����5�.�2 @,�����1>[9��Z������+�h�m^�mf#*��ؾG׿�3a; l%�3Ȕ"����]�Ǣ��!��Q��+����0m�����Y���9��T[IR@muR��L�qt�M�����'�3"=�Cc�n�,�#B��՟%'5���v���m�p�@Ip���U�<K[n4>֚V�|�[%�q�c^�vd�\�h[3�gO��,��ka#�<m���18������̖}�7k��Uf+l��ɬ.�j��F��xum��r���k�wq�w��J�Ct["�ѺC�q�B:���SLd���&?��,��Y��N���I�U�:�P��)Q�mOӇ�_?]����z�jr��lP�Y͜ΔA8�ss9'�ջfgci�t�B���e�w��Ll�T4ױ�4uPwow�!�ӓ�'�Z��E��b�z->�P��lM�]W���3���|�w���|��S��2N�6?�钻Jh��1P��?�65��l�E�Ԡ�Hу˗���=ݷ�%i�l���n3�:���̦�1�{�S֮��h��\�[Z�?_1���w�]���J0��j��,c������tMΪ�כ��<�zi��-���ߛ���o��&�Vt�� ����٪�"��,mz�����5k7T�.��CH;��"��#�����,�����_��t1��e��}�{��J�A�gEV�t#�6�u��`8=��l�k\b���-�.��Ɵ9��T��
p�}��S����Uq�^a:3k���9���������*�����H'sԎ[wVg@�(�N^2w^f��-�&�QuC_ᄷ���_)J�i�!7��ƹ	�����݂#j���ɼ�+:a�?��6?��z9�s�g'i`4Vt�bҨ�UN�7��Lh��T�2Me�;�z�M�\&TIz��<���yo��;�8-=4��qm�l��k��es'f�$E��=!���˞Nև&̧>��0�8�|���ϩ�g�*-'}��Y�F0�n�����E���r�k�X������	S��	Z~��[��Ov�W�x���ا��5O�	*M����Wh�u@�`.�x��Om�+����O�&��L�2�	H|�8p���"�;�먘�17��Y�}���8�����Oi��5���d�)��+FX����t�/��1P�m��g71�SR�t�����`����'�ҕ'T��nt�%\�譶��D�g�	o����2�k�J�%][	Z��'�cD�摜��I��7z&=�^/�3Iѫ�E��g��H^�x!)��
p�*L�5�5F0ҴiRw��s;Uy��{nړ��BC�R��8��v����Ifr���y9\��_�K^i'�1ХU����U�;�7'��'�|2zQ�z��B��IW/h������"B�E"��u"�a�\1#(_�;���NBÏ&Tݩo�i/�*~�M��)�{��&Pg�����!�`�P�����#e��r���l}�_d�7��N>���r����ֹ�㓎3�2uGXٮ!�S'̮ʳ1u�颂�L�j���=&��2��.jO���:I�!�N?��l�	B��][��i�[�r�CĎX�LI@��.�}����,֌f����}QL%����@w�"�)Ӻ�JA�	�y��;Й�@������{�!=�dj���IN���~�+�&�a��EZ,֧h�������Y;Q�|�|���GDԷ̝�p7w�aV�L�u�x�A?�u�y��XRL�������g[�n���!A�F�F;���=�¤OZ����p�.���^���{	����;��JסL��ky`ג|*q�qch�չ�͌��_9��*TU)���ص���[9��=���J�Ո{�>�i�ǼўX��Y�J��!�f@�Z�`��0���j/�/�i����b ��:!O�_1ѐ�'���$R<�s�>c�Ħ@aÀ�<2�~�^mO, �oe@H��3�d����΁z>�M��+d��
�6_�&
m��qM{�#�!��-����2EM]<~����+�)1�������ڤQ��!/�r��1�HJ4�'nZ��t�
@c@��Ŭ9f|�B�g��5����{eP��=0�}�"��u�l�u�k�h�E1�}UF�l~3tp4& 'ʄڲ��QG�g�H�2�7���c|?�N8����{{ʖ�N �^�k[ۚ��?����m��}��Q8�V%Q���z��.�\8�{�ӗT��o"t�d�1���Gnq�+�V���tlX��_��ƶbL���ۡ:��	��Z +)c��?|`iwE���!��#X�16LT�X�╽i;�\��Ѥ���-��}�9��8����7c _�0~-�U`��x���Q���\�I�4�w1����@�O(W\;���@�·;g�����X����>�<ɛ�{��Ԛg��&��g��
�q7>mr)n�4�`60�sO?s�p�x,�,�a<�������TY�����J��f`vM���":��Ct�1t�D�Tʇ��`'GLLr��߰�(�_��N�CRS���)�����{�6�7^YCS�wu��9��	E�;ؙ�]>���_-��������g���3-�V*��۱RVx�����xe@H��:ȇ�xdb�������#o��+<6 2z.�����`O%����=�0{���/���Y�w2�Ĺ*_���a��x�ɦaE�R:��@�� X�L�Ѐ1����x�2+8���r�Z���K��Y�~փlA`��&,Μ8l=�/YB�Lظ���kt�u�T8s�`����sZ^k#�c�ZƦVx�(_qH]��(����L{��=����+�.�四�#:;R�&>U�V��F�Sc=��L���f��$��u>���s�x ���b1���
rt�r��c�O���읇B��9����Mw�z���8��Z.	=��)����;%q(,d�-��3X�JR_}��:|�4	���v�Ϣ��(��:�Xš�K2l��r�>H�p5�~�K^ҁ0��*��6�Pv�k%�R�<_� �h�Ҫ���wI���F����I�Kx�
`�t�
}�g�46�[�J�a^u�`a����2x��N�'2y��f������$j�a�P�@937��G�5=���@�_�A��A����\�@���J@���Y�éd�ꚧ[ġR�����o鬧��NFY4������bg!^%�ޡR$}�l����Vj���k�!R���m�	�a�Q��wO�3ާ�M��"��XJOS7�d;��������+"	੹A>(�'���jZ\��R��HJ�	Q�F��%gh���r�?s>��Uʔ{TRa��n�;���֭��G�mG��#�4b��|�G� #.��r�Rj�a����X����"m}[z/L �E8�����6������g�����\a�;����(��?{o��!�h���]�}2�Ll�!�oes�f�:>�y�����A���fK,h[�C�e'Kí<P F��%�pD���n|�j�;�I�Y؇ 8F��H�w��2z԰���0�p��u㌾���.�����&�&@�F�R���-k�X$xf�
]��ƽ�I�/�h��Ha�������:� ]������&�b��T�_�?�>�4�!.����w����pR07�g�or�{�\������y�˼���r�F<v��eO��V��)9DW��r�0/�~��58Sf}��2���I�&�0�f|3���DC/�8���)g��`}��0��V��#��F���~����C�£���Fw���-��%ɉ�"U�U��5x��nX�5�ۣ��T�5�fC��!Q�A$�;����/=��\�`����#�x�(���`��#�e6����� �l�{V�:�����^U:q��7nI���ÈA]�unTv͖�fia ľ�d^���1�����n�����I��W�_&h�(����U�k�v9y9�~q2�6�
0�������:�-Lj�%Bm�4��@Z�S��_^�Y&���7{�i=��a�WHi1]� ��l�<[��e�*A�<h}$��|G�Y�I��P�,5)���pρ���ă)�T�t��r,q%:A�7����1��m0�@=wY�x�힨�=,"!��*l�R����h�ԫ��A ��qLn�_ꅃ�*g����"�Wī*S�i(�vG�fg��s��'��U�q^�BT:_���������*I`�q��o���f5�,���r�kK����aG^M�U�������^Z�_��G>̶�٩�7wG�Fc9��'d�A��W=hH�B>�g����(Ȱ��c0�#D�s������X[�!�jz��r>B�5���)��,�ݐ/�R
Ƶ>���!����P8�?���l�'��X·��
=�S��G��v��dOLFo�}]ooLd%�۸��>�)1�Ϡ�1�������j*�=E�a�_�O]��}�<[[n���,���a��^����E�q^��#@���8�A�r�iÆ�D�o����6��;�b��\j�g�W���(t��U�=��1�u�������Ff$���I�����9oH��Z60ǻ��c-S�Ik��������SV�-���fe��J�VO������zCg��0�q�S3e�9�**P����i#1�D4ѸGӸJ��ߝg+!�?��3��j�9ys&Q����X�8�����LJ�H�o�w�I��������E:�>tU� Βȴ8�Ͼ0�ޅ�8Z�ju�u�CU��mӲ���PZ[4��)T����5�t�L2�v||EȓU6��]��Y�_����w���ua-���y�8��/�X�a'��g����t-VCxg�1@�Xv0�����Z�ܥ�=J�Eh&��r:z}���j��oƀ��U���Dd�1���J4�rs�8��zB'a��;�魃�UMW�2s�W�rH��	S{+�)?+��M.��#����[$�KL������j�7o�g���$?���������l.j{덴��֎�"@��2%���A(�$�^Ok�@&�&q� ���Y�$�T���PF�Nr�̔!5-6f`���+��H4C��:+)Cd
����<�*�hi4 ��s���K���m�??�jj�I�2r!�Ь�RD7iԖ¿է�;�@D�o�
�\��Sr.kI����DZ�ƅ����qy������u�f��8d�<��n����NaHpcO_�4��f��v��o��<
ħ�Ɇ�X��s~C��F�7,�ŁT`��b{!���qՌ��T�����b����9���>F��.J�cA�=ŋ��4�^���)+f��Y�՜k���&t��DY�ӛ�����J!]��ھJ<���
h�u#�v�#�o��-64U�Q�F}��?n&\U*I]Bb�J���P_��C�-�K�~�[Z5�y�)뙼�>��|�)�y�W�������\ն�����:�W靽�����0H{�Q�Y6���hಹ��r2OTę?��O����(0]�j��ޕ���E���a�t�dR�5@+#q[(�e�p�n� ����f�W:~�GL4 
�'ϣ�I�]�rw���$"���a��J-�ȩ�X.�����7�6*�R�4Eg�A�y�q���t�p�Ia\B�WK����/��B�����|�`���L�ĵ8F�z��G�
L��!:��i�S�j�r7������\�@@���~Ռ[��3bH�����E4��!�u��)�\���MJx`�CQ{_s_������O}T��1?���e�Lw0�`ٜD��^��V��_=vڂ� ��������M�:x�Q���
W�����[7�>+X(��;bED3��s�y�t�Y㽽L�;ƀ�5K�Y��*ͲG�-����2�A�_�R���{we6̹쯦��l= w����.�����u�D$����ߘ����|P���B�i�Ӗ�`~\��ҍ&˧��X��Hbj����^�}�滈�p:��"�����Q�G{e��~x�װ���Q*���v�2T!�s���p��8rApUyH"��Ֆ2�=bk� ���,��N�v}ƚ���m�B�>���?��Z�bL��E�u��w���S�,u��N:@�ijr�P�����3�{?��S@`�6�7S���!��~|�$g'� �u]SL��u}4T�^�o��h��v�y�\��jV�'��}�qV���X�uׁk{ef������\TW�$���g�o$�ᎍ� {HyD_�1$ca��!�����K�ZL���Uɒ��ʗ���V�z�Uv�oI޲����&�9�A{�5�q����_��'��	���KH
���4��5gM�������H���m�w�<^�v��B��XcEM���y�3!����'��9���n>�io�#?�cw�\�����AҚxt�U@��Hr\2�u}.��ڢ�Wrɓc����q�b�8P��3Jy�n$��R���� ���'�vs\�bĜ�.���!���G�E'���Ƕi�� ���P���H-kFح�?JOo7-���x�٪�D~��f(Xs�(+\J�أ�" 5����6�9$���{Dv�J5����aUV�G$D�N
�q�RZi^S�Ҕ�	[���o��.��sQ����	 e�8Q����d:C�&�a��67V�)���ŧ{�qj-v��1߆A�V���P:@:��L����fB���Et�-�ސmh��S�,��lX����) l\�jwPi���Y��B���/��2�X�0ަ�h{B�C���2������~�r�V4�ٺ�]|��'���d�e�P>a���<j=��05_�i�����:�@�-<�!3>:o�79�G�Dn���Y艠���Ǚ�mv��}��C��S��l�n��c�Y�&i��p��l����m�S՛�Jj4�F�C�k���Υ�爮͢�V&z��L�����5���2R�)s��Cl�_�Ɛ\i�n��+c�ED]�W
�I����û��=����6�b4�٩|\жG0[����0� hӔ4��7 ��6����G�K?f�PF�$�yiw�Q��|�)��s`Zn�|rU�WR$M����w��T���-xb�Q�#�m��k����bYrCX��[�⡸�r���&���6�`�u�D����Rmn����|J�D�}i���@X��ο$Є��}��?�`�y׆���=�%��;��Zl$����!�1Tӂ*�`����*\�'U�����z U⯴�����lT(/���4�р�Y��2=N"wVaW�ՓkT����k�?�ّ�����h� ��s�+���銮���ƦE5ٰ+
���n\Id��j>����a/pj���9�D�*�3h����޽ﾷ��2��X�x����� X�������iB>l�_�G#A���:}]���}���[��5����[�̧��u�ϔ�3�ۤ�v���0~�U����uy;����ݍB*Q��sS���ӥ,ɫdiz���7�x˝��3)b��A@��;V�K!3�k�T�>�[��f}�����0!rW2����A�EOka�Rk%p�DT�m�pZ�t��?&̑-�~'b�y���*������Q{�%��<����~=��V#KW
�0���L���jȫ|�S�7Ż}�ӗ���N	���#�Z��6�m;C�^�tQ��p�Ev�·������e��T�<-��,aw	� o��m,'��� �Y��%(v�X��B�����	jO0��8{���ܹh�ݽ�j��u�*vE=ch�4��RJ�I�n?;jXE�
.` ����w�]���9�t��81����W� ����2���71��
�KR��B,.��R}MD����u���?-��C��Pg���ǴGؓZ��?+�w^m�Bw��#�&s?L�T��H՛ er��C�br�ғbf����xɗ>^�ԓ	�$��to���^��V�D����qk�G��J,6������Q�̋�, ��n�\g+�)�ۡ.��۸c'@�8T�~���Wo�6R�4@�K+s��@'T��m4�n�5]�K��ͅDx%B	��! ��%u���K����6.>r:����ܮ��\������t�O-�+2;
W�;%����m��s����p��������Qt��@�������Lvܚ	�-�!� ��J������b{���o�ܪ�%y�.U��W� �m	�H_¾��ñ�D$>V:d�N9ƨ�6����� ^�N��n�\}_5LJ�/�-68�r(g�̄�7 ��E�@hv^���������Q�Q'�Bu��.G]�+,��'!���-�W�U%4'�$ȓ7ٌIIP�Me������v�}��*O6d0Fcr���dq�������"`'Ԝ��7:l��Z[�qO+6_��ה��ٵ���6�.���z7�E�Ӈ�eg��~&��(C~6��e� �2�T#W�m`ǂ�3�M1�ӄV�!�W|��_�$1�9,��x7a0�N����d�B���20�p��u��qW��?����_;��+�}L�^�ڶ2���>5�_��=;����d�3��Wy���r�X�q޵R��C~"I�9�Ɋ��D�j`�Z��}�3�o�V�{����xsǿ\'٥����kg�*w�-���P֏���"o׊���-���0~��ʥ�og�N���:���<�b;;~��F`�+�Z��
�3�)��<�+�w{²>�=|a��o�h8$��x�fƛ5��wUL��[�I�X��[H٫i?) v���
�)���W~G�V,�Vk�'�E��_�Ǎ*�2&�~��h�-�u�%t��a��$h�) %�2Q8w�<����A1��@���P�-|5�����Ko�S��g��Í�ri6)葔x$���1�bq�Z0��!� @��
����<��z��f��������ͼ���c���f�q�I�Q��2Ydd�b�l���]ȌE����A;��<�q'jT��~}�X�"��σ�^Z.iX��
k��0]e��跔_7�������B5l[N�N�(�z��`p!�²1�1����l�㉹��*�+��. ���3G����0g7��,�2�F( [�(��3B4$�B�@������B��y�!��rJ�'����A����>�����<��]���EQ��kmz?Z	���J��t��U"E��&bja�g^���E��L�`�����ߗ�����\�?�g"�����HF� S N�/��;�#���$<�N����l�	�<����RU2��6@��y@T	�;-[�PU�Qn���:���$���:�[�}�	!H� �g3D͚����慨�$U�����-JS� ��/S #���1�g��\U�ע�J4�M�����LB�	9�:�{��G�|��������qX+aX�y+�r_�n8'oG�׉�6c��r�<d�R7G��4����_����x�7]M��)��_�n�1k5�J�.�ԅL�T���\t�@��S�Q�W���� �/���gF��*�.��K��K�(n#��b$J3�(���c��y �)ޑk`rWɏM��&O��A,Qy4�V����&_yߢ3{���]I��\�c��V�T��@�[�������tzqG��8Z#�M���ᗪ��d<���Ѐf�bɏևc��e�[�̳<�o?B�����a�x��0�Un�1uV�W����دxk�h�^?4z�_�N/��>Z�
5������>�YٳK���	t����{9 l�F�S;8�
Y�ټ)�]�\��۵��&��>�����R7�K	��S��a2�>���^�4&H�!NϬ���*$0�����p�:�M�]H�Y�}��J9����Z�����S5z�2c���C�]@`���Ŝ��o]�r�SƄ]�D[>\7I���I�*P�u2��6P����X@)x�)%_�gC�4;�iv�A=�:j���#��~�h�"�0im�����G����!�C��|���l:2�μ*.���}��8����﵋����6�ە�R�Yp��*4]�|p��=D�w�����$�/���F�r�}��O �?���ò�!��1#]�w`UE�0$�&.�oH�kx�:��`/�E\���d���Ey�:�c�S�XF�qhY�zEKa<f��5u���7)W/��K�U�����Q����'��$%MS��oKQ���8`$�K�}�2�f�yꏳ�,c�KkXS��:5U>b'�j�S�J �>?��3x*ѹ#���e�� J���fV=�ʰ�]���r	�j=��<��\�Bl+���_�"�$���ߴ�=?�X�a�`}����-M���z�Y	�G�hrV�˵o�ٕ��$�G��6�ïZ:oI�*�֬�7&B�Ns����o1�G���O)� ���аX��>:k����V;Ό�w�v�A����ǥ���G?IҺ�~~(�_�R&��(������6�2|�:������,��Nwe��٤��|w�'u�nB{�� �a�\��g��[���,0oW�w|3d������]�z�����̴^ Q�ͫ%~쪠\oSg��jv�ߩp�ɔ� �,2d4���{Yɰ{1*�f+j�m�kWq\h�uT����3v��T'�L����Zy��Wr�|E�#���KWrz�ߦ���й����zx��i܏�!a��\@������7�Hh�^��f>�W�.��8�����۔� 9�s�ݴ�J�L�c�/�+/]3�̠�J$z~��f#���ǭh�� �vc���mf̐�X�m~��=�t�i۟8@�&r\+n:d]i���%��k���P���0��p����@�\O5�)����8�?%ĕ�7(GNh�-W�Bߞzq�4>О�q�J�x��o=�p^ٹ�ż���C�62g����d�A��������.��cp��x�Q�}{�qd��N�fKR�U�#��;(o�XZ����X��M�g�����[%�����{��M�=���� �A=d:�	,C]�ٍ%%�I+�1 Eߧ[M��8��P�G�� 9�/�6��P�S����}y�����K|���7\m&��?�|&��3~����ט���G�����?ل腶��YC����ɼ<�����ZH����;	V�=�iN����{����xOI;)��6��sK[5ۢu��,n�[r]2J�I5�c��O�nۗ��EF��N�D�m��7��;�Y
�,�0����ވz�;5mVTY��75�/o#Ѣ]߿�B8�F�%Vn#�-�<ٽ:F���5���e6�;+�� c~�hH��m�A���� �̦G���O�ޤ6>o٤�"M�6Bh�|&�UƤ,�R�#�pf�n��&�L=���+��wgv�	��W����<���XV�`(D�KP˫�WacZ�!T�H|X!��0�{��8���e��С�������ZVa�\s���  �~���}�t���~���1������_����f��TP+��:s�"9Mz�s�?b�̓�"c��o]�j��-���"����.�e�	��e{�d��g��7@����p��4��ފ��?*|:��I��"���6���B�BM�]E�a�xP
���Wȶ���\�Z�&���Rc��4"��5�`e���vF�>y9e��س:D�%'���&hyE��a�栠��i��!�_����i�������P����ewjZ�M�qD�iXq��(pE�Cv�Ժ8R�[K$���o3tu��5k��T��4:xeS�����=���%!X8~U� �=���F�Ʒz	��}Za��)\���5	O�Y����/��"-��	y��Q/\!�8�h���^�
�h����t�{�/��A�8�s�P�f<��;7$�⇭<��
+�aq��t��1�Y�F���V��:@V���w.�㌱�l����4h�[D�/܍D���j4��d <�j�ye�R'�C7n@�򷽷A<��h��A�/M�ƫ(���v��b��F>���� E�^�A׷��Q[.�,��~M�r$B+"L{���b����	�Q�U;�����[	���?���X��F�ni�x}��h3�IҗB��|�n`@O��}��̺���:w��pwW�oc:�zN,P�1���jJ#�^I	5!��8��|,��p.���>��c���e�w��_�B<��i���^��э�	�~�㒍��x����#�$��:�uP�R$�t���?��)a��n��̼1c���|��N$���+f�u,�C�QC6��9"��!ԍ��_+}�A��ں*�coLO{Ĩ/�0̈́��1~�In�rbV0_
pX%���jx����f[k4����p���ѥhԖ:C�5ȗ[j�?	}�m���%8�+���D������^L|�;�a� e��x�nn��ﻈ���Lƹ��R|lC�5x�;c�e%r< �:����5{�6n�-E�U]դjŘ�;��Kzᯀ�7uԾ�� S(��@�q��irj�D}	�cz����_آ���lupn����O�\���%����E?1�e��gg¥D01�����݀��u��>oZ����
�
�[f�،h���b���ŉ_�T���9���">����b޳p��J��{t�1 E��w�'�b[=�G{�o� � g�h%�J���!b��I�
��;�cH6iv(#psN i�aZϸ�N���i��(}����e1�� �'˨��e�#CB���c9l6Eo7�f��yi ����~�wD���D�$ _β����Ec�b�4j��̩ޡ�E�hv�d���G�k'&'#��ݥ�c2fb���7
������R�]��R��'Ň��+/�Әݜ�/v�<")I�?�ʉ3`�����!P�iM<P��3 ����%�<q�Hg]��0��I�U�K��fH�(4�h�1�.�B�Li ���z��)i4N���~(�`���C��������3�x:�V+��l^���(O�0Xi���R�x��8�*}�6�B.ON_��\hA�l�G$C�-c�$C��z�y���#qu8p풀�VcM���{�2ǎ�m��lH^�'=�}f�yjP�шN��p5�;0Q�y�b_B�~��פ<�o�~�W�I�k����T�0��l�ΐ�k�_�Hpoc2��'��I���?��!*�!<'�FTC@!1
��˾Įoł�
�+R��X��w� ��PD����fsR:k��	@���f����W�V�<U���Cn�}�������FPzJ�"�K���i���r��M���v��}<{N0O)z�UI
�3J��J�Z��q-��u�y�[����&tQ��iE����U�,�2�!����3z��J/)��}u@�:
��cM���B1�H`ʡ�M�j�/����΄������&6��c��L�Y�Ƶ]�9k��mm�	��!�U?���vp��!�y)���z>��yI�y���1��8I��:�����>0�vmc2����c1-�	
4,���yW��Y����ԏ/{[Fl�]��A�0�j�I���%�Hz���2Ȕ�a��RX���_�Zi#z��4>��!� o�4W��G~^AF��Zm�5TsЁ����<�ر�b\7G��k;��{�5��Z`.�Nt��T|D�_i���?�YJ��O=�iR�Ź!���QMg����U�b		;���}7b���Y��_>XL!o�=��SE.`o�+Ri�5���x�$�&Dݖ�Z ���t��9�3?a�qDQ��0 ��X���i���,wR`c��Iڶo�3e����TX��[};b-��LJL��e�a��s:����&Kʁ�w�t�Za��m��'i\��E�܍jI����}��y������}˛c���c)P�R�Vʹ����%FWl0:��$VT�o��<�Pǰ�pv���_�9�L�J ��\�+���Gz�*Cc�F�q{�^=�����tꀵҸ�&	���w�`i��B�TU-k�zfPgg`ߡm�d�p���Ue	��� �F@Bb�t=.Z><;?�:�f�ÿ�.6T�G{��l�3xם�x4�!�%�,�8Z���\��둘{X�\V�ӵ�e��gP�׉)�3���K�㐩w+�ݯ�[X,�M>z�u�4��-�2O�s	Qxj�۲�E�o�����Ěx΄C6��:ɂү��#�mf���(�H:+J�屶�wa���s.���fř��7[�怇�^M���c,��#�kC��e��YWi�Dt�l$!+B�\��uG/�0,p�k��G�v�F;8�=�,頾��w^	��o8Vv���#��U�ϻn�Զ$�Ǒ���;���DT�r��l�}���1?�����b�5>c�EB4�).�oǪ(i~�Tn=���P��m=��={d���+��ս�l'8]mX��T�z��c�`���~�'p��.&훟 ��B�~o@K�K���)����߱X�E�
��R4�c�ӂ },�$ �!2��� ��Z���}�^x3���RI,9�ܣ=gX��UX6)�ST�w�b@֚*U�߾W�ҝ2j#F�8}�`]�Op#���scD��:-P��X:���2ƫz�*l%�$�NЎ{x�§�t�exYn͸��c��+�D�Wy-���k�ԌN�< ���_$��ô�q����-xs�B��m��C���x�3��萪�sU��Z���s]��� ̑G�e�A	�s�	�E�Cpωұ:��B�@��Z���w"�Tk�W_�@i��xy^'�i�s��/��|F5���}j��qRs'7�­���5#̄q$��=��A�g�d~�?�$�� ��
Hᢖ��_S��&O�����k����d�_~?�5c��G���i����f��$#L�ʿZ���]���Nr^	A��n�H�x�S�ğZ]Ǚ�wQ����Ϊ���O�Cٛ2�H�AV��o�G]��r�Ȝ��iw�~t.��pE���D4e�!I�����q]d>u6`����~��$��Y����x+Ck쉻�����7���W�Z��!�uo��J:�I��W�w�.��D����MlG;�<�ރ�,��ra/���[�:�)���t=
��Z
Q�Ǳ��(�t�:�U��st��3D>Qr��y�u/+HA��`���ϩ�$��]�ѳ4+x��͌�8��^�[��=*�U{?nF�È�v򲘸�F�$r��-�oWa��#K�3P�N��L[�)��y�'���P9�=|��sט��RP�?%��Wz��+�Kֆ�/r�O�C"B��o�jh�I�R�(ϭ.�*����(:�k�(B�+����Nn
)��8�͐s�2-�9H��y<�f�c�ȓ睧��S�vS�S��kߦ��f2�3əs�8���C��L�(��g�R��o?@c�%���l�$�E�Dh�O����;�F��q�ٟ��)� �D���w���p�!Cz������NT�ݵ�Ą��g16_�aWJ���g6RJ�Lm���2��jj�w�;@zԃ���� 	��_�z+��FW�z��1��9[��J�F;�Ơע�.;���|wRqĲ;�:^041
������%f�/�ƫ>Ej���4%��4��{h���y�u��ҍ1F��#�,�l�d� �r�z�MjX�-���s�Bsϴukz�{�����/�����3�C-�ԯ,��L����EG�f��)4�c�࣯}""�����=j�Oe�'f|�H�2$iܽz��W@��!����t������M�������-|�8q0fVjJ:Ο7�Ų,�D��mfܿk�ҧK�NW��#tR8S�;�M[Y"���wh�Ҵ���{:��g!~�2E�y�5��z�#ʠbW���φ�~g�]����vs��]gz��'
5�� P5�qr+��<��2[�"����S�J�#�h�;��d�x����=���X����(.�9sr<��\�*��C�e�}U_p�C�T�rT%�s�iS�k�<�?���sA��HzF���gˏΚ�l3l� ����d5�-�>W�ҩ?�M����v�����d��=y�iЉ!&�n�ܷ��<~�8��y-�l�V����D��:���I/N�T�Q�4���q�9C=I�����Rl�ڮ}��\�Z��]��x���o����,�ɶ�c�~�B��w5�nQ��ʛqTtŷ�'�
�T����	/�fFH�cS��n��x�� �
0ӝ`�;��b�a[��$�,G<ʇ�m)�_�ꡖH<}�_z�r�OV��|�֯�.g�ɵ����9L������TҢ��0��$�Iu&-m\jNE�\̖��we[P�.�@��³Ǯǥf�}�lxz���aM4��z�� �{�cK�_	m�a%�=hٞoi���jn|�>���#gF��VG�C��Ł�əɽƽ*}ɯ����)s��\�
��2��P� ��?��{ ��2���eje�c�f�M���O ���xaP9�Y#��͸ �D��T@����Ы4�we��җ�*�W��n�� dXYJ����9U �������.߱�4��~j�����d�哌�[���/(H��S7��	  �D�d��Z�!���,�Ɠ���=���P/.�Fd?˽�c�l?�!�2���F�,>��nDB�^�*�Qp��*>��:N�Y�Ký�Y��i���k�Zq����|���~�T���>���̮cN�Ƭ^ŷ�@oJ���θ�/t����oO[S�)I/�NnG�p�$^���\ o�~�~�F Z�s������J��:0g��k������~۠J�2�']�u|lBaK=���RU F�G/L'�RCu7�ܠjk��b�D^���ks����;���Zao�m�݋m���7�C���~S�3�Ur$����ן�h��	3��`������|�X�5�<�HA��ԍ�j�! �]����A5w��i5h������B��6���,\��ޗ�jM��3���^r]�E�����#�3�qґ��5���ӣ:Kp:�I��
�6Y�-[�ŝ=��2������đ�8l��Ѹ�5	�����)�L��[���~��I��RL<�!1zf��Uϝ�]�p�u��.]IF��,&��{%u:*5V���<���K��B�é��F��\P�L�.;.a&	'Tu�/�hZC�[s١���E�To�����f"�xE����6\�ݻUe��KR��=~^�x��e�כ�;_jxShw' Ϛ�(����o�M\�g9�A߱8���[���]���4e�R��*ԣڽ��=��c�G��{^�>��m.�z{��p���-�.y���<Ѳ5�H̚寫��&X�j�r�NQ\,�����&�T"�5b�!!Q��<r��鶠�q�����ԫ�8�I�;e���	{�nc8���0Cvŵ��?� �_�f`ɲ��@݇Xe=7��&P��m���<e{�puL6�oÿmJ�:�35]�7c"� 'fy�A��C<
��7ʉ��q���|=k�R[Q�k�DáB�Y��E�>��t�\�U[X��>xR^�o-�&�.���L'��3�K �����G���/����,�
��S?Y�~L����m3�sI��3��H��
=�QH�n�Hv��8
�VD�-o,G
�,�=������o��s�H�+>ﳝ�Ɍǉ�2WV�f���i��F� �--�&l`�qFPt7�ȈrAx�A;����zw���\m/�%�^ $�1N��Pc=��+͋�DmJ�jW����L!�w�z�Z�1�O��>�p��+B��D�ϙ�X�TM�qZ����T���=ԻJ�΁z��G73.�gZ;����?�i?i2��3`��ܣ���>n��_1�|��
�w~s����I�c�&V��;!ʞ�;���j�PQ��R�]�J�x�Oy��]�$��}T�������_1=~�Dહ�E�V�����t�'�|��m����J:+�U(c�ܝ�+.�?�s;��Yo�]�?９uΪ+˘ �Pp1�5#x^�ڦ��sx�<߁�{��t)n��Nan��kz	�"
Aĕ��P'�푻�hy�P6�$	�H>�hJ]��Z&]&�dj`)hV��1�����ɶP�w�=�\e�j��	������Aiɫ�F��ܡ�v/��O#B\B✠�7��3:���V�)����=�k�xgh�Z�E��?��,�U���]��Z�nj�8������77��� �l4��h,��rt�SR�T�M�0��c��	���Զݵ"N�ծ+t�?����.v�9������K)k�/��~�w(h���X��j{�4�Z��3��{z%�xs5�0,l��h�7�V2����%�,���;9R�J�����B2�
�����_僫��Lv��w0-��۾������b8@��B��;
���Q�T���
�Šs��_B�u� .��K�c9�kF�j��ӆ����&V�R����4��������觟k�8+L��}O?VlN��TB���$�����;<7R�G琋�=����O�/!�B?ψ��I� ����D�/��kv��#��\���r�!V�R�=J��$��9��nʝw&!z���S�k�������ERC�I,��w3��_����^�@?L�93��9~.�����h*D`��j��ۻ��y��%E���4���[�Y���L����dP��ͯkj	� 0�	s����H�� �4+�UCx{��ݨ���T6 �ph�%	)�NN�[�I��%��Йȯtx�O�)ܑH�eCX]�Z�^����K�<uR�`sa{�q�%���Z�/��L/�������Z8a�?�m+�
�k�s���\S��,ls�
��#B�p��A��ǫm}߭�X����5g�}�к�{lOl��W�N�i6��[�2���� g��.��i�G=8Iۼ>U_X��2����i��mWJb�y�7��q���L �A�hX���ʲO/'����/ɷ!�q��ѡ�������� ��\��L�z��cڨ:���I�
J�u�gZO����K� �J�u3]��S�drX�ꅜ�O����G�(�����k�0j����V>�7�����#4e�638��L�������V�e6��E
������j_�bnk15S�d��e��#�i�'e��G���R-u�o\.&�M��Ԉ���6BT��w�G~��i�A�e$�؊�u�O��	Y�Nہ�}>�ot���[�J��.�j�w��k3���F�4��+R��W�s��솸����%;e>A���� V)θ~��(��M�F�Gz@5�$	" 8疁�~\�B���Ɩ��ѴT %�Dq�8Dy_i:�H�>�s3��U�<.b�<����$Y��w�.�W	��{{�`��3]�Q��&-�C��B(�}$�Պs�����5����=&.���db�Tڗj�n�q�Q�� �\�=�A���V�$��z�C�ҋ�0o����-��J�wQp+F�i�y<�ʮ�i���a�E�*���m@�9�j������'��kw+���Q�]:�EsN��R�1L5o�����aM&Y��H4w?hAI̚z����A�����2M�s�y��<��%܉�#�\��	i.o�9�0Vڰ#/D$���M�RX9h�Gar|��a�s���V��&%��3��(E�Cb�-:^�y�6i���pj�(+�Y��6�6�_�@�@gP�ڠ��楕���tB�h�U��N�sg���q+3ae�I�+�.,'��x���YC�iu�;��TC'���� ��&�"�惇	�����+E���ޏ�����������_^@���@ 5B ũa�Ё9���rQ��j;�M{��%e�%矕����������B$kl�y�\�NfR���*[y�)OQ�}djq�ZdPV�L�_��A{�wx͇{��ݛ�G�)3���V�#�/h�w�S�a���e����, ~)��m-K{,���!:0N��w� z}�z��xA��.Ԇ��T�D�Й/d�8�bX�Q<TcԬ�Y�mV�����&�=�O�t���!���c	^x�|hPΤ(=+N��ۦ���s �P�2���.��N_��B�aA���x�>��$�z�L���~�@�QΙ��W(���uZ&����͈~r�{��.�x*y��$�Y&�;T�.����*U*�o�`G1Q���՗��L[܋��Z(���+�K@=0�^���vmp/�jZ-L��b[�4%��	�݀U~��3��{��&hˊ���0��c��0�*�	b�)nQ)ʩ�V��m��A�h_$�1m�q���cC����Y]�U�\<>�:�h�cM�F?�C�n��3�`k�oYګH�(�>�8˒���mal8��r�،�e�3qtt��ŔV�}��xeb�p݋���m1�s퍁U�D?�zCS%Shs��5�.�~ا�S��G�n�
w(i�0�{מ�e��H��Ȓ���S��pv���&q��8s{w�)�H/�T%�����{��T$�F����B;q��]f���3��y���D�梚�}�Ԣk�f�����R�Ct0A�\W��%�<�	FT�\*g����.N\Ģx��9��{�A�_Zj�QU�\��?Z(̠6@�J-�>��^DR��d �鍜`������H�Z@W�J~0)�Mjְ�+_Mq���Tj)q�ַ �3t�{�<�E������}�c�VY�T�Kcu�5���;%~�\�U�4 ���q���U.�Kg�l�O�%�N]�rg��6қo�»��ה_�W���D�곲��oe՟H�7���O ��m=:�Wf�RV�'��b���rR�o�?��� ��^���'bf��L��礂h����4���S��?���.P�\2�3�c�n-�+�!,��=�<���
E��Io�0��f`\q{����8�۷�)�߶hq�*z��;A��-[�MY&Ɔ�|s]+��UE�ڂ%*�~{F�.&���5w��5$��G�4�Y���	�?�Y�^7a���6FVFb��(Ef��8r3�ʽp?���2��;�9�&ș-oΆ:0��nu�]�����ښ�{�;O]���8�2��$�W��N
�d�E�/�~��'�wOp3�!���>b��Jz(b�Fs���.��L4�=S'�3��D��/מ�����'���t�o$��$��l?�ר� ��Wt0oC���3��&尯���ɥY7\,��4�	ͥ�ҁ�2�p�/�JVaKJ�����wg����m�f��uR���5y �J��)%�By���왑v���q���-4���^��*V����(p�����j���%�ѭ7�P���@��6�XDP-ي��}ʐ���WR��/�3�ñ�4Al�����J�-���2�(I�)g`���B�����4�q��
@UE�OY�/)#�-�V8�D�z���A�UDU��j�3P�	|�vk�,�b<���ƛ��IT������|2���m#w�&����R�N9�(��e̪N㲐G��$�*UЫ��-#j�1)�Ǘ�Z��ӈ��d�����,
2o�f��u��FZ�~y'��w>5��������ԩ��IX�i�
��'ީ;k@�9٬0n����}��7�X���{Gx����t^;b��؋��&N��c7Z���-{�U������IA��{�����s���m�|�J�@�����k6!w�Jˁ��B]M:L�D����MQ�[p Ĵ2�uY�߈v��*��	S�B�0�p�.�����Ͱ�Y��.����I��9�-�GT��|#�>6?��ޮF�>�ץ�����u�'d,PL[B�������\c��K�2*��䇿����g2ә�G�
ڳ��:=�p�"�+���) m�R25[����F�C�M@j��ق�^�50�I>��Z� {Σؿ�����̉���)���ʢI�k
�cMC��g���]$��E+��b�V[\�d��eck}�B=�y�S�`�P#F$g
$Z�V�Sb�F����}d�⎴���7���������nF��cd��K]��fO������j���P,�l-�!��[��򧘥I�m<is���g!���+��Bȧ��Y�>�!�6f�	�{ڰ��^�:�e[&��~���U����:��]+<kkVk�h
ܰ �d_�/����8\����tT=]໒L|	y��N��}�R�����4)-Y�A����]�ut��>�	������ne�
!���n�?R�p)d7w<HZDݑ;�z%��z����>�8�Q���$a���(.�LڦqE 3�a��H.@q�%5wk=��q���9z�i?��8���hO�1�����
{����
ǒrŒO�}YtX%��I�X3�5E˨������p�!��rk���JS��=���1)�9�S��6Tim�*)�1�9�CI��3}0��16Pn�	*�a�ܣ����܀��8���`%��J^o.ۄJ2��Itj2`&��&��˦��ݜ\�h��	W�:V�W<Rl.\���3����E)�BD�;�6aa_$�D2���7ϋ;��q���ءHi�N)�~��oۦ׆!eݫ4Q�plB9�O.��cn��peU7:8��^��n,3�B񄃑��e;�-���Sx��Ip���%u\)��kh�B�V��	��?�d��� �Է�ךEa�����"?��W�q�<$ӈ �!�S�Z���I�QK9��l7z�&6�2�)���������(n@���
�I3���<j�a�=��cTqT{�a�?��8�]���k��#� 죒w����q����C ëED������'��>|@!GZZ&B=%����z+�2��E�����n�M1�=|�͓��7��
��Ng|":{���$�n����O_T�ƭ��Nd5#�w^#�K~gu ��TY50�Q��0�g5zV�h$y��zR�/���E�|.0���m!p���8�x
��7_r�&hH*�~T͓�$� |��B��)#%�l�«�p�f�>��?Wd�4)�ٖS����;��hda[����sQ��pV7w�(��0G�!�p�=��NwK�2nz�9/�he�S�j�K3W�3�������wx%��F��Ы'���[M���@�S��CW�|/s֚5�D/7��>~Xݘʊ-��6���������dc`�ц�>�t9c*DZ�wH{�M ��%�9%�Ö� 8_��ȩ���&�E�i��j��tơ��9����]�O�Һ��u����;+C.�{���&�M�t�T�)^Щ��lx�AH��B�d�<�p*��;�C�|�&���a4t8��woΠ���I@[�,�#�@�f0
�(͏��M������ +y������C#�u�����n�}*�Vj��5���R�g���̜�jX �ڍS});}����*�ܬ W�(�����d�A�N������+�*����ހ�����p��#��
䤽��cC��ؓEAd`���Č�b��vC@l�oFX�8EtB��{���� �+1zq�1WK-�pZU�a��sc��� �F��$!�,�2Ƭ���(>x��@�1c�P�l�G� �r?�e��T����q��ls��e����p~���tmRQ�c�fS�)�z.<���|
�4[
��c�c6P���Cb�^�q�7Ŭ7L� ])�;9UBu�����XH��-�ƭ	xRv��4��B��΃D5#�v��0������	VYM�S!�ý?sv'��ì���??��p�)�1�b�'
���f�&��������p5����=C�^L��}gS�J^�շ�Q��}�r��/r����m#TP	P�PL�
��Ea��s$YQ��[h;̀�j.:2�o�"xWX�08�!�����w�;�`{�U�j��fRu�Z/�$0oF�y1shrG��@�q�ܣ�0������:m����� ��fRs����ױ\�F�,��@�c��Q)_���b����^c7�y4H: ���lg��u"�Du���v�Ȳ�KIgeU���f�^~d�!��<1�-՟m��[�My#|�*H�`��;�Lb�)ަ
Z��(bPr{7�l��*���"3U�F�6�9w�K�CQ���A��s�ш�T��G!غA<@�[fwJ'D\B����	��4���Sr�t�˰޸C/vD/�@��O� ����U�	�K��3�휍TU���X�o\��2+����6�c&�`�G�Y�Kz�`n�eJBRQOf"�so	�
�ߊ�.�B��5��O�qn�i6
� ��]��0�k!8ѧ�muHk8����?T�-�Tu�`���3�DZ��x���}�3�SV[e-<�7֞�Z��D�H׿+
�	{���V-��/�!�pi�Q����?��7��b� (�x,�#-�9�ᠱ�:��ќ=]Qaz���M���T�u?;��RX>�v����������^�ӂ�ڃ��;���y�"J�G�a*���l�>Nߑ�Hw���;���\:#�ݭ�j�h�{��xTl˜m#�<��W��_�|� w����'%��r����5h�9������Ak�<�hڟ21I���p_�`-��_�
`n�?�%�wQU	�������=��4]� ����"���)eظ9t���g�@�E���V�}�A�ݛ�[��=#a�F��20��FF!��谊7(S��v��\
A�ȫl����a� ��J��8w��odRc%T��ҧ��v�4�PB��z��d��!3��(V�bs���N�1�D��O�p?eX�|�S��A�-w���c���h��Z8U(�E��-��+�tB��s3��A��eA^�џ���~�%f�?�t�b��m�6-���6\����̐F�-�밹}�=�K�/�Q�L��;����z�)��R�ֽ�{u�5�6�4��������j�עa͐�ɦ�����K�Ho�L��v3H�8����b(�{�om�d�1�+z���?R���R%[���i2��M�:�B-}g���%�9��b��&T6��!�����ʅ��}i:�u�4+$o���\`G(�`Y-���#�/��X���uZ�_ccDet*��p�I윆�8 "�#� M�11|�E�"��Z�W}�=�p	 	0">�Φ)8���C�*
�?f=Q�T(y���� ۆ�ҭ���f��F�i�V���:�|�>�(�k��E-LI���	l����{nym��)Js�����Y
#����!��ɉ��y�w�(-���ܚ�kuEZ\�V��S彖3R�r�Df�p����Md8V����58c��4X�ٳZ�G_`P��z�� Yc��� 6L���g��;� Y� ��Ϸ���0D@y�?!��g��I��t�oa��|�VeQ�w8�f����t�g����%�@���K��ӱ�A1e�;Na���Y1�p!���B��-����/�W���sm�HX
b������	��G.�S5B������W��A-<S��G*� �q7��ܬ<���60i~U��"��P�4�);�:U�������?��9Ў�sF�U8$��&<�ȫ�#{5U�JbOdA�����,����b�*&��J_�[B�C?�`s�z���p���̷X�T�th_Z$�	���+%�x2�W��4T�B��\w�òz�=���1�p��[��a�ܨ3x̃�����D�J��brz\Xx
���4���ϳ���Ƞ]j�k�;{B{��e���R�X�I����&N :�:7IS1g��W�A�Q �<@�Ǌ����W;��T"^�����̒|��k�;��$���� (����-8lɑ 1BH��1~�?��/͏��|�
����.���Eɭ..��5a�CK9ԡ��G�i�S��_k�H��EG�QD�F�x�qp�Я���J1A�Cɧ��m{�d�~(o�tW<�Ja-�C*���ڏ$�"=���1c��	�k��-ky�3��AñJlDo��$i��C���qo�bΡJ�	L���W��C�����E�$�ɿk�xi|� i�.��>6�d���0����>���F�{�r脖?�?Ҋ���^��yG+�㻸i�c�����Nqp�{K����`�!��/���`���5����	3�1+�0U�<YJYƟ.yw�9���D��y
��-!�N�[�V
���D��3�.˃�~ǵ�7�Ns������R~�%������$��鷨A=��459(It�N��|��&��_�\���9�X�)�Cz@"*A���񸲗'��w:����)�����	����gã���sT$�7���(g�l� ��ٞK��USDz�����RR�{�{d4��yc%�P�V�Y��/[��F+t��n��%�R��KӉ���ߐ���2��g:��ggQq�H;_�P��J����,�_�z�,�XA�1]+�:*�"<�KO^�z��x=o}���+�N���'
��r���a@����}:-:ɝ�S���a�qЦ$�Zy�ݗү9a~EZ��đ��%>S��S;9���+�^AYu�u�7��[J�Z������t��􋌑>��>�X�唓��H�Z��&3O���r�쁩R�\t�qO:�4	��8<��>�=�ګ�R�,H�b_ybQ�#�۞��cn�/��'�i��Q�I(��FKSR�D��ut��v�ve�y)�>v�w�CLC �\9eE�V�O [��0���)$��h��V0��ޠy�X6_I���X�{�k��N�$�LVC-
uz���{>�$�
�OC�
�*U�;�E�:�W�	�g��jaHH6��,]�_��4j"E|��@���)@>L��S&�ZX�Ȇ���@���O��2���uL�E��V9Y,vV��[����+��i�.D����ҫ�p"ʞ#����Ȍ�I��i_X��ЄN����Ox8s&�Ae^����f�@Q�V�]]R8!��ah��/�U�8Z^���U;���vn Q��gA@�)��>��e�u������|-���k-�����$�Zt�P����,�͸��� *2jps�*v��1�#MCo�ؗ�� KV�F,]x���`�}�������m��d*-W<=ū	�/���\HuX]%����g�ih�?nBL>d��ё��{����a��O;d\��b��k��e0���L�/�V�|�-[Q/�o�ZvuQ�+�໢���������e�-[*���E��&��ŉ �X>��II��x�h�;�W��GT̋ϯn�^J\'F�7��՝�T���:�y1D�� J�
Y�Þ�@����8�H��|<��szˬ?�ᦎ�B����*.\���Ȥ}8bŝ1�,�V#�ch� ɑh*Қ�ݔ�;х�?�``&i��Ds*��Ix/j�UD��t�.��/k�&�>�nG`��~�0����*��_n3��v���/�I-#N���~����8hFY��V�[{k�C0�̽�Ԡ�~��>��܊'�B����3� ���)�Z�*���x+��>}�|�U��(��w�����u���H��H]�L���v}B�.BI'RH�&Yп,=�������3a
`��M��郣�A��u��3Ag����il�C����$�;��g��6�n9?.^��:&�,`h�D��@�aln�hcD�
B}|> ���*���a���� ���g��D����s�b[�?X��|fb�IE�4��p�4e�֖0�ҕ�m��j��v�#,������;����R6r�^�a:^�NP��ZI좔�ȥ�_k�	|H#��m.��������F�=�d��	��7G2ҭ&.Z�c�u�ߗ���Ū�[v�R9[+^6M�ʚG��+��C��Q�k�ڝ�?qO# ����oUχ�t��̸�O ��e�1�с-�'n ���%@�7)J7�������h�&�<�Gh�0H�$/�Z�#�;I,���!c1��=�pd�a��Ʋڷ� �¶aR���據h+�Z�S� �_�Lc���wP�(i�1uj��ӔG@7ӗ�IhٛCܩ�k~�*Wt�+�7��y�]:�2�\oL�-M�nr](s�$=80t��J����1�3�;�@�oH�z+29�Ʊ�80�^��t��FB0ŀ'�N>��PPz��R��i+ќxQ���*�i]�DX�N?��:�� �:E^�?���_:ޣ\�� e��=po�7����:Y�3Vc�r)�����}6�7�$ˮT;�:��:��ɑ��ڴ��峭(]y��/�+�<�#�Ky���?`.���̘��髺�|���>+m>���Ee��V"sA��E���q�m� �S�׾�ڲ��׹&����;@e�N���Z��Xָ�>�@�ycvU�[Q�o���3�Lǻ��T���l$��y��_9r� (��T����KG�=��%!��~���.�P�{t�����tmeM�.mvb���& �o@5Eq���w�&�k���t�<+��`����{�����]-nh&�Ų�m��f:�u�8����Me�r��-"1�-�u�s��27U/�dw��;���vj�� Z���q)�����q�H *���� �#��QD�+�\+��?NHHd7�!)�[�ٺt���!'��
��'e��)H����ȃJ�k�s��!�����ܷ���G�a�)>C�-Wc`���-)4�:�/�0�~�b"f���Yi#I�*��n%�d�c��>��0����0�I�����4]��e����ЋX����)�fw<��^�N���@&?�ޣ��^> ?Q
G\?n[�-l4�'�
o��q�Y.ѱ�F�����?��mݫ���6�J�4��ְru�+,=w��~A-�w�qlr=���Ċ;�L\�B��/xG.{.��W��4o%�T�h�
�3*f�Z��=�Yl	D�Ø���K�j����]]$��fFݍb'�U�mC�FW#�',���_i�ӹ���Inz�y�g��D�3�UO�~�^_H���U9W@},@�!]9����D�Bo�<��(�7��?Ǎ�����9����ڌ��Я�")��F�Aڂ �.yzL#���.*4_>5�X��2��t�Vci)$�uR���}��T�Ʈk��=���b�Գ�����w$�Qr)�)�3�,|�V�@�������v�{f�]�d������4<�,hڽ��f��nyS��88����RY�a �Q�.b���R�c䋤�l~ivCa�?p�֮\��s�X�^�/Dm%�;����|��I���]�y--c�`g�l�&�ֈ0�c��TP�~�IO���H�Ī���#邙m��H�ͰW��p�H���(�a��5k-ϝ������15��L��1h�b)]Ȩ�>m�� �����Q1��k�o���Y
�Lb�=�Pj�4V��v�C����!}o����2˕p���a��~��)#t�,i�]ċ��MU3a�w���?U����\,��Z��4��A�Q��c�2��y�'? G� cY�=t٣/��,�y��A,o�
����5�_�J����C21�Y�f��eac0�	���V�޶V�K��!�����LcdԨx���y�I��9���)�{V���g(��;&��*��m9�R'�GI#$+��q���xwn
�֔�]f������&&M�21cI�����B���/��_��;�@�dת*������q{�3�d"(E�������c��"ܑ�4�*lǦS�ތ��hk8ޚ������gHU�!$�ZH������$p�� E)�qE)o<���嶯��N��j �n0S�h�$9c���J�&�G	�'��I��{RPb	�ʫ"��*�i��Ԝ}C���$�n�����ጦ!�!A�ac�JV,�z��	�2Ny�ʒp��JӘ(|}�Qdů� �:�ILX:���4��\K��?�D�+�f���K斊�o!�ן=\OL�$e�g�'D�49�x6N{ݿ�v��;�M��1O
���h�w5` �h����z�&XW�V���m�@��SJ���x�
���竬�i�h	� ~P�C��|%_�����	�۝	�*��vY�}Jt��ڣQB��jB��� g�^+��7:����б�D/�#�5�֞�N�h����|�+�j'GA��d���>�m�h�b�ۜ�0���օ���+���E%�׾��
� �i�;�RCZK��^K��7
�&��`-�R���G(e�R�����݄��k�����Pp��2?>�)�,Ml��a[(-�O�x=4���e!;���k�@���b��׫�M5�xm�E�}=�\��~!%�����7K�;��Ӕ=�o�蝝��MB��.�Ab��7x$�|��.)��Υ*.S���Ip<��D@����q�!B�K �O��sg���g�j�����~6�"��Ä!����U��AJOZ>6�~'A��[�<�HkaB#2�N��{%���d�FɃ��rߋ��f���G�����۹E|�o?��A�%�Pf#K���_N�	ۚ�}D�'b��\��1%�Q�f��pDn؄3������~DL�:+�>�X�����IͣSIIf��8%�����:�o>���(֥��-O�*�'A��������;T�i�p���]��85k� �g�u�Ŷ�M!N}�5yVgz\�!~_�ih+�q��}�z@{Pu�ɀ�6���
���W�բ�3P}�>��}Ǒ�/�RAd�D���1>Fxh;���Y�04��:A���߶/G̎�j���A}q�cx\��G0��X �,�n�_igĦo��b�&,$)CK�j�fʻ[���~֕2Q:4���hlph�4ӵ�lPֺrK|�M��t��CB���L��S-��-V��25d�J�����q��yԤ��Q��'=���I�%B���mH.^<���z��鍿���M��l<��[���D��p��,<�G�b|oMs-��(;�O�z2�!��~:�.��z_����@�����𐶲x6�DI<+��(1bRqN�?�wY�����9f��i��~¢�L��	�)��7�U���uy������g^����b-d� O�#_��&w���ʏ"XŃC�Cf���@��&6R̈��1 _�Q��F�����/�1�YP���"?M�{q+��o�3]�,�ͫ��4~�
�c|�j�N����{z+J_f[O�}bI]��)#2�:�d��I���g��]������,�9	"�>MM����iOG�t�cnU�B5L��lR%�*��d���ivZj1�yQb��=��&�P�q���ڠ�}�d���NW��F���n� �Q13w���Be�U_k��#��q?�V9@fAAz7��Lv�c p�&~��쟪�CAsj�Vׁ���l3s�KB�������y9t��<P�F��^�,�"�[�PL?tp�@�k
���o�O���5^�G�߹4CB;O{�E��Sr�L���q&�����I�eMKaWC5�C��Y 5q��^��YD���噲��}�%����FVǨ!v"rp����/'�2�����Y�[��]o��%��!�\Q��`fi�|{�Z�G(�DJ ��D�{����O��h	sLb7$@Oc�����p �P֯4�n�B��_U`�"k��'�\��;"9'���cޜ�U�U�8�o_xFt��k�y����4��k�k;f'ľa[��?�d�!� (���]�%��Z��'5>|���J�
�~���� ͒%>*��t�8�z}+��2pŎ�h�|{)�/���:��7�>!����P`��רv�J�a�;\ �v�#AL�F�\������#���y��z:z��)g�YSf�F�*O���k������׆�N���yH�ʡ.�R>�ф�-|���C����y���֌i��}h�DPƓi&��m��n�.�^}n������pP�~
��l�������hf�.dke���Oe�j�eW��hp��,��@��Bn���/o�]�`թ�%�N��R�x���Th�_��0�; ��S��M?$��mH��U9IQ���x��G�ﶜ76�C�{���c!���
0��Ժ��.ݠ���>r{�w#�����plۗaVXț���3�O�P��rs(w������}�!��6-gB/��ȾP�Q�Q��)V�WM�at_
�t>Љ�۽�2t0c0��NO�~�yK�1>'
M}b3���R�d�2�h�ȓ[�)�0ݦtd�?�H�>h�qH9Q.:�]�N8�N7�[�-�9���P�f��ark�e�z�e�h�H݈C��|PŘsBq�Sh�n��z���n�8t�?�L�~Z]]�Zi�^�iǟ֟5~�������u,V������~�M��$4�q����<�N��/>y�/G���j{����Uh顂dӿe"�5��T�LW��_]���n0f�"Io�/	�켯�Ve~��Qx���|�w�@�"[���A�)��Q��	��<����v��6�x��/A{��`����a�F���|��C�^�ݏ\(��&�)L���W�a���X��^�~���������ͫ8ĝ�3.i������_=o��Jd�5�3����8��u�A�^������Z�5������z
���a��?Z�czŘ�������FC��B����lsK�5���"1��t�d�C�G�\[���3[��_'�~qM]50{%�8�Ƙ� fg�p��*%z6Ԡ��d�Ћ(�$Y�H�ٲ�߼�q,�(s�{@ܚm�j�ab7�]t1��
+8��c�_�����Dz ��i��^�Z�>��uġ:n���Im�ph5��������Z��ӞZ��G�"T��]�^�3r�i!jM����?R�9<��l
�s��,0���w�L�HA�X�Ɖ5o�7�'�(B�KMz8�t�����<pVs�Zr1���,��d�Ԇ5>�\:��Qy	����&�k8�bUb�Z��[PP@N�
֌KM9;C��h1��׳*�E)����牨9U��1���g~�X�ݝ4���D���b�PgLT����bhd����|׫�
7G��l�,��%��ގJtc��u$�y,;���Y�n ��n�{�M����S%�ԻcWm���	�{Ƙ�/g�,X���:�Q]���#�.�{�p�t�n�I��Bo���jV��KA�����G}�I��}���ߛd�,Y+���Q�s�d�c��/��o��Xo����_~5�~���yr�>��U�E�,�����!��� M㗯����u�E���޺Zw=�h�/ھ.���2(9ؽ��pN�L����a��G�kec#<%�9"�X�dN��͊����N�|����D��X31�@�!�C�>��Ӫ~G��^�E�S-���[�	*�'����5�D*&��3KH$��i�@��@L�}�_��N��8v_*L?�WD�Y�q��
�ݶ��0��]�j5[��7�n�K[�sd���4:�&���0�1�T��A`$�)�m5�<�Ů�COc�K�/�%	�Ma���2�����֛�q9��P����<������P����l��Z�W�j憧��{Ir�hߢY���}��'���_��sd���NxY�D�i��f�c���⪅G��ohC��6�GUa��Ϙ������'̷�{����J����L��KV����ݒ�LT�EaR-p"F~J)�u����H*F?:�������׀���޼�Q*�RS�y�LxĨ�(���hd�_��U0k��o<���ެ-aS���ÿ�b/�@�z��*i��h�%4(YkLA
$ω1;1 ��i�O�	��(?�X��,�d3�v�Cԟ ��ݘ>#��1���L:LT ��?����Tf�sk����B0�5�~��C��`��ׁ%�;dC���I��po+�WfWA�p��E��r�<��׏�$
@U<���]&Q˾
�Dp�X |e�[b=:�&����ӧ�q,�$�q����>6Z'T��w�6G� |�G
,��ct�%M�"ۛ�7�-A�Լ�g��x�m���=N������o��U�֙�@\�l�Du�&w�ck@
�֌�#�K���
M��^"Fr��WX�3:Uf�|��(6��%������m{���s[q{�&�Y;����m�I�N��e#{��IK�F�d@��d��§9��El�Gnϊ�s���ﱮ����&�&s�6	�����-�vI;m�5ZH@5ޥC�͛���\���CSB�����X�	FR�BY�����ѱ
�рv,����K��n�ǽ�JBѶ:Dq*���4���8xE��Q�a|Q��Re��]R�*d�D����
�72M7�!lW�FQ4;RS��dqq[k�zf�鈄���8��{��8y��mՁ*����`�ŗ��O[���[G���ϓ�&�`~��#���2��z��s��{�"m�\w��<?��N�s�@^Yr�1�Θ�����Z`�����.����t�S�gĺ	�"jw�Qn�۟�6�Vj��x�~�M�l�tqeu��@Nl�Sb�ͭD���_�>���>^�4Зe7�����M�L�*w p]}���$c���y<�"P�1,�krJ�j���M!�$��I7U�hl��ިs�� ��*�9|͞*�E�D��(��L�n4�ڪʖp-�|�c&-���h�����n�g�_h��%�y�ޜr �b���'  ��Da]�3ngp�
a��)k����8g|�3��%>�T��T��'r���C�@]�s����_��,LSeq�F�ww\���;��;�}�~SC]���=L��������0�W��I�}�T�b�y�Bb���}A`���`l�b�7'���|t��j�¤A����1��z�-@��L���m��}� +�Nr�o�&��'f6�V��ʫB��՟�uL�>펁4��'����Q4�a2[��$ؗ{��Nd���k��k�
^&%�d(O���N2$��v�A�rг�qk~[@q�ϖ������3U���@���N�����j�יz;�mF�e���!Q�Xȵ���Wb7�v�A|�-�[Ɔ
�cU�R�,�M��\Y����^:����2/߈J���.�����&��	��TԗX>"$���ͪ���E��s+���jLF�z@��6�7h	�г��)z_H}��f�{�o�lQPv�*1�t��i^��j��g���/�ۂz$�K�+a��ʗ���&�� Zi�R9��fu�������5���/
��D�P�^�W!G1+��q�T9�u��p�\��*���gˡ�=��ի��_=��qN��������>oX�e��M��1� <��d]W����b1"�L<��\�O��Z�t���E�4��ݴ.]C�#̜�Q�gr��B4�0A��aͫ2�n��ϐgQp��^l#��TL)�?��^�����tX�[����K2��^�`�����M���+�j	Ņ�@�W�ܷyg�hOI�|����c`�k�R�ӃމBK�!*��֭�J�a��%���d����K����$	���:��vΞ�y鍼?Hu�rI�L����� �4�p'{����}��P�NV����>�jcS�W�I9}�'01�o�0�w@�#B��q^N�}�1)�ٟ�Ru�m}Y�}�1u�;�Z���fW;s��{��w��~a�$��� 'b	�8x�+��h�.��Gv�S���~M��|[�7j���w��J�W�=A���Q�ql`՘�����6�*�U��<�H�JY���v}��Q�[�D����R��6Kf+��XB�j:d7RS
���*�`Ke�#ށ0ش*�}����@������ԃ�x�R�;�W�^����@�L��h��4�ی����q���1���������y��>�$���?�>�br���bW��Yߑ8�t�O�m��w��`T��& �U�|G.�_!O��D��M0�%v�v7k�B��5���G��ϲ��`��>��t�8(�p��`[��G)<�/K�$�CŌ�L�z���S
BL�2Sڍ�'>9�,3 ������i�l��x���+�f������,�v�qCf=ҟY�[M����O^$K���h���ˏ����{�x��I��2kYq����}�d&ҷ�[j=>����o������M���G�+��3�vMW��fҽj�su��~�\�W�R)��P|��L�{b[�P�ﴜ��5�.~�WtΥz~�R���L�BQ��D����ܵ�iN�=�}(�լ �x��V���'Ը]ߩ�q3!!�/.�,#h���^�M<+�?s��֜.��=��w���,Z�����R�䫒�VC]KN�^D�Q��N���X��;�|��p|��@��cq}�·������8�/8P��M~���(+������)ԷO��Lͳe�ގ�?-pwH�!�]mh�����#�d���W s��}ƅyw
�y4eD�+�M	��v��~���=�[wz�|:�l�:b�����!�D�f��ɒ"��MS^,�Ζ���D�H��.r�@��\�wQT/�7ȴ�U��$�FYS3�v��'t��|���ϵ�H[�5��M#9��b&B^�s����G"�=���9�{`}w�3�"y��?��>���!C�\�Huc��=���At���"j�j6�hn�NwKE�?a�����W��,
p�[��
f6�-���@^z;R0����ū�Y��1\����Y8z�\�/`��O.6d�t��X{�4�yt+7��'i8�#�JV�^Y�il7lG{�魩�{�-���/;���&N"I21B @e7�S���I�t�q��H�:���C���bp��u�<_W�F���)(4gaF��8���"W���v��	�p��NL���D�7��?�^L�^q��U�-X����}�Q|_�$�/xz���{ŖLolR�G
^�&��>�2/X��W�.kS�y���:aF���A=0��O���p�(`�|�y�����gZ��A�W!���2u�ִj��>�C[7�D|�B�Ѿ�9P�����G�Oh$Ì�N�=5R�Y�����)�|�R�e�Y�vf�8>J5�a�7�ڜ5� z{k��kZ��'*<P�+ɑPR�hU������*Z�_2�:|�;ɂ��  ��hm�о�����+99��䅞L�-<U�c��Ch��s/�V9ҫ4G�)�ـ�t6��!i�i����y'��ۣ�ս��9[��vJ�=�?;�L��7�'�/������V��5���A��a�(@���]RШ�`�N��ll#����e����X!"�M�y���k�=#��/1u�~��L�|���--�j����ē����5RG&��&Qk���9u�+q��/@6��bSF�=)�6�d�^	�xC>�D[�B�ë�\�&D�P���sb��"�B��q�"k�棹�|���Rq�ԈW2J~j��K�3Mܳ�hi����2Q(��z��B�]���b�c<�3&���2뜴�7�'��r�C�b��ە�3&[fbs7�Y:۪+,X����4h0������%-�
���\���L�0��z��jD�}��<N.�T���W�L�nR�O)&E�$HY��O�2�h�.�cne�A�L�U�˝<i����x̖,��>�j�?eGP���$�}��)'����}0P���s~��qþ��"�@"7v~ۙ  D��}�������m2��,�K<�lvy�|��#�Iӡ]M�1�q��2���8��!W����p��9(:z[�޻�χ0y;샻��6-��@DS*$���-BhnO##Qעj&>���8�V�w۔Gd�a���,9k�3���M�߈��w-3�K@��k��G�䤪s��m��U�����7e��A�ҳ=���[�wSy�ew��Zm~�(�e����e+5΀e:�Q�bk��D���nٟ����1�����4\�4�A�mq�/��xyܖ=�~���a� <�/D��T>:o���UU�c��Ðb�a�18155�ѱj���7����3�>�{��U]κ��~�Z��t� d�K�m
'�U��c��V�"��J)MNHLm������z`m�UR���w	M-�Y��|W�%���̺��b��N���������?�yZ)2�km; O��� 7�oVI&h�)`5���U?/Rŏ��ȉ�S�=:����W��Z��1�Z̠p�@}���?S��h0��E�q�gL���§�?�fe�VbQО�0h��R��� H��_��a$_Rހ������;K�|��d-��ԫMK�$����l�9�-Fȏ�Hź�r��B��w�����Lq��fL`�SjHWS��a�{�L��R���:���-����u�f�|.�3i���_N�{\�h�@�%_�D�[���^�2���Q��nkk��0vN�ߦ��l9�}��/�`vi@���H �T�7M����qZEguNhqZ��F]�SC����9'E"���U����@�9��u^�Ȉ��t���G�8�lp�����y�烲�"��+4Q�6Bc��� 
��Q?󧈏3{3-�|�!���.�0N�W#Ƙ�d��Բq���@e��I�^Nx�(\�u�x�^ލ&���y��W` 3a*�����x��8N@����	��i%?"F���ܴ��R���L��M��-�462���=���K���M�h~B(�Y�[�u!T�[Ћ����U�D�@Ng�~Y�f����0Lh%�ZV�]v)��Mni�F�o��!i'ő88Cg�{�v�������pf��1v����ʯ 7j�QVm���@3������sX�_u�m�x!y%�L������X�p�9^7|~�O�o�ua��Y���~��T�(����:c,���"�*`��3D�L�%�4Y���&���ɡ7��G��ܑ�17�Z���q�͝��JK?�?��𜿟���0���.$d׵����w�4�
���ķ�21!U��.�.�|o�P��3~�����\�
تo9����X]p�6Yz�Gh+�=�"W�8Y{�u ���i�.-���i�g#���K�-�F�O*���T����@2(an
I��q�f\|��TJ0ޜ�y�����l�K�-�o}b�E�yQ����mP@%��'Ȃ�D�c}��}c(��w ��qfҳн+j�!M���l���f$�)1��C%�y�&dvj_���c��NK"��L��6�r�-�6�f�_�y'!ۥ���,n�qsLt^���R�ͭa�&Г.'�������0���S%˙Ela+�`��p����Ϩq��Rc�9�����M��i���<h��Jm�O��|a���S�1!7�`�h6TlDj��eHhh�|����d,oO$ �ؑ:��/P�;EL���L�@�?��a�$)�y����ў̛�7ϱ�i��2���l�J\U���aĽ�yÜ��y����h��pm8g�UJ('^��W�E�>#��4���|#��1B�p�B��#�뽌U��ӿO؁3����[���^4��A>��K�γ��XzĒHK�j���������J#�WX.n_T�Ue�~X�_��X�̨�&I2�{sƓ��5��?� �eU�Iw `O��,;ɻ���������~�҆s(�hk�Ow��cH��eK.��쨫h�	kðM�WR�;�<���!���M��hQ�Ž��1�����L�G�0�:'����^C͌2:���'��Κ8�獨��r�o�E'k������o���*�x9V��dAY��y��D�8�wF�l���u�h�~*f̩,zX睲���W]Fvoc!�6c} B��/�	�1Bp�$�����m��`�ڮ���j7��Lym�zA#������vSe�`-z���u�9���A��0�`hÂ[}o�uV�ޓى����/�x�IZo�L<=<r
�/���D�,>�~Ã��3�v{�'H���0�<�I\�MS�Q���C�%뙕�Jx��lt!�_�= �_άapHm*��k�i���@꟰�U�򅶅jiɴ����K�VM�(r�z;���z��}��'Iꙝ�]�P:�L�@��o� �1D��gK<���֊݀�o~�X���%���D����*�E7�LtOzđ#�k]������tfKMa��:��˘��p��#�y5��n<gl����*v.C�vu����,F3$z�N�E��E����`�H� e^��1u�������{x=� OZ-�Sj���e�"]���\В4�ʓ�*\dӡ���5��m���hژ>���8#@IyՉ���)��icuI��F�i�_�!��a��'n�O.>L�3���U��ὖĨ��{\�buGM=���S���O�1!���$D�7���Lu=,��,����v��ˌ�6����l�������tVXC�G�F�&CE�a��0���$q��E����A�#�}_
�u�啣�ل��$��)�{��|ѤJ��1��e�
܎,�1�&�N@��~)r�`��?�V�n�ɻ�K�ʌ8��+�q�v�ac�2g&��c�d�I٧��I���K��k��O��{�!/�/λ��B����T1}�*Ⱐh���x�����Myu����3��Zx���Z0��«���J�<�����]p�ތ���:�ثZ4�d��Վ�͙Ǧ������A�g�Z�>G�n�(�BF���W�����?���Yc�zk�'�Wꕋ��ۨV��d>��8�4
O,z�%k�|��4���������j3�7�?�T"H����+��bi���mY剬��0�k}7WJ����
��Q�K0"�[b��.�$����_9�X9hf����,��|��w�e��0
]�q�ɗ�J+D�A`�]��m�V`4�5�j��.�J�hX}�HW�O�	L��a
IZi4�gN>���{e�3[�&3?�mw�aМ��J�Q[Ȃ�M�?�s��.DP���O�D�e��K��sݼZ�$CnjN�e��������� �N�k46�
λ2��Փ�v�e��h,�z'�e&���'��KE� !�͑z�`�>)��;f��s}��h���a��#�a�R!�8�~?�l(1ݒ�K���5s�]�<�4l� �P�#�q��%-H1�wYfR�&��ީCkq�Ղ^a�I��2�)���֊�֘����%�&�>�OPW�b�(�E�=�L����q�3�;�k���yU��qx�7 L��[�~��~����\���b=�T@�qp��ci*�2�
��zM�1g�zxm�����
�).��o�/*��S�+�c�q�V��BG�"����G�#O�jI�I������Y>Y�U��KG�����v�E�Mu�)"��y��|��v���݂?����;B����� ������7��m�{!��M�w��uk�u쯹����fF�:�1��@@ou5����c�Jre�)M��N ��'������7��@�+�b��g�d�0���LW o3�g��m]-]���9
��7QThF�<�sʸ�LPj=s�<V�kJ����9��H�e�`�}���l���'��4s *�.� Z����u�һ
�r<K�g7�X#��%�X�p���{3���� Q�py �����R�ަKU�%)�q�Kxr��{ �Ha3��3Ivp�fՁ8H�EMp��r�3��Yl>zXTY=]Ek��R�n�_����
�4Ec2e�ޢ� �i�P����p�����^���C���\ B8��S�t��Rg�>���X�|�W���u;�|�j�oL���΢L�9C�m�ej�#m���G�0>_#�� o�L��8���faR%�b��}L�/w����~�T��UB���<<W8�C��K�(���Z���B"�()s���T��3�ᘗ���O��JJ)�V`(��pN��-,T�X���w����ٯ	���G�Z�=���~�i��S]y�RVʒ�M'��&V�0D9���9�`6I�K4���kaY l�>>`��A�٭���Z+�4�?x� ��n_5�1xrM�G�`^�I�.C��7�g������+Y�Ё�+	y���l�<��+d�!��D{'����h7}��Ҁ|�U@����"W��W�8�P��F�ߏ(��g��c'=�}>
F�������͸����A�?Ի�u����^���]����c�8���o_-I�V�O���b6Y���/�wu�6.��{�)nܴ��$���;z�����x����\tl_�ރ�
�-���6w�ŉ&=�<�
�}}v�ο�������_��,�W�S����N�S�j�U�޾�; *"

w���ӱ,?w(�i!�?u4�Fڙ�2��V�������0P�JN�������`����x��Z�u�?"�/�
P�6���:@i,y;P0�"Tx�V9]TF�%��um9A3�]Y(��Xs���r����O&`�R��L�2�:��e�"7	�'k���Bu�2�nj�+,�������D��k�w�������ؤ�5�d���^�<��H#a����y�Ĵ��Ɔ�q�vHq���������������^��Љ���y%݄<|V��T(��T��âc
�BX���=(�ݚi��r�|?}�2\�n&� ����'bsmq;5����U��w�!�+Sq��.3W�Zq�b���BVdW��<�^\ۦmvC���ŽRo���O�6ˮ�K�:���x�o�늚8Z�E��o����A�Ew[����t�쐖��_�w��1��qrt+�瑆׏�#N5��������^�DZ-� <�pFn`��lI������U婸�DwEV?���iֳ�2�YE4x�<]Oy���>�{�5����|#�nx���*�HG��d�wL���6�F,%�ߗC�1!�w���O����� �Zkr��Wv�f�{>�\�e�ʹ�~��\��W�ab�ȸ��Ю���r8�3��E�6
�� �^�tdX�H?U��C�f�#��E�3��O��e����/[3���jW{Ʀ�D18�.Ӱ�:�&7:M%��G�PG���a}�pz���u[':���>��B`Ԁn(n�ק,X�*֔��ڥ�b-��?r��z�WdN��o�r-��<�o�k�(��\��B}�Od����),��~�#B�`��uc8:'a�kQa��<JJ�]�����'Iq��\��I�
w@<&�w��g�TDȷ�_r�I��s��v_���3/R%|>���߫���&���2A����<��U�|�?F�p݇juc�{��}���{��q�y�%O��lm���(�y��&s��2�~	�7�gELY�J�F���~��W�Q�{�e�����u��,�[>�t�4�t$����n(�*��&�g��r.��=G��˺�� �(�b|=�@�ۑ���p���7�`���Bԩ�� �� �}ͼ�ۼ��N���(&O����s6o�t�nB�9��7���m'�/���v�������`n�{x�pzC$v⺙��i]�49,h��Hn'К�z�'73Vf��4y�u'ʊ��>��'Z��̫� s?�4�x$epZ��a���*��_g��剳����L�߲~|����|��&��I��Qh�_0��QJ
G��m�"�M�E����xP~Xe~H(����e�"uv(��t�|^����?��|�)��3�h�!����W���9��+��0b.��<Z��^�ޖ���{� 5=ĵ �K�?�U|��>���e��=���!C�g=�����[�7�Tkݽ���n�Lcu'�J��G0g�s��5��I�^1$%������ɍ��}�c3�����(^BrJ.{x�����ѡ�>�S'�t�>���m�舶���_�����=kϲ����n���,�~YI�' uoj�wM�zl�oZ�	� ���D2�.T�؄�Mܼ[�'c�}���-��78}�Y{}�o���"XIn
����輏+ޱ�=�+�Fj�v��<������6�f�}��Q�,a>Z�$��lqLƁ�֝k7��G���m�a��s�^�̍����t\l%�w!�B)6/2}:_/<��5.D2k�F��R2����A̮�,�}_l�m7Z���G�:#/��*֍�b���yMh�(��Z�)�F��{$�;@@�F��E�N骫��"��SvˠFӭ�쐍�]-�� �!�i�U���-�Ѕ�s�u�b٢{��]�)�1�^�ڴM.	:o�v�@H�?�/��@~&�p�y8}��ґ�o���d3��^O��KN"b��D��V=)�ӝ������!H݉�k��J�3�ljV��/�Q>EE~��I�e x1�!y� �W��s<T�Y�����h�yMP/��=���.�p,��Z�,bZKcW�E���}c��rL̆�ן\�����W
��]�k���z�B����J%6�TaNՋW��:=�x�j'O��A u}Jf?}@!��yP�8,x2n��_�d�{��$�����wq����Ù�1��]dS�x�n��1$�/��5qh-&��)��4[����CX�Ʈ��0�""���߱�[���|l��6��l3AP�@7vG"�?#x"�^�H���:�w|_Z5�H����G�j!� 4���d��0����V�?*��<|W�.��{�����c[<9�����Д�F-h�7Ƨ����3t�&]`>�7X���eP�Eu��Tu0��W�p�Gɘ7Kn�.���z)uq�Z>�n\�"�_�>�'NB�j�<�5����)���p>{_�����e�^ ��jw�	}&�5�� ��c7=�����������W�7�	:����*Ed����d���t'Ek_��߽�xN���aM>2�n��h� bZ�c��k�ɲ��2t����I?�Pۓ�?�#�z׌B���^�<���5m�T(�sp�$0�h��Ӧ�V}""	1�À�Z�q�81o��I
9V9�����e�]���EPg.˱�L	��w���]�] vZ�{"��.(�����`7C2�έ{!�t$J30Ƀ���6�H� ����r�D�����0,X+k��h��F��9H�V]�-�Dm�B|�eA�q���ݴ�����+&���В4��\?\�/q�2&���r @��8A�j�BLh�g��	�B&�6��h���RY.�x�C\-����2<�e�dB^�˸7�u�H���,^8Y砨Jg�k��1�V���&�X�)~3*�7����|���D������w����9�F���W��_��GN�[f��%"����:��i�2�}
O����nsGqlء)�>�m�J[q�3m)ѓ����+n�O��i!�v��/F�2 ���+@q�`�G	�1G�*�6a�����1ྯ�Ė�zV:��X3u��-�ญy��1_j��2�\I��Ծ>��H}� �b�M��ܠ�
�rX`!�,-͊�a*g��d�(5߁c��X7;Ie'WU�:~T�È���͸�ġ��3x��ԩA.�+���3��X;�L|t�A���Ғ�E<6�����;�Z �q�V�+������<`����r��;ڨ�ƣ}�(U�B�j\�?����A���e }�H"2��p�$mɥ�	IXN�<���
N�Pk��pGo@��<��X#A��+�����~��Gz���{z���\ͤ�JSwI�݋i`��8 ���TS_�z��Գ�@��i������9
֛)�=ד����7�����RT&������2�j']�|5Ł���3�wEb�q{���P�ɝ��v+��U�8\`C�m�ϒ��]�ȑV�����7e��Rg�`ĸ0�p�ݤ�ꡃ~yP(v�&��#f`�ؗb�ib��@���5	8�U
�j=L�Z ��a��]z�!'�_Ǖ��C2f)>|O\�n��]Xe�X��������*k.^e~3��].����
�S�!*v\�����pir1�4��nq��Zo�{�џ�K���d�T;�@-�1�� ��R�yj,�M�� ��e���N�[��ӖQ�៉z�O�F&>(��Y���9!GH,&JB̅Ek�ݐ�E�}�ý	~֗�g"�&u��6zmX�P�[��6B�uClZUȶx7�	� ��A�E*h��Z��ª�d�9`7�9���xr�� k���ڋ�k��&�j�2.���+u�Xj�;��*�:Ud�w�~ߗ��Ƒ���Hɾ���Fw��a����݀�eW�R���%9>r3Y����]�D�|