��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2f����"w� �Iv}�aa�*�c1̫'$�qCiD�������A���6�'��['����Oh*`� iKx֍036�b��Z4�V��r��Kz p��cH�?L�s΂���Ad͔�\4$ �墍ZS�q��@D�����QdM��Ä�����m�-z���o����}*�ڴd�dd�bf���� �Ȇ-���Uj ���#����D=�P��"<��\+ki�S��A%�Z������*�JT�Mc��/P���˶�,Yʡ�8 �)��.G3?e{z0�z�U��s|�ƭ�Z���{��J��sNy�-K_�(wWh!r�zܧ^��������ʉ�w�ac���/*�u	>R�P��C��h@S���p�U���5V�B��1i̚��C��TrQ���w��֣�2���.`�X������;K���@���.g2N*M��+(;뮘���u�fuZ�\�]���[�"��G��5�>{ncǫ�p[MJt@LQD��4(bQpR<�%CN16�Ac��Iu��6��E���b���P�w�h���!F��~>�D�i�I<���[R{�S��1�v��r��jf����+S�T?w�`h3��+ƕBEH��L�"-<>!�HKZ�1S�N,�(��.�5�qi��嗓(�n����g����d�a��_��N��� �'�7�bP��f��xP~�&�mvz]JjM�:}1�I�0��)_S"u��ۉ�X��,������D,�}1M�e�]8}e����j��9�(��?�{�v��1��&QfL��G���L$��Q�`S����y�w���
��07�ӂS���05)������M��Uw��� �j��N�dц̍F(���}��w40��-%�=���}���f���~��8WBLЩ��z���d��bͦw��P�R={qj��27��FB��I؄T�p���+&�5���J>Ka�
�&�P�,*�r__�_�,����/���_m;`�͟@�U�;B�y*`�O��X�cݐ�S��Nq��G�_jh(���t5�|a�3�0�~p����E/�~���؇b瀬�'#���GG�TJK�/�{u�)���f�_���/ǟ�C�/3
��c��)s�~�:Xe���X��4x(�K�5[����I0���5c�!g�x���,W��Wy'����r�#��vz��Im�D���8b�'!7L���5�5��=}h�+ڸ;� ��;�P�����aN6�Sqӈ#/Zع	;�+��#"�{�P�ї�G���0�⽵:�K�E���0��Ma �k�q�t�Ε[���A�a6Ї�ܖ=���@v#k�&=wS�S���4�*P�12��^q�ކ��3��m�:�"n�%���xF�KT^b�>� ��!�~0Ц���!Z���%�H�'�G��*WCf�y�g���`U���uV����Haw�JgR5�j�A�ݬ�J��E��/K���N�b�E�qp��]jّ�7ш5@����ݙ[,^���'y#�	��5���j�KX�u�ӻK�QG
x�%���8�+� �MG��L�M;�4iah��L�sW�ֵ��/~}��D_�� �*���՞B�o������t���A����8w�G/(��_��s����e�s2����A��z���C\������T�`N�
/����3�r>�@tND��]ެ�*א��S�|7Qk[��4Kt;���!��ڱ�Ԝ�}Ϟ��59[,� ���ӕ�k��Ʈ|!�<	����"���'��5�N�tVJ��K�Q�QsG�P��~WE8Zz���Q�FCY������n��=��� ��:
��,��y2$d�i�gj���P	[p;{��3��Юa������'��l��9�K1_<�]}��ʾ�q���s���k���Pf���&t��$�O����<ɹ��)*'�m���߶���]%�\�\#��J�����{^CѦ,U���o�.dt�qV��tkR��ݠ+5/����ݳO�w��������+��^�Q��? <o	UvѩTm�[�q1����A^��]cV���D���/f��z��#����m�$o�ˁ��@aCٲ)�G���L2�+�?����,P�h�����u�|�>(�ɥ5}h$�׃S#���i�D�X�9����i��ڼ�v���?�w`"��Z�������+7G��>�X�;��%-��C_����H>-����F)�m���p�S�"�2I�d�����7H�i��g����ǣ��.z�B �'�<�ޫX9��<�4=��@�����f�>T��y�(�72�K��A_�8���B5�v2���%���rj�߻�=w�N���Q��"�N�Xf��FQ�����@���/��-��t���� )�:U�w��.5(��I��&Mb�w`	ZXGX;��9#B`;~}�tX�|��?wN�׀����3á3��O=3�&����c#�G���l�Yg:e1a��9��gaA*���}�Z!�!��~�IJ��H��v0�[����1�*c�J۬$D�Q�DF���`��\��'m��Rm���[SF[��?��g��h��_U%
R����b�46orU#��,J��M�9�o |`�1&��߱�ߠ�x��j���E�U�V��E�{�}��	:�y_�<BE��´�0�����vf�*���2+S�o��G@�U1K�V��:�)���T����cNUNh��߷��������(��>����?�;Y��C+a��U�V�S���D[*�cMjGMZ�����J<H�QG���HMO��"��Ҋ��@��iq��۱!X|�nZp�#���&e��3u�26=�ˁ m#֬�����:<~`H
�/#�>,7�A�����HuP�'�đ2������a�K=��1�&�v^�>�.;6��Y@!~�7�\������!`�G��hp�uv�9��O���\�p����UDĤ���|�|��C`�`�'>�V֣�WO8�@p��n��O<�k��~F �o!�n�[A�`y��
�m�a�T���m�J����L�1
��[�w�9t�q�Mvr?Uc��T\�eU�U�$���}ĮW�$3��(u,���d0�s���ifz��l��o�S7��S�'Id���3	�����YA�o����Y��$@��aY���� ����a�m�G>%P�z�������Y�j3q*�r��lـĸ�vH[?v��Q�R���c�$���ek�i?S��4٭�_�X�^��Q6��q׀�����ĊX��b>3��F��fs9z�e��7�b���U�JKRǙ0X���4P(:�\�Ng���9�C}4���WC�r��&�18�>�v�S���^"��?�ĴK�ѽ�k]����.l����e�O�SJ�`����n�ʜ����8��Ƌd�i�o=�<�������<<-(-u̾Pލ�?��>���a=N��MC$w�uʄ�*���}�������r=޷_��l�,nم�4����(��R�l >}��O�興ӶƂ��F��
[]k-VW���5t"�]��!`ͦ��?�=Lt9���}�e��!Mm��E<t�22hS�fqNn��̘�©������7���8���.��Ț�j�7Z#��(��ϺZ�4m)[�q��˜
�堝� ��#�����ϒ�Lh���T$��. �ԡI���/d
���H��P�i���¾�@7l���a,}3Q��z�P�����Ɨ�m.�n���L)<��/Ap��>!��0ϥ�_$G�Q/����غY�U�,N;6
�
�e�Q·P��铲��
⾸U��|7��̣b�k
��F�E�O6�����*ؾ��	��"�]�"x�9w����S5I�%?�M�&�k$N �"�p��>�r1V�2PUp�5��wj�c����t5&H$ Y݆,�\��`	L��^��Q�Q�L�A5���8ɦ᫉Nz��ہd���-;��{�D��[�>k
c`u������ɛ����;���I��׊�Tv�z&�*9D�W�L,1�NM��a�(ڟ��F�*?�F֫.d�0/�
�
@����_7��ž��>�
�tꌠkf����5m��� �M�&�D�!!]��EQ_�8�uc����G��P�U��"��!����K7�7}���P��H��%��g��t&�P^:d��Wz=�M�j�/� �}����i>Z95O���{L�����U�����x���m'_"#)#��E\�V���M�E`�5�nl��%iD�w݇��.ofws��,}Z�����
"|��,�๟�������ʋ�ػU�?��u�L��$CZ<A/+<��=<	߫�������e�NN�%�K��fN�R�v�	6�h��I�2]h<�� ��x�0�||�M�~xrL���K�E�:�h����;k��A�c�Q5�.�k�D8U�x��T�)|�3$^7"�E���JM)zH�l��q�g�����*�8
�	]�Da�^Jw�⧸�ش�7��m1��'t�4�m&8�f�/7\��p=��H��J�B���)u5+"#b/�?�}u@�˓��8��ڹ�`6�����rs�D�������)ls+H�lR�i�2��� P;	[�qT7�uF��������~�������!V_�bC��K�]�ޖ�Z[���T�\-T<"l?P#\�0�X:J�,�]2�s5<�Sk-7C��w']���U���|�1�i6��c������"��0��H��r�-�`�\;��U@��~���u.5}!!I��}tzg)�Y�|�r�Zy��|�_���E���	��S�HX�-��:��.a���S�QlM��t�週���,*	�ۋ(��A��} ��AR�?�~Ɏ�'ǚ�M
�k�RHN��D���Y�W0;���4�>��� ��h��[L��b�79�Z��|�4����U�tz��I(w�1z{�<R�����K`�d�R�ʠ���"�h�XOAy�s�b ���b�sh�l�s���ѳ�w���#W����k�Ea�̠b$ΓE��#��=/�
\��<dՇx�L6��os#GZQB%���9��)���D2bX���Ju:�w�5jMB9ب>�7ܯC�&���tq��C�
d��x��g�߱P��HA�-�.roe�[�H�ƀ*	XZ�,̰��	l�֔:��AIt��k�k@^�ŮՖ�F��>֨��ջ��6ǿ���0�c��>���W�l�ΰ�|���i=%{��inX���R'5T%{i��n=�%l6ɏ@J�?/�8�}6�����n�����K�b|J!�����\�JV~;��6�o��pӧ�X���,��&(�[��Bc^���1m��b�Ҥ�GdɑR#�[i��Hp���0�����9x���!v��}sk���@�EL��t��ƴp�}�/q�4(��S�Iw� ��.�L؃�}���r�Z��|��i2��r�C�*�իE��d�|F�at�J��@o���F�M��L�  H�F(N�����߹��u�i� �~�6��k�!`a4JG{�p�=vVBd��c�q���� V��>:�<�%�b���)9t�J�c�W�Iy��7Tmv�),�2�V$w���a;�R97�u�-��;�����SmD˨��]W'uE�VH�9��i�=�f#�b��%�ĵ@�ȷ��J|�i�b�'/����n����O*�v����D`���E8�uXv����� |jf��g���N�v���&�Cv�T�
Lbd�:r������$�g o�Ᶎw촲L��_!x��).Iĵr�E�y����4�A澒��*�?Z`(�M5é�-<~[e6�4k竡0Wy6�J��22��h�x�����A��r��DQ�Z�؇�J�����xi��{����B>h
���ի�O�0�_�p�]G	��J��dp�Y	�)+��뤹���/īc���`�Y��Tv�������5��n�
\�.
�$�D_�d�Y�Un�=�gu��M��<�?������j:��d�7p#H"iP�%~���+,X��;��+7p�j�H�-Lk(�`�V=ǝ��"J_`��"�1���n�P��r��@��8�ŏ9�� ��@i��-v@���;ۦ}�!��/�Xɠ*��O�z�y�#�"�+ʫ$���˱z�f�)g�D���m��P
2���l��s;�Q�y��_���ȏd���v�	��Cw�K�Ais�I����З���V����+?O���6zj�龴�d�m��ʉ��x뺷Mft��>��I�GJI�[P�+�
�� �`F8�&�@d�(
8~��w�s���	��L�����jY����K SN�=�?��V� ���q�oa�����> Fc#�vҷ����f�([�"q!��"���iʿ��g���w��'i�U��E�+f���E���H���((u8bhq�>��ֿ�C��V��/���UB�V������I?��縏���#skQV!��5�ޢ܃����,ɡuY�*D��ͼQ��Zk�{�fk����D���.f�J���N�6v��"k�(g��s�EH�]]M��h}s�CbT�"T�'xls�����J�p�����},C�>& Q:�ɩM�
�g���o),�X�R��b��&Ee�{<4��+�:�&��*��,m���f`l��"���-�׉��=n�"�I�l�%��`��?�+�ߵX�q���>c10Pm���h������OhJ�g��3��9 �+�5��Hh{�j67��=��;�(MLS��x�%��"�x�Q���B�V��ۍkp��;���]�&�.'�4��i�4�����?��T��I�h��9W>8�]wp��՗_\L���ПAO$��{t�b��fb(}��+��ټ/��G��=�p�aI��7G�ɘ[2���]E.�'��=�#��V�V��9Bm���z֎zZ&���;���K��N.W����Y�D&[��"��K���y/u����dO�C5��8���QbcI_�~�?ʱ�(��b	l/�j�����5iq�7	��"�>-�pk�U�m��,,Mw6>�QơO�N9�H8b+�2C���F�]Y���C��?K*f��Q��Ad��Ah�\���-r��C�{yc�@j�հ^����t/���]�G�?Psf��{���'�D�-Q���&\s�$�������T�dA�3ZGO�7���Pf�AO�TY���I&SB@ӽ4�(z�!�Gl%Pgˇ��`�N���=M��U{ը`�i��֜?�5o]�Is�'6�S�s��ZwqS_W�����>�����GTML[�d��a����R!$��Q�Ѧ�K S��{]�~~2s4��x'�"�����S��H�����j,Ŀ97�[���C���}����]�ύ���t���-�ՠFR��d�=<�"d|:�ձ9��z5x��&�Q8��k�6�ty��C�N�T���ʺ!\(]=?��y���|��h�
����{V�����l�;[n �@-�����})w����5�����iJW\!��V�!V&#��;�Ę
}�j��Y!�����6���v򖣅��e���$��a J�O�4)��)x%�H�lH	�4r��YJ.�x����˂�v6tv��ZS�ʒg&Oņu���/<>�/ճ��O�"��c�o7�&L��Ḿ����>���_����$G��b8�W���p:pl��5KY�6��9Y�F���}��"r��f7��N�+��Ҥ��|Y�J�=�(�m��Iq{D^A��mg7��*]1�?�X�g���7N0� 7i�Hv[����HR�2�5Cbÿ�
$Y�N��\�D�76 "z5C�(-�Bm��[�����2j͢����ez�+dP��
tz7/�����2���S@y���n���-/=b>}&>�ە�*�W���7�'��@k����JӐ�-���=��Y4�x@ �ʾ�W��5>VNW��d5F�����dV8du�?�OM{��n��>�*�w"���,�o�� �ZQ�ɶJ���S����B�5���mA:2���e�� `3�<W�\��U�	
���T�Ֆ-Pr��p.�x���m�)����^��/Z�VX3�l�s�H��wD����n%K���@��*+� ��z���.i.��
�|K7���V�k�k���ni$P�ཾjVNy�'4Eihbc:e�7��u��T�e+�Q������AH�"f�8�QᾆAϸ��+kh��eZ��ٶ��vwG�v��GBD�$S׮8x緊Y�Wi]���=T �`�lB��/�g�X����N��3	WA�P�\��mS����<��c��A_C���ҕ�H�&՚�2����b�\�����i1�^b�۹HkQ*ˏ�3�@��5RU�HS�6+��'���w�i��e�����.r?�m�V�Ȁu��l�+ ���r�!oJ���ށJj@��X(�~I�
�+a�|t���Ş'���k���R߷��Gݎ� c�J``)"9������sD��1��p�gc���n�G�o�C�<�ٌ���`r�գ�-�/�k�i&���4ѷ�8-9*�S�R�u����^e�w&/�)��%�6G<���c?��@]�?���
����-o���c	�Ch�铣4��|ܐ���v�p��.;u{sI��w6�_߫���d��Ի��#nLKL�;��-��q�����$رҐ��2zE��!n��c���f^>�0Pz���7�g����2 躣��w���.�(�m	�*�a����]��̇?�I�c=Yͺ��?>r�1X�o�t�ߩ�3���5�#mq}>��1���X l��>��]d����[w�y9�sQ�I�#�)f4�n>bFe�M�Ղ�}�Z�Ce�8/��S�=T
8�LC��E�V�D���m��L�!f���:��4�X��.��&�V^n�J�
��t^\և������j��Ro1�v� d �hE����@h�I�4�H�4"D'���!�bH,�� �~�$�_�Ԉc���f�����~���έD%rH��nm��x&�A�v��b�A�oJ�#u���ً�z�
r0����p��>;NE��p__��m�����wȥ	��p��CG7�B�0AT�1Q)�q���@�Q�e�o�43��
`�U�4�5Ztt���YX��w��O�F�bi.R��p:�jeX�����O�f�NӘœ2o��gr��x�E]�c"�X}j2>F�a4RBȃD���� �m��"�A��f<1Oh�ڃ�J53۵{������|BC���}D�*B	=W�94�2X�{�����)���4zk�Hݺ�*aD������fT�-w�P?D��[V����!���`l��K�2������k*����&��ܺ��i7�`6��W��ù/m����2�\hT���M�d��C�E@�@\m�4�a�`Xrt�f(���>aV��+�;�����.��$lT���c���mLЫ���`�oѦB�g5M�3Y��V� �1��?{��ξz/^Rlg�*4��6J��W���J�6n��Ö��XUt.����q��>��j������.4��}+BFw7n�»��q7�ui�J�8�2KK�1�[_!�t
�G�t�P4ud	�
�����d�O��cS��봽--@�,�v����\�Gj�Ij�@5����uw��8���K��S�1tI���L4��
k����X_�4v��י�"� �J������E���������%"�p�F��g��Ӌl2D�r���a�M���9<���,��k<>$2��.�n����moe3m� �DAw!6�ʌ�Yͼ��I���Q��F%ΐh%\WO�Y�@;+P�~��'wE�]��_�]��{�w��}x�)����ǃ��G�3���+���I��Ԣ4��"Ҹ��;T��t��7���ڦP���5�X�v%����;������j�]���RvG-f�%ħi EЂW6�^Ђ`��,�Ԉy����I���8<{t�2I��Γ���x��+Q�8��m���OwR?�4�<�&�}�j<���������Q�L��%���N�6��p�C�1!�E(q��ǵ�TJN�P��$2΁$\tsՅ|x��]O��c�� T	Fc&!#(bZ����pC�S�$z;f^zGG���ӀqG��-[�f`04���T���]U�oLv)9y�({��Od���5�%-Z�eQqv���4�=�=�1ߜ�0;��Y�֖?H���:b���1���b��������!4+*o��u�<&T�C������;�Kp��W
l8�`��jn!,�� N�Ue�)7�W[�uM�1�ї����ns8�U�����/H�;�k�ļ�WD��E�]&z(�Y���~�����E�U�Q�	�a+u��r1���<��$>��k�xs��Gk��?l�Z�]U��N��Z=g�wٳ=`��S%�c�x�G��E�κ�E���#Hu��'���NƵC�
��:�lፏ�Q�]�u����v̨��D�nK8w��Iv�&����5�t�*�.�B��П��l�O�K05�?��ܾM���O�u;�S�ѝ�<�=<�c�R������'w���Nr����bX�	0GL��j�*�����^�&T|g+/Q��@���>���s�G�`��x-�z�|V2�	,���^N�}��5&�^36�y�9���֛����>��8�d�#�f��+Q_v?y{(�7� _�$]�[w�h�w�U�ٽ %}"I�� ��b�=��k�w��C�4	h�u��j^_�	�H�m��F�(A�e`����/-��k#tG�UE�I��[&Z{V����P��F[�*͞��z&�+��iڏW�y!�E�b�_��ɨ،�g�������� J��}��q���e�F����h�!7���ŏY�B]^��>�!�'��W��۹�L���`�=�'��
={�a�Qs��$�Ҥ�̶�ʄ�O���r�O!�5o�e�d��n�o��BE�9u{k���(|O�Qps�<l^��^����ݞ��qIء._�hr8���-ޥ#u���v52׹j��hLҘ�F��M ��ئ2��E2����)ۺ��T���(k�S��(�:<%&^*���v0x(��/���&95g���A�f��j�A�K���=�����1�5����G cm{�eZ��ݛD���H�iG��`��cS-| l����ȟ���V_&� [�̺�!��v��;?u��T�2yZ[Ec��|Q������.��C;�m�ۋ���cwʺ��oc�oL�O�ϗ����.���)�]��y�t���hʏ@=
��2ب+�AJ˗���	��ww���_^�g<��vn*},ֱ��h�|�%��c�{����	?&��A�$"Y �����a�	�~�<�m���F�Ղͩ�ڎ�u�w�Ywv`^ؕ�