��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?Bk��nߨ\���	--�2%��mB'~̰�����0�ƛk�w��G<ij��M#Ȥ�]�Z�Q�iF9�)P�}⃒�e�\��rgH����$�Aw�.����9�U�ANH�@��4K}����!��IV�jqIo
#��nL���Tv�!��勈(yW�����*�n17V��O��B�_�U��`�ŘE��*�Be�P�I�P�:g����G}���X�˒�M����%:Q�g��m�K��$MXE)�j5X����	�۔P:~��I&1�`����h�z���Ps7���Ct�L�9^#�öRh/$J:�4/D���K�m�,��6c��娗ݪF�����f��Q����g�xYD��N� �h�k*��\����٠�K��9
�Ͻ�ܙ�08Շ/.j؀��t���[:����f�Ez��S��Y�%��L��enF��zؤ��iM(¤C�T�̟G�H�h;=�8�<F��6�a>lŃ˸>�N؞����^��eǑ<�N�rL?����YVF\9`Ѡo����e������$�gr�B�����fP9�-�Hzڿ����Ǭ� ��ҌÈMWYN�L�+#��	у���a :
���30l~zZ?
`4-Bzz����
��tF<l�ъ��8�����KX�i9�������e��S�|���+K1��X�|g1�� ������!9�-_�ײ��˓��xZb�O����(��R�A�o�~�{z-�$8봻������0�9���0;��]��M-_�G+���zF�7�E��~� � ��P!��:�;�J�� x�M @z��<ʠ�{�\D�b]����<?⵹?u�pkm�w�r����L�Q�2�ۏ���,k/��?�� N��7�E� �T[�o�����M��r�B�h��fnm4���Gdm�	�Fz��j��YÓ��?�����$�Mhk�M�i������7��?��0��}[\���5̛nL���l��Ve;~X��O0۠��m���~���儃���s�;�]���Ӧ��Z�S�'-[3��yё���2�rx��<���		��-z��mk�u������K�#���׾X�s�P�-�z��!Òs��������6����5J/�.��(���@���HI<B=�2U��q�}8�E���$�e�;�/��vC�Ǖ*���A(?�����G��AU?��e�2�&l�W��HO���;���G1���if!���o'%@#��l6K�VH+X�!���u�9���X�C=X-l���0�����ѠL��pZ=��Ļ�N[��.qˌ�E$�m�G�XI��}q+RYW�[Q�V[�N4ja��H���q��
C�����E�3߯F/�����`�U>*w3���FU��A8��E�7���O��<l����<�I��l��O:�[�4@h�,��f>�V&�23�)R`)x�7�H��,��H{~����[����挠%���B!+2�/��&JUn���0���%�����1�ٕY̠
|����~'�B�9b�m�=�VP��m��o�����d�JF_m2��z8�-��^��$4���g��d=��?�A%�b���	���|w�
��҅����vr���������H�*��W���E�4�ʥ�2�~;�2\|U�'ǟ���'�����_eƴu����qßJ��)�����mV�-�A����4A�)R,d��A�Ǚ'��w\��s���T�p�j	F�H'vn
�`��z䠆O%�;��A1Qy{�n/���M�VAH_b���V��'bȵ�h0��~��#���aZ6 �jE�⎪��\���E�!�ܓ��"b�K
I�X!�1Q�Zv�cj����?��m#7^��IϢ����o7M��0ƕ�Ifjn
��Ŗ�۶b+��F�3�uq�\�ƒ:���γ�뮕b,>H�������_Y;��	n�1	fԘh6}#��_��bY>��k����2�0�2q��m��m���4_��Dg�e�i_d5����R�~Hn�A��M<�,Qָw���Х�z=�FIٞR��G���D8��>���.؅Fc���&GmEⓦr����{HtV<����0��Q��iMZ\�p�Bp��q�-�#�䗷hd��1�)�>]��Ef�X�8�j�;q)� �wM����D`�p��m�5�/���`"ʑܤ�M�J'�6�W�^��R,]�[Xc`�[���&}��2��'�W��Z|"��i�z&�R�O���['�#D}4&���nX±Oe:O�:�"Frlt��P����Xp3��_��u�+�w�5��E�R�~Ys;4v�W]r -���X����Y&DFta:������Ky�c�Z���Ny���@��6���7�J��t'G�.��oT����s���T
Q1�T�B���[3};,���ޗu���IOs�p��5/,��V1�t�][��ʏ�u��m���%G&��F����͹���~E�S�����;���0'��"9�;�O��IJK8�#�Cڄ#o��=)��xy���$�t��n��X�뜏�Ƞ�Ğ�N��2x�ww��((m�8(G�*Ϝ�Lxk����E�Of����i��^I�"��s�a�ـ��n
T��d����Pvݦ����W	�H�R �������㋏��w|E�1_���7����Y�3�#�V��m&�,cr�ty�J�ә�3���7'oPe�G^5��2�VO����,@�0"����;:R\X�~�Jp(�L�HE�cvH $��ѯ2���������|�p�"�P<�c�^ǒpZ2J���YA)	��֎���Ŝ��7���'�C��[&BE�8�X-���qqR�Kx�3n�0��h& TR>���dH�t��F�`���]sg���B1�z,�"Z)M�}�P۔��U��(/�.��ei�}���$��|��-Ʌo��-n���te�P:��>b�Pρ#p�9&d�0྆�r�1�b@���bl��3�nS|�°��'��+={����M�� ��/��hG̷���+���� ��+�����WC�o8pNi_����Z�g���_F�Ο���Av��zl/P������n��J��`��?���θ�pA��ݑ@>"��H�:*g���jrI��r�.rO���4��Y`x�����xt���1?Ȑ����`��f��
�fzF�I�\zY�\�G���'h�����c�E
F�Ԧ��h�¶�D���f��&���%��}Q.����rV�+�C�v�K�xO�}Ѳ,�a�F|a�#�I�B�W��>7)N/;�D���6Z�*�&K�V%��+K�( #o�[�N�R˦�2�9�����A��7Q�-�G��_+�w��c�6d�k�f����u�Ȋ���oV� ei}Lm��d�P�>�^�v[����4<G)BK*��A�s{F��8(�I}*�3�eQδd��*E
:���@���ߦ4:J��o�{AF-1a>����Uv���Q
�&_�o4Y��S4�@��d`��r!~�ᅖ���1�@� ��ט�� �	c{�Q�iXGS��,O�cj�"�'SfQ�������4��p�4�wi���4h���7Pj�ִSs5�6mpGƄ������q�ԯ<�%s��{Ϩ���A8�C$IY�1�.���6e����|��'&&�{���r��9fr�E����#��VV	�����x���F�#����R+�H�j���1�߳�9���7(�K\t8g�q� *�.�?&uT$���"�Q���������Ϸ�{�yJ�DB��0�����y���d�h,�ࣻ�#�&��Eg��@���!�i�X��Y��^Q_:p����B�����Ҡx֎
~7���]�=�H��(P-��t��A��2yʸށ-�n�[a���BG���S�-%�{v����cX��xѬ����@ja�i�oWd�����?���̾�}�v��y��W����F��ѐ�=t���)��Eު�dh�唀s���ڝy�r�*���`��es�$�_�i�����܋�2C��OqF�M>�~�r��I�wzm=}ordt�Z,�0�$tU������&���o���֗��;ԧ֌�C' ��1o%)<�ր5o?r6�ʫ�e����J�2c��s�6��׽-�u6�[��D1�qB����.�#��JȲQ�Yv1ϡ4YfN���
�|�v�'�޳D�&��R������k���'B�<;��ޚih�@���]��K�^�f) �����6ٞ�d���B�2RY)B˽.�C����Ɗ
Ֆ�R������	->�z�_D�QO�}��Ј���b��'���Uc��;�x�����^�jQ��s)��Ыl�z�/c?�� �.���)l�&���s|1� ��2����u�w_k~ۺ(C�}^x[֮^�,�
�h��µ"�e�M"������LA�(��H��q߫�	Nۼ�l�S�4���L9B��R|������ttTT$^�I��D��|:T�B�E�W��3��xSdw�C��ϯ]t������q�����9�nLl�gw�3�� �\�A��!�q{��]T�2Uf�*(��ɮ��(����*�mIg�I`ާ�wt�����r�\�נ{Dx~��f�VC��}�跌l�-�b��ճ��U�ɔV.������p��k( 1@�!���o�N���!�/�ʅNzt� �\� �]x۸��s!'|X`���S� �?��C�n�V�N��7�<�V����x5��]Q=���?�����g�����4t�nZ�ћ��@��a�>X���*�ZH��f߿�?���%�+�[*^����e�q�6�����;X{���=����/����1����38�TP{���I��S�1����d4qے�귊���73�j�~����y��w6�jqH�=�����GP�#���x��s� FG�9��8��P�;�3��P^�	��(���D�������y��N��|!Jzz)L�G}~$qO"�O�s��� ��Ϡ>�k��p����8�yJ��`(���x�^�5L[%Za��ȷ�������g���:b���1��`(��*�OqA�c$(��a}i�b^�,k��{0�gF��u%���rtXx�$)'��=��FH�t��]��PM�����MT���~�%T�Sy�\��	���&Q�<�3TJ���(^�4������a���90|�����b
r�8;V���ñ�q����#2�9皖鎙�՘�_���.�l��)�hػH�i��t��UEZ;��^˧�WYL`-�š����h�yDf��(�hE`�u%��k�g�*�BkD��Oɒ�$o2C`5"Ș�����N�]-��#�����g,��(Ο
���
<�i|T�E��+�j^ (��!E�w���/Fx�} �=����ίc�lFNJ6��^��Wf| �c���[�}��K6��=GW��l@�Aܥ�_Y��ೢ�-�&O|9�	�I��$�l��{����@�a���vf 6z����P��%AF�9�'�h�?�B��`����>���3��0Kn��)O�b�#b`+Y�*L (X�v5{��AD���#��|���K�ӯ^b�C�*�@p���W`g!�qB"em�M��9�%@I����ѪzG�Ԣ\~Jp��`L�a4�R�|�
�P�A���GhKO�}�k���$lʚ�� .N���݅����,�S�?�sF�ilK��� B��-8������ߤ%�w< ʝH���Й;�WW^��-�*TT6�Dh��χ׮4Q�^�*���,$�l�tg5��\X�u�b/@�w��/_�,&�O�K
܂�!�-(�g�BNSb�|���x�І��|�X BI
��HJ���c�鳒I�[��~��3� v�20C�.0�[�k�uH��r8'Dl[�e�Ut3��C�At���2�L��?h���6	��nn��I�;Tt���[ɐ���u�^'�V8}ߠ^�2+G�yW�)i�A��vJ�"�+��W���ԙV�1[���4/p��L:��LC%�F%h�7��
�e
R�5=kW�C�}�]s�)8��u�'�4���d~7���n���B�o�1�Z�ʔ&��ͺ�S�~�햣�6�[�̱0�z97{G��� �d��g����S�����[�>�A��+"$Ê������n��H���aO�F��t�A�]�Y�:��lړ����fItnIz�;?��ə�Hsn�Bjz�IQ�i?ǟ
3q�<�I�_5��[@j��cv�1�I����Y����Y���"��Q)���C5�����դ��K��fY	�0Fj�L��U�9c1���l�m����Yc���yo�bp�{�3y��S��(wȤ�G�Qe%j�D;=4�c�aПx��l� ��۽َ�B�VV�k�D�w����������,?�2"�%e��^/K9�04�Kl��.#�L,���<�.������qA�HW���$&[�'��S^���t��D�W�Y���<��* U�e�)�Su�m}��y�ݥ�S7�R�Y�mo�|�m�}��F��Ŵh���j4ԍu�
��y4[����@�V3�ta=K%�ޜ�69*dϙ胃z��aVՆ�q��K;�!��FꩲU�:vC��%�`"�l�[`�/hV�g;��g���/�&����5k>O٪��z��>h���Q���D�	�.��e�KC�f�a��X1`�%?���K�d�e�Q�m]�*z�߆ro�$��j"ב5���ӭ[��� ��A�ݞc�.��W%p��)��5�->�4�V�,�#�~̾'������6�|b)`��X��T�Ve)I�C�$��a�N<���#�O`��rP*&���d���=�`Ƴa�SZ�|!c�~��R4�(��bn*��9�qO������x�w\�{D�K�JR{���C���.�@f��9t���))���R"�S�Y[�nP�T,O��i��W��wp��C�2D��oi���q�H�O2D��=�r�-` ��R
m�8��2�_!�&w���P��� ��%��/T
���:���R���_CEU�R��|��F�3�Y3~�ST-�Ey4���#p���R����'�6�����#v���J�&��s�s�c&�{��(��e��T,y� ��%��+j[ܽҐ%K-7(�(�A�qO%L�N�����8Y����_D��0�qUt��~ފ����Ƌ5W�oC�ۭ���rc����}+碝k�W����ѱVa��dkX�D��H�%1� �Uφnj%�����?��?��X��&|SՋbOҀ�6��B���\���vxe/'��fU�Ό�N� �Ӏ�Tʻ�m7c`��>���K*��䤈���A������&�d$��g�����y�9J�发�D�}3;���H+��;�|��mS
1
�YW���E3?K%T����!ˇ�&��i��ʽuj�S-	�J��T+�������߭".�n���^+�����lᲳ
G�b!��^R��}L���.���6a�"��Ȥ^iq��U���?.yyY����\4��*EğG*�Q��g�ژu�����WY]B�U��Fc*�4�z"��+*#B��*��_���WQ�1��h<�?wp���4�j���g$��I�&����[4�G����6�4��ɂ{�dƕsN}�?0���v��	j�b��!.��#�Ѥ�"��qh��A�V������uK�E�#{�	��0���#L]L���<�;P_<,@O�AB���.�	ۤ�īD����|'}u��\���������:���q���K��%MZ�������!E�5'˽�EJ�Yy�,kx�J�f{dP���w�H���M!�1'�`#V�{ZQ�;��eEAj8d\CC�#^�w7k���޸��ZM���Z@_HT��̂�l�r���.~��%�v�ws4�s����E�T%-2�S���~�|�{�>QzO���;_ ����4��ﵵ^���ݕ-u�Ժ�����tq�.,^#b�����٤��d��U._�?���G��QfN0)���	U}r�\��A{J��� ����_V5�����t�ڏҍr��,
[TCI"�P��d�Q���xk:{�w����l; ��A<�~=��^8����DHJK������m��Q�����)fCLq���$�H=��!��i�H�4�Z|�L����ܵ���h%�����w����� �d~�ҏ+�=ƛv�hTב%���hd�Qn_�+��:S�.|R���\�4<DO��Y�UWv�s�ǲ�M&h�4ʝ����"Іc����Ԅ���(�;�ca:z��d?cBM�H)�wikgd��"�&.j�Xj�{Y<̊"qMF86�We/�8d����3�$�0*n.�:L@�.��Z��61��׭=1�����&��XsLx%˄��-6���ӷ���6&��Z�:~ySi���'�_c�2����
��	Yέ�^
fi�o����*���׀� n���xط�^��d}E
��=oi�%�=� �3VZ疳7ʪ��"�i@�.yK�h�|b-y���IB"��h�bѳ!^�z��a��;M�UKO�Sn�i��M�m����$�:D�X��v+<v]�hɶ�]з𵦾�˹<��^
�i�����QQ%j��Y#���w� ��D�}�6��^{�9[LO�qh%ڒ��@/ze��[�8��Z|(���>�@O��b�k3�KЂIV��A`D��œ���tNiR��u�}NX-g�#AK�W��p�h�g��|;ٜ�$$�R��;/"ŝe�W>r��, �\U�L~s��Up4�+�d�3e3�k37�h�}�!�����-��;?~�;ԙ��_�op�`¡����g�JH�U�����O�c����T��6:����4���HɃ��XA��o�k�}_
B.q-g�#��I)4���$�-� ]��Ax���Y��b!�Oz��7-v5�O�a�M�}�
�����됓�G�Ң�[����,0�З�3RR����l+L�>�v=y�������C��\%��ȵ�}������E�g%���J�Ǳ�8E�LH��$��=P�)���%}O�t�K�|J|ՋJ��r���ʷ�*2* c��6_�6���J0s�}$��A�M:e����bu\J��uޝS\MI�=:#��$,���U���0XUȾn�;����m��O5����D9%������%�6��QCd���h���-l)��ۖ%�̽�"��f�3/l����<���J�H��7�h7��Ce��8wm|;����(FQ�����?k�����:���������q�U�[#J���鷯�fx��#+��I�8F �T��z�(�{�S)F�I���9	�D��d*Hy�J\��L5y2(Z��S�y�ѠFL�s�X\%|������4S!��(W}�J�.�"9�����LU��jH7�;�Q/��KCӭ�w�O�H��D_�¸�W�'w�F��h��	��	e��]CsѦ7�
\K��p����y"��q,[�w���o�_�Uޮ+���P���ׁ���U��^gi�__�� C�䦧��� |�7�*���t��M*�o�G������Q��:ͳ���������-���MJ���i���m �Nl�흋�\��]5�=��+'���S����i

�"�>����P�K�2��?��/��7(�ó�e�!�_||��jL~d�Ȯ�_U7�]Q���捝Ep�P�7��^2J���8�/�??����d��V�9���2圔����JQ�G�c�;��v�h�ެ;-C���xV�8�eY"����	9��[oշ���0���1�2��;eF�US���-�zJ��tQt[���
_ݧl���r��gG_��/����Rա��ʤ����O���̓�X���GD��3�b�x�|}S47��T���c#�}���Y��W�J��93n��,Wv�Fb�`��<��' �;�˟��u֦
�g��:���V�S�!�D�me�]�ˠ�aU��-��G#F&��:@���FAB/?vk���0��v�*8���.UP����<�eK�E@ �!�p�@"��f���������q��� =�"�5�����>w�l&V��*�TM�ގ��2��tq �ԗT�LM�!
���|

[��dt�y<��LI��J����Á7�h�_�I� ��nf��X�F;�N'� �:�ޔ���=�+s�TW&�6����=�P����e�g�= �� �����b�ch�U�!؎�Ȁ�����Su���^��
��摢�Qrt�w�������˽U/?sh���Uu��0�?Sk1���dMЉ%F�-�k��atoY|Z���O���64�
�Q�������+�7�Wڑ E�EljĤ�N���!�K�8�o״����X�MGT�+���X�������c�i�Q։lM��������vrO-c��d�����]mgq��4"ȥM~(��L͍oy ��X�0r���W= .�[	����*�)��F�C�(#�i�5������)=��4�k� ��<{tǭɔ�<}
 ��K'���0�����yy�!^�|$��x��Y��Eo35�:��"�^�x;����7YJ�R d(�g[&<�h>��I`�"b3����c�f6߭�,�$�����ZVQ֓���AS��4��e�Q�\����1+���S+�<��|�mSp,R�3{T�����B�qʹS��S��,H�8
j��gn��<�[�����������BoX��t���O��#�mxWQ7�	�4�>�������2����m!���AD�\:�$9"<��0	 _�5ET��Ў�g�o�|kZ��Tn�VVVlϦ���3�y���(�D�[R��(���� ��������&gO� b��i��
�ʧ"!O$��_}t��WA�;^����
?��|�;6g�=��ګ	�	�嘴���uh���5�R�?��	b"Y�j��.��m�p��bv���	OAN�����H���_�<�����3��p>m��(*�������!/5��`����1(�C}���+'�2N�d��6���w<�e��Jo�T�[}��P��]'�4���h�ށ���ױ��<@�?�I&�V#�$b�3T�"�\!j��j>�}����|����Kg3�G5;%���.��x3�t�0�CfiP������^�:k<E5��t��ϽOt�~Q�,f]W�,�^����+����]�Voc�������*����,�t	����2�`���W���1c7�(i�� ��$�C��Q�:���į?hٜ��U3bf�1��Ǘ�0 ��� ��\O�(Z��G�����6J�wX/�^����� �`_�U9C����yH��5 e�4Z�8Վ"��Q���u�4Va��/q ˍ1(n�C%�an��-O��\qm�,�?@�&{��x$=��!*����M��]>�Σ�H��k ���VF�NN��)O���NC����ݻTqL8����v\0+ˌܨ�`��B�DS��,vc�O�ۢe#0���E���_�k��e�BM*�w���Z5��?
��W�$�kU�K+��q-Ј�XS')�aiAewv�G�^�Y-� (�O�Q�L�1<���Z�R���I�f��L�j9"����H��2�,ė-��l��Br�q�ȑ]��@l�hv������ M|qN�q���y:Z�s��@����r�u�fw�9���)݁�p�.�S�uݍ��s
t$�5�i���p0�#��,����
����O8fg�����^��Ĝ2-�* �'H�0,Z ���u}E��Ǚ&4w�����ĨNj���o�KyK�6�jC�����y��%��_���өU3�މ[��i�sU��aÙcx�`�5m��2M����mv�=�*�>��c΍VCu�H�Х��m�=�&��lL������[���d�e?ܗnu���Z�����!ø�ڥ�
���g�TM6�γÁ���w�����!�U��œ��5%��X,��C%�f��� �/D��	����B�)�Q#^�󙋫[�FP�oT_�h����4^����shyf����h'&�99��by�N�e�0 ��΋��S ���.��)���8K`�R�^�S-	Q��0���\��I;K�M��?*�V?�:���.�A4i�U�j��\����"H������Z���Z�&�)Sy
D��֪�g��;��u��M;�igi�������1'z���y+��P��ڸW)5egOF�
�a��c��.��#/�ĥ�G�jG��N&<��	�sq�"G,�ĕa9_Fv�� ��9&��].dq��g`z���d��#���ɇK6y
���R>S:#5��@�s���,��!�{���}��1u�d��J�I�\
�����ò 8�B*�.)oy���\�7����lT�����I��V檰1^%	K�+l&�Gz6�n��-(�%�ܿ�ރ����eb\�%��L�;�s=�+٫����n��'�l�t���d=If�)�>��3[�{�͡��&F�K�"$���w��o��o�6�靈X���r����6���V( ��A��x�s�=+��/��;(P��fj5��Au�%L�rAb2_﷔' Џ� '��4v^�.�C寶���o �S�e㎰��-2���e�����Se��&lЂ��^�< �~�4�8��?+�>�kP���'�#�>P��V��9��N�ʪm�!��]��c��*�2Mf�dU��F��n�X�Is���l���g�hmw��~�M��QD��$P~�,�(?����ji��(�M�QJ�g5;D����a��Aw�~��$� i:�染��nz "5W�a��N�v�_�Aej�1aՙ���Uj2�ņ'�۬n�p�єk�*T޸!Z�@e���//��4�ϡ�"�U��w=�^��M�
1���k1�U<�m*i�
���FC��1���&M,9�A��v����}*9��W�#nZF����Ӛ�N��[�q�qy�ipc��I�Ǜ8�iȖ��r�j�!� V��_x�C��
����2!7�9�?���'.c\�Xŉd��Q�g�A���U������,�l���.e�vm�꿃�=J:�Pwt����1%}{f�#�9Ľ���z�^@�S�+ƃ&�!0��`iO'��t�����].����k�y2Qa���ɲֻ b GWr���I/�?0��4/rߜ�*]b@KQ;�y	��k|����)y���m�`k8Ua�yK>|�"T��vM�z&�ȉ'S�ƒh>�GE������
��ЇM7_�Y���������n�q���UA5�Xv��x'���~|2�Q�F���.�L|�0BY�@��h�[	���LNY^�EBNk����ꄎ�66k,�E��ԫ^
x#(��jq��CΑo�!�ǒ���-)oΘ�3�ts�� "��WT楿�$D�j�O����q�qT�R���?
/�~�3�y��Ԝ[�	����q�c�/�e^�ޛȽJ�͟7u��������%���C���iCUc�?�)Ȱ�U�����B��\��FI�|�@�S�AIO�9g��FAF��*��:�ՔW��Kke9a�I�|l�	�]}�`��'���$��D?U�x�4�Q���L�|e2��-��5��xx%L�Y��K_S��?k�:m���,D�����I�͕�'�g>w,.�ӯ�7�D�����'^�JJ����U�^ܭ0mo���Y�|Fx�`?V�ٓ���p���������y����ޯ�N�``��"�Э9m��?^pH(W/s��ה�VOtPS%����_�I����D��bJx�Ȫ�܂y��w
�3����4��H�lZ����=�J(� ��O�m�3#H:�H���ƀ���Ʉ�7TIEz�����;gV����O�::���c�GU�	�n��*�V�:�
���
k��q0��s(�6�P�&��R)kR4ْ��a�3y�3W|�,�b�̹I�!��d����?��qݰ#��a�x?���'�~��r�4H���(b�P^g<t*���"��Z�е�PS���oq�O���پ6a~�h�L�_�v�n�~#���I V��b���B�N��Q�яƊ 1}�Q��Q�҆+�k��tN�ݼ�9G�g;E$��ۀ�/�i�o2�D�� ]��2�T�z�l�B��~�̓`���ax���^~��{+�z�M𧲲eS\J���Y&Ifo�G��k-
{�x����h�r�;����+�3՘���0:�k\ �v��p6nc����K��X��"��k��gڟ���14�d������V�:�8��}a���=����H(i�F���cъ�1��S�ѡ�]���z*g
)��In��X�mEޟ@�����W3��d�Jo��u���Ӕ?v~��)~��?:Q��A�7�q��|
��5���]��젗/�J����R҈�1c���,�X�g�k(H�s�x񢾈�2<���v�s�pj]�&�{|j���l���eɠ���d{��Ŗmn�d�e]�'tF�l|�uJ�o�����l�"����;����}<::?y}��c=;������f�����#t�y�,S�0/L��8Ͱ�5Wo����+��icüD/&>A�eё�1�}���8q��轏E2�f~&�:5�J�)��c9�0�L'\<�J!�A?���a"7�B�5��=$Q[-�9���bݔ=��'ś���(�U��ٌdet'�8��i��2��/}�T�]��H��\@��n��h!)çu���o��O$Z�Jf ��5�Q�NT�!�2��_�b
L����I�^0�(���喗gh����)ײ�J�H�k�U����!�c���-~�� *v	�B�����o=\���1Z������b��"��&oEZJ��0xm�5�,�U���gE������ђ^[��<7� O���P����h>�Nh�t�K��.�l�m�d5�9��8����m�^�3�4aUpܜ:�ʱ#���U��x?�H_�DD�Y�3��-i�ڽ�X��)�y�f�%S��.�i�O9�ӟ�&�~�0%�Ҭ�=��حF�ѽ+,��f�[��иw����N���VL�k�I�ͮ��B>8�^���
m?OpSU�è
Z��*I�il�ˠ��~v?�