��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z�����4��������8xT�(�h���/�<�F^[��V<v�Lz�=q{���ˁS�=Y��y�
��+J7�‿��(��ߑ��gƄ���'�j����/��b	 ���5��G��r>��T�CF�h��PNdi��NS�rd�j�FN��!X�fɅ=&t]������0��R��1�b"�܍��#��LJC�G��o�à���zz��c��Iq#����s�h��wb�¯(�"I�h�.[�Q�n�9��<:ܟUGS� Z�b����m���E������ЏǼ��DG� ��}�M�:�.6�Y�K�G���K�_"hw�Zd�b�\�55�3�p�SV�����{ꍅ�И6"8�YR_fC�?	�X�<D�-��9����Rp�4,�ඒFA���tQ0N�c�(� ��c�7�����v�$o5�h�ޗ.�z�`h|� �.���v~`��j�!�l���y5���؀%�q����!or��~���|�kH�Z���e&^	��P�c�N�8�}��a�:_���OH�@����
9{��㢒��T�Rs�]]I䘡�t�9k�2t���'a�Ơw �'-.BR\u�R��x����	�ǿ>�[TΛNG��(��"&hߛ����^�Փ,�/Oq�!b����D�S/u1�}cF`�C�:�w��-Ơ���}�Z����SP�����ihZ�t�P����x+�bZ2F\��$���A�u�
������XAիs2�(a��+T@0	Vi���^s�l��̄3� ���|���
+�h�x�.YNO�x�T�u�ζ5�� �̯�����7C&��<�\�&|�@ke����v��_��3�q�m��u�s��u4$φG�:=�w�i�"\Yz�$�ī������i�n]h�FP�߯��Ph���2��
*ڛ�6�E.w��_~���$JRc��G���D�D`x�M;nl#��� ^�AZE�#�NLl��G�����8�b/,I� p�30t�0��b
��ՑD �+n�W���x�s��G�B��ߝ�l��L���n�>�ޑ�Pq�%Q�T
�f��dc�S��u�7)�n}M^�D�v�(3���\����ѥęW��T�������N��=������VGQoU'3ЂQ�#�>�
�'�����9H��ާ����R�:R�-*jzz1��}�H��Kl�XM�J�����_\��#�Z�u����̄��������U���z"ۆ;��(b�iD�Dms	�1��g���=�]@���C�.cT��󿶭�2[L<�R�L@�71_=�}�,�[�KI�j҂ƍ}È% �?[a�����[�G=P�ݙ�4�(9������fR��WU�$ Qc��kkC��&	�Φj0�1C�faԿF�x�^��	@OpE�: T��<2	�ʪ�|�P�6y5�M\ԇ�	�q1fЅԍ���R���R޾B�����N��6�Sh�V�����*d�1�w��RC�#9��E{���x+TON:Q S��M~�b�޽�տ�3�K�U��,��E�CtJr�#���Cp.��8�
}��B)9�B9�菩�}�C�?7%��1�:�:yAz�m�
��c�I��h�5�^��ර�ĿrR��?���V��͒R���T�=�,n�Y���h-��>w��8w0pɰ1�Q7Ͳ�[�.[[�RT��e�>�q?D*�Tݏm��ވO
<@�C@��5S^׼�� F���Z�*{L:��5�5�y���
�u̗֒n�iI�����N�:)�?��p�i�͸�PT��R���X�� l÷����C���a��?���Ѳt ����@-�[��P�q�(��Ik�u_��`�h`<eDH��@����W��&����F�c��<Z\ol���S)Z�k�Ϲ!������≠�}&r�mQ�H.�`�K�(E �a���C2�x�����L���u#�;��Xk�E��0��5��}�-<!3�Wo?^�aV����0���Ȱ$0A�&��W���gc��Ǉo�v�A2V�8�\�J��hn�������I;.�<n���x?uV��<����p�>�uc.�e@��t��#�`���㦒�e��_�����b�߾�JO{�E�f��^<�SW;�g: �B�����1'�	o�}L�Bѿq��)�bZ�Cn�ّ�GWp�i�ԯ�Ž���Gv#X��(x�J)|���B��R���+��g�l�tĺ}��������ț�b����
��b�K��r<���P�H��]B�N��!h��6��z4b$��.����P������$��Zk�->A�[�6�a���o�fRC��~�zbN�E\/������C&�����������P{�6��p�:���E�a�y�󥪌0;摕sWr�����,���Ҙ7��0���(dST	
{����1�ȜwJfB�v����1��P�3�����Y���<Wc�`��2 mg�?ÃҠ1�Ob(��{9G�ڵ;݊j�6�'VP��VX⎢);'�TO���C&��y�2����a��B�Tk	��y��\<�q�wl�[��K���F�@n.���1n�V�c-9�fQ��q�@�����z��1�ӕ�M��Bn�Q9���|d/�k(.��B��/�e�����U �������i�.��8��[4�����3�~[��n��36�#L�8�s]�[���T���ر���jG�-���J�.m,��G��GC\�Z��F.�W,��t֠&Vdq�%Ut�L �r���t���p��}Â�~�l��A�D��O�6��{��dnYeh�ud�6Ұ
�L��׵��,Wg/�*$A�
����'�!p�Œ��0b�KNpi���:iWv�^�p��;o,��t[����5��������#5�XI�5ậH=�?\��:Я����$YrÆ���^���;��ZWZ�-{�S��u�V����V}W�P��f�����y����dt.�!��_&��zA��",R���
�V�Ma֋Ȍ[75/��߃��]���Cq�D�؝����4Vf��7QC/�k��Ⱦ��:�a��$�N�@�5�X�}�.��|M�vZ�i!vnKa�3B��~C�q�Z�yuDO������k^��~�+s��p~_����,��K62�r��h?�I�}nJI�.���1�E��3h�?���F*�7����̛u)�N����|M�Åo+�9���w������1�6���K������:>�R)�}�ʉ�M�D���M��JGFd�}Gw��r�э�k�X-R\�LQ�/~�	mx���O��=�8E�^ ]�3����?�)�z{PI�C߮��J��k`f�����M��!�gΓ�a�4�?������I�O�,����j5����8����(��%y�~A6�רP�'T�+�zWRɨ��'� �����hC��T�V��ת��J����ނ�^EBr�/qa����v�m�2(��O�W�E�/E
�2�r��l꽷��M�`�L�Z)g��>m��03��]�U����%����� ��a̛i2�Ut���(�O\X�"��(�|�qF�n��&��$?y&��a�,	O�g�f���x�dKA6�k���#x1(�R2Bf�yrV)�f7y0<ù�z�N�o�w�UI��:ɒ�J����AVi_0����G�*@�mB:v��,��x���2AK�>��������D��(1�MP��:���,�Ξŀ�P������0`m���{��?ˋ���1b�o�2j�?���j�	�I��>G;�%���	5JimpWgi#f� '#(�S�`ꏕFK�׆��aވ�q��\8��4#Y q�s':$�NI~����j�D3��7o�T��� 	ft��۞���+z���3,����B�	�,7�����,wZ�!��D�.+� ��yd!��/��}n�]�����Kqrvx[��t�O�w�6�3��k����Ø��9T��g��KV�QqT&`�జ����'o /q�佱�?c3|��v�G�{p���I��ǓL!��!������_`��<�q�d^�!8�n�`���B�p�P����TN�^�*,�d�/� p��K$�<=|��ZĴ]�?��̙��n��lҀ|�3lL-ic�����䯔�u�zĸm�"�����^��#�xp��Fo����aPDq@��_j����><�7��M𨀴��"k�����z]�6�>v 缝��aC�er_�*aMZ�0���|�|��o�]�IvѰ�ϗЭ�E7����3eԗ��=�o��ٜ��~��Í�Ο��y>_\pd3s𛏮\�Ek%��A��荛�}R����F�F�8�YlUuN�ْDyʦ��.��w��cM�'(o������ů��OB7*I�����^V�X��zg��.����јP�3�o��N�W{GĢ*�zse����{�}�o�������Uh��)>%�lyY�(G�v�)	!�����A��K_��~��7�*n6̭ݯ`5z�vh���@�_�˟ɼ�x2� �t\�m��~8ND��~��x��7�(�k�Xb؅Д���N�v���$Ն���'��,�>�4����eq�v�]��w����ο�^:-?zES�/�X(v���F��o� 1��P8�䘢��K0�����ɺJ�J|@�5���*�P	{1vF��f�Ae�ṛ�o!w($k�3�ek��u����GF�#�-�s�zAN�u����hm�Vyq��׿Q;SD�e�h۰HG�B*DR�T ��gL�Do����D�P����YD<�҂A��c�&`�`����
Zl��1��ϻn�˥&��O�����R���X��CP	%�2@�R�hF�W�,iܐC����݋��Qm��ݬ�{W���dK�ƞ�_�m���:c�J�ՓQ�8��_޿�|���Qː@��?��E.��w2�E���Rˁ)A�V
ێ��a��w��X9ǡ�ÂǤ*jr�2���/:�d�����0Yc�$}"��4�����Z:é�X���͏���;M�cE)�sc1��6�M�}]�#�s�XS�S�Y#7��� ��'�#�~�a+Iv`����\J"��h�ି4����
E�_�͊�*������d_i�H*��7���<:�~���?S�øez�� E!A[�n4����m;ۙ CN�x\�m���ě�C��ِy�I�:�'���i F*f�V'�����߻��;֐�C�y���K�oF�}�cTԲ��C	��w��1�\�h�R&w
�o¹��tҫ[X�0����-)
_��o�8��g
a WO.Ul~�]W�w�ƻ��1�f?�e$�4�K��6'��1}�"q�����\ǲwT ������s�Ra��G��Yh!L] �J;k��fG!,�%���M�_K���{�j�s�Y�2���A�?G�Y�� W1x{������J����	���&́�+�� 	� ��<K��DB���A�]y���9ݻ�T���i� �V��~��#ܶ|c��U3>��KS��>��[MZ��q��+�,y��р%TH��ZfLy�|�Id�Mb
��fp�`�@���/{�W<���٤a:Ӷ�C2Y�*Y�S	�	�^���_�8�O�[�)����X�<f��w���{$���H~���+}k��$-K����0�Č���u���Eӕ+'��&$h�����r�tf�]�b�F��g���Mb̻`9Z��n0U�
�}b،�jK��`x!�b�(����|c��\	g�8��np����9������N��m�Qʥxv����,Ů� `�jX�e�0�1�� �7�r�R�����?���	�����і���~�i�]�Ѩ�i�x(<�wG��	g�v,�\���,��T[�,�Ks] n�+g��v���U�ԃ�v����10yh�1̀�����e)��^�+�ߋ�I��琄�vy1����c,t���ՖI��d���욌��?0O��xů�������%ߒ^���X��-^�t�P�(�g7�Vo����8�v�.�޼�>Z�	L���*�����Qv�x�;N G��fu��D⎳X
=�9Nyې�'6��5���c��X��~+(_�Ho�"2pj�цLG=C;��,lT�L&(&^w�ɬa`\�(�.�	�\��8�G�mH�y�$��(;����)��p�0L�l��G1Ԛ}K9�Eh��0�۩���N��h9��TY�La��{&���F�^L����㏫�tָ���*)�l|4K �����b�
����m�4R��+A�Op�K���۠��Ane�^��*"fd���+�?�e�{#m�8������L��@�*�][py�#�G(��R��B���;`ɢJ	��)2obw�ey�P�!
*��k%���	����_X�:Mfc�գ y�G],?u-*G,�S�Kv=�
-�W�E��a������wJ%����gm�6�ꂭ����ꐶ>D�~�<�ZW�TP��Gp��ځ���s�E}_풉�W��KY����F})���2�=;�T7x���5a��b�o9����.�ŰN8Ʊ���8Q P�
Rۉ��;�L�n	<��z��C���t�1"9��R��(��Wz9{�!���}@g��i�����{��t�\u�f5S��(����$�=4k]>^°����x�~�"�9�px��	w�C=����;�;����~�OJw�k������-���ǟ���a�O�b5v�-���-�6:d7
��Zejސ��k1�"��寤�ސA+�U�z�RP�j�`ٯ�@}�>��]D(ܚ(��<�}e�P���s�fg�_S'+�f�	ȯJ�"za������8V�qYە�j,��[�}�f�H���
J^�o� �ג�	V ���;c{�&y���3�}N��v�ׂ�n�qqq��R�ǎ�fR@�X�Ev&�F�X�N?xo��9k+�7��N��(I@��N^���utS���b^����6W���r|�Q�4d�g���\_+B�dIv`u���EܴzƟ&��4�~�G�6�j���T�Fxam
K��r"R)�]v�|n��Z��.���[ƞ?�_GMʏ$2M$�
��TQ�bxN��ڭ�[�Ock<�+g�X��Y;����d9��~(S^����EUL~A��D�pH�y0��Mj�(��3���0�]6G�WT�[�ס��;���w�cz-~;�F딬p�
�.��q��an�XZ�e�xD�p2ati�6�i1cOs�� �2LeO"�&�>���A�sm"X�F�~-�{Wʻ��'_7��!��}�ۭf=\ȢF^��T��>�����ۖ�o��v���<�߽k��+ψ�����*�Z�/�n��S�{���0�S�7��*�O����_�B��Έ�G}�t�Y̢6�%�Y|�T� �`�2[�n�E�S����_u|Z�+��ۊ>_��{,�k=YM�����'J%kIWx�ZI�����S���/�]��k��L2K9���?����2��o/.P�*;�2k���}F��������Jj�~�E�Q-��p^��T�Ut��1�4�[�k4:��}^���`E`j֏�k3����i����\f�����wܻ&�[�ޣ���]�} �Nz��83Ph�ϴ[]?rJƌn���NO�M��ʙ��:&ZS��Q��o	�fq1ؾi5�_&~�wX���T��D�Io(�[�4i�c;�)��L^V��l�A3�<Iƻ5��`ܡ�k��g�ȣpM{t��T }o��>��eh�t�ժ�ܷ)o�I�Dў����f9;h�%��Vr��}�nݩG��+�%�z*=��^뤻�����'D��Cx�1�����i��0����"*S���}�l��<��d��֜�d$��y4J6s�����=h���;���h��fZ����H>��C���P�~��(&Q�[n'.0���{H#��������T^Y�un
<���e�"��܂ �T�jrìds�3>-`�^��V/�F��7�P�$*��T�5H;��HW���{I��,/kE�d�N�0�j��,}y����ME�O�~_�^�t�e.
��mme,�VP���'������)��?�4������p�9�/�d�~s%խ� ������t���OD��7�;��y��~�GR�J��LCccU�	{+#r ��y�>�!�[.ъѩ])w�ut�\��L�)8w��Q<%�r�0�6��-$Y�&-�D�H�w�Ea��z�Y��H��8X�Ã!��/�]̿��^�*j.C�	}q�
F�+�0�b�ѝ[v�!X%�OI�,��K���M>y0��������¡4 ��g��8D��!Nr�f�f�ӯ�_�*F��ۢ�_�e|���Xϓh��L�����xUyc8r�k&^?�;��[��1af]�2����l�k�ό���I��y�Q����,2���� #�?��k���s������hN�٧�+8�?x�"��Ā�bh�oC�����=��ܽX/�~������0������@�"�2���.e��(S��.a�?6����C���s4�~4ˌ�bŏG�U�kS��Z��\3i.�X��0ԋ"0Q`0�KП���N�i&�<,��N_�Z�G��Y�h�~�m.~��H����2��ٵ��[� �c�����;�SF��M?*fT�V,�Q��� P��O�z��|m��]4��??hG;j{��僯��q�W��p{��������LrVE���Ȕ�M\�T�Cƪ���r��=ї�/Ag�k�F�;F��O�-�YEC��%��+�������5O�*���$JI8$9����?�q�6V,��3�v����B�!�2I xH�-����03��
&�����lT6��y*,U%ǅ�aZ�#�2 Ǌ.��MI}�}�q��âR�?�-9ӟz� �kk����2��/}a�Dx>%��w�oP<ExǑ"�����!Zܴ�;�@E��룒ʞ� �ޝ����}�<o�5緼�|ݕ�̋��\��5:�� ��
�k<]�D��{�nd5HjE����T�5������2G�!F�l�|eR
��B�(��� q�!��l�h��'1u?�p��@ߝooHU�0t�!������n2�b�u�^5������]�	��<�L�~"�)[ ��fX��s�P�C�d�Xuc����p[�!��Hx̷'n��k��R�&��r?��3��cOJ��	��\��|EA�*8���_:��d1��j�/��T+�����8^�a(E��3����k��_ދ]Nymt�tc��k�8ї���_�o�F��-5d|���'�4��GDb{w�OXCI��(��f��}v���-[w,���xÐ{ݰ�Z���{��Ϯ��Tԅ��Rm򖹌��������f�iJơ	"�� 5_�ꗇ��:j��1P�@�F������[I�ɫ�j��I����2�iwj.Pws�H6$"�fr%�U�rS�y�i���H�]�" �sC���p��[(i��@��RE��	r�v͗�_�c��~�{�m�]V�꾀G��
���W��m�-ɑ�6�y�g�/�	�rc#F�;k��dvԕ�yc�W�(�e7�2�G5H#m�W�q�\�^\I��#I��Zp���:����TE�� �'��<�Mˑ��5��G>Wmo��[ "S�^6������al���"��+�B��u,d�E�=�t��׬�U�8�M<F�4�sa0�J�V�+�)�
8�u
b�����Cjx��+[�x��X�}m��WV��ᕙ�{D��n�x����q�ίdv�μ�����7a0����B�.�y��*1��d|,Х)y�p�Vh����@P���0;7ۣ�K=���'��QJ�v�m�\�W����^6^��V�?�[U�d+'�A:~����;w��uؚ���Ky��R����Ю������}Xh�4[Qm>�$YX"��a}�&v�+��ۃ�İHK�x�x�@W�X3�n�Ǚ��ga۪�y�N܄O�&�w=@�v���guB��W_?����L��-&�AbrIڋQ���*S����Sۊ�>��{�J	���X<��<�I��J��:�S'��u5�&�+
�a�*��D�I��e��f*m��_ڰ�/'$��� �tK��a��"���(�
����o�g�et #��1_�Ȳ�2ɢsHKP-��ۄe ���V�\iPO��V�`�7*�߈���#�s�s�G벪LUg�t��A 7� ��<�R1�ޠ���3ѷ8u��e�2�g���rb�xY+e���TНD0�M�m5.o�&	?����4À�ad3���!����G�}hAK �:�9e�h� ��6*\g9o�Ro,�#&�C)ݴ��rn��v0kN��]�D��&�h�ng y<���,Z�	p�|=�Y����eB��Q��"]�I9�l ���o��1�C�[��KkÀ�xDI�~��t�@\�F4�n;�	�5�&J�������
��0�º�?�_�}8�y�#Z���k����@x�o�d�玡>�ደ�ltv˓]�Z����T�uN��Z-eSX>Dj:cpJ��ui9��!Di���D[O��}�����_�1��Ѧ��1V/6��*s�a���dNAq"�q�����ms-�*�u?�k��B#]u�Ao&�""�&�(Ŭ�M8DK!7pތV6N���n6mf& ����/Ʀ�@��߿��\j*�u-�U������t�m癳�isq����{�7��K7� ���s^ٺ���r�۳�r
'�R��ӵ�!�:[��4�>+�$ę��%�oy=ڢt=��x�t�.UQ�xڄOkMnU��3�/Y�є[�u>���,섿C(�?�S�XG+�h��"�z�R�Y1�c׹�c�&��󇎔�]N�0~���LƧ�,y�)��=f����h�3��|�!Z�P[��@"�FJR�h��iA��!@>JV�,V/@����]�)�i��g��h���[I�"+��C��ӗ+ś*�f�Pđ����..����W	
�X�*nIz�t�� 9���]���J�A���,�t\���ږx�BB��e�ܛ��3Gz��?=H�[���aK����85��L��_J�*��p��M!a�"��}��L�㫶����FkzoayEc]%-��;����t��Br[��Bqmg�n;l�QK��`���x����xy�jg �qe~/l4!%��#P�X����y�ࣂ�p$�p@ۦ[��r��M7�lm"0S�$o�օV_fBIJ�Xs��o�a|���	V��O�;}�1��3 @�@X 7��r]��L�Q�֫ 'n���23���n��kon�<�q�d�4���,0��f�C�d�|��z��5�&T���7Ϳ1婬���*5�������Yz���N|)Kc]���_�P4�hh`.����4�EC	��%f�S�gȫ�����u���i�Oڀ�k��U?Idq���� ��"tn��!��5S��n��|*'�\~�bF�X���z��
�\+�-P�{���[�C�Vva	&��8��w�7��ݨ� �}���u��F0�;��޸��:y�Y>�p',�T���ݞ]��<�`F<_��]��ل��"�����K����N�˦��͢�S�xuȌw ��/�5jq�-M���Xd�h|���#'+T���T�.��l�o���C%##��r"��蝖ͦ��y�T�Z�js�.A��O^�� d�Wne�-���]�a�u��n�B��F�R]ͬ�c��ǆ|��1u,�3L�D�t�o��뤢�Q&%�c��7O�Qk"~���]+[)�m�Y8��p;���h((�F�҉�<�?X3��oB��V䬔�+R+& f���b>����������g�[�4$\�mknW���&wkZi�`�a�$!��,l�	�g�����&_��p�.���G��
��u�w�=cy0]pϟQ�#�>���I����اt�l���	�-�)�t�E����b���+T���=�&M3~�Rt��S��Myއn�\YW�Ni�k�x�hd1k�k������*�E|�� q¬%��h%�X r��l����@ij�JG�.�d{*L��n&v<���Ly�
�����<�����<2��=�Ʌ����_Z6���H-8��<�ޭ��5�Z�����La����E�X|by�a�Fo<���Q��<�y�e���\g��Y���e�v^�W�*���� �;~f}��&��[����e-����xH�r_2&�w<0/cg� �F+Y92�4-�TRZ[�W��׀	jD�,��!�H�+y�_m��'�]"�f��Ԇ��b�mVm��~	R���[�hMF�	lH�HJ�ڡ�@�d�hS�� Y��:�7S�FcV���������w��[��(�?-y4<&�b�H^�{�̳h����j�bbj�τN�&\��1��WX��٧��+�J\����W�"�2L�˅ ��y<x��/;}4��+��$WjZ�l�����0�"�_ۋLKJ�^������؋/�!�٠��3gY����ez�7��& �+
�o5o�x��
�6�K�\�3켤k��j�����W�XUZ��S4��4/ߵ��8�E�_���XJ��c:�\�cO�ĥ_��;�{ʯ����,dO�t�@�z��{5�='�0�Q)���d� ��ur������z�s�,��Ё@J� �,C@S+���"��@ʹ�4��z��6A����(�v	=t��}���ɥ�q,e>AoYT4�M�$N�����rz9�}�M���]GP1�����0h	��PT	GݖJ�P�}���|����y�����ƭ�kWYxJ�hLv/��ەS�#��_^�ዖ?��1 ���"@�醗F��$1e���d�hw�=�i��7`��Xy`�%#�Of�!��D��z���ع�`攳y�_�۹]��G�V�Is�ߓ�S+9�M����+��Iˊ��E~Y�X��(��>�����8�Qm�?��z�&�ӆ�������!`�S�+-��G��)��Ĩ����T�b��t�`��2���rZ!А߽K�f�Y!{�����W�� ����#��ʚ����(�B� \*�����` �@2ճ�?�� �q-�7�?U!��4׳�
��⩽�r��#�B����]s�z?�w�(E�"#��w�7�D��t1K��(mj
�Z�8���:'.Wߣ���hE&?G�˄�c�</f\��YBw� ���RX-끾`Ʊ{W
�4�`�֗�□9	M���MO86�OǬ�h=����P��p��)K�9v�R��z�'m��Uj��o�]�>U������+��2؀c�g(Ò��U�ϙ7�|^����@g�� t��QP�Jl��SyzG��EO��$�E�>���aw��F�%I��3杋U�7�Y��Co���<)�'5K���6]�p��We��G���zH����)eP]jV�Z|3��(�i�vpR�m���g7�g���T�+��<rzu��=��͘%��������
C7貱����u�ᇩ�b�ic�{B�[N�C�1��)`�=�W�33��ь����&) �F��ըVGa�k�fψ��7\4�	��S(;��u`�A9�,c�׫zP�"g�Ct�%��l�DB_�2�yqӨvXg`�[Gǈw�]>َ\���>��L���-)k����
\ϫ�Ou��"���2X��v`H�������n�ﱙ�v�&�3��n��]��
���o�҉#�)�J95ҟ�c�h׳5�������Խ2+�^�F	72�q�)�F���%�j�Oݞb]�K,��71~"���^��)��6vi�wi½�&�~z�4=[2��:��EI^�����ד�Ӆ ��U�	$���J��G�e9�|~��KB�@i���z����F�;��xZ�B�<m(���ǂ:���(x�m��:щ�p��m���$�v1�oW\�s�z+p�y~n��Ηt�{P��a�(*O��9���rc���d	�̦x4|�VM2���YL��(�%��%�ִ4��|g��U��\z��#����x��]mʿI�p}�J����e�~x	�&�Ct��:�:���9-��Э�\���WЎ¸j?��B�s�o��z�y$)�Q�Y��6֖󯒓 ;�C���W���d�����dp�V���;m��(�$c_�$�-�)
�|�?6��S���)'\-�g,=�n��]o%c�[]��͹X�!�~�95o����F��u��Ʉ��~[��zxS0���1)J�@Zf�.�Ƙ��7Z��K��o��0������t�ݍ&!M���� ��9�Z8+Z�WQ>:�d�i��(�>7�N~��p���Ԟ�bO��b7�pB+�.�J���#��8/
Ő��������Y��7H�����O��r�"���HNX���kP~�^� �1E	X�F7T���b�/��NyX�~`@�/���:���
�r����!O�'�;鵹��^�w]|�]�kЋ(
��컲�/�����s��R*�6��e��6h����w�-����#xB���_T��t�!ߠ/'8dn=�ir���&ϬY�yS/FO0�,�����Bv�iw��-���-�L�F�-���e
��k���'�e�~4�!)aP�2����Nf�)?ԍ'Ф^�^^�~kX_���SՊ%���p �D��7QH��sow��voS2�46 mK�cM0�I�b��+�f�H��uf;�S�9Wm"�A�@���7� �E��b*�V+Px�R@*�R�B۩�[_rm�2q5�D���_��7Sy��#91���<�6�Lc�$���$d��җ&	
G1Kvq������|����vLl����YsʁX�K��ˉ�h��FM|���cʟ�0�7�A����_Ʋ1�7�(5��x[@�$0w8(��رvIěf�E��hSP�����R�	.(%郓�'��Ar3n)�� A�~�$�L���rK���R��Ű뻝�z�O)FЭ0��
����%���.���3�E� ���W�+DXi�Ņ�T����H9��UKĠ��c&|�=��?�)K%�����Ę��(v���|�U�p���W��68�>4��u��E��T�؛��$����J[z
�)�B����������&#R���� #F��%�&}��dT�m�L6�C��%?"���X��t��Y�M�U�Ԯ����^(��%�vV3r'�#��2��j:LC� J� =[e�/-�wU�>V14�'��6�����
wl���,� ��ev���0���0Пg�4-3Jf�RG,�
h�V��Օ�-P��D	8o(�V���,�G�x�ܕ/F��@I�e��좮���V�ǷlFT�"�K�4���ˇXRǱ�zK�	R�DJ%Y~�Q��f�Y�;o�F�Iu+�>��x7,�c%iwE���P�ug��ʈ픲�2�$ <�������	���i�u��&t�N��k�k��2\0�JS�J-�qE���#C��j;�<�C�g�|�i3;'�h��4܉o��r�Ч�������Y�YA�����J�ù/g[�/��Ʀ�0Z ��=|H��NPTV9�?U_Ո?(��[D����	�����8�@>x�I��u��Ň�K���Ș��{Q�,��Y	�������:4]˾rJM5;g�-	f��_���7��.W�$����?nf���s��_8��ן:�-V��ݍ29�x����|2Ϣ^���-J�8��V���m*�~���P��#��\�+�{�<$�~�����` v|Sf�d�*������.���mB��p_TK� �~�Ԝ�k�b����&3�$�Ft��j���Hs_��I!��$e�6x@�C�r�2��;�y�N�]ѧtx��0���$AG�G��[�Lf��ֈ�iLR짾 6��åb�c�$���D��w �mɡ�*��&�r�!�o��#��#��@:y�������@:įVѝ�ä0 ���������C�o����|D�� ���=_F]S��3�9�;�P��	[���'�Pu��Ew���� �Z�H-�G����@�w�rO�ݪ�Ԧjg��KPx-��U��hO�B*��}��	�B�@��M�Q^�{��1#؊`����h�n�G�-��U1��'ƛ������W�v�@]ȕ^gI͋I(k��vIIt���yPm`e=�4����>����9�vd���;����4]�U�C�����w��E�&�]O�w��r�!�6��^��� �F����<.�h����u����:Ԝ`�o,���}�`m�8ka0�B9A�e@���F&Y����#�g����i~���:�=�7��L���j����r�ݳ��kH�Ä`�ڧx?�d���r���6s����D��������%[�B��]˝6�L���Вx�?��S�d�P��U�3Zw�C�_JFn:Y�~���I�6�u�<��^x�%�Y#���yD�[��il*
o��?*TD��_�����iź{���oD&�k�NRUk��$��Ҝ����L���vʫ�E��:� g����� o�An���T���wӷ�C���o�o�/����୉�Y�ꍲB���+�=Y���㾀o,��H��	�J܌����ӋB�A�r�k|���;���{��BIΣ��0Ou����O
b�	�j�琩�(͵/�E����L�Z˂�*=s)�D-i��]��ɉ�R9���3���2�$.pe' �d�O�~�i4r)�5T�8鬬�WpPS�T�\��5W�p@:�`�4k�==�$Z����@��B���>?T�a��f�kԘ
NZ�:�y���6ˠg��h��&�4�Ògt���g�N/�����⚸з����΅ݴwE���2Ғ%�J�� p�.=h����4%u���R��<Tkf6� 	g�����ٵc bc�v���Ϲ���eZ)���=:�E#�(�ε���W@��!A.�Aa����O[}�[��o�lJ�s���)�=�_���G�����G��O�ۊF�wEL������M�ir"P(R:�U5�{���[E�1�����I��wyҴ�
�B�M�x���)'��ۼ��<@�-E�Z\��Q3��QF�x����鴧����ϑ<��L[z�^���R0�~)�Ͼ/p����5_�cyT��iY�
����H5�,�|��p��|ZXIޅ���(s����
,�_��&�y�g5ε#��&
S3�z��يH���8U�����t{�Ȭ�Ύёf���Vo��(4ys����HvgE�%'�p���5��%��՛���y�ì�1������zI�v��枖O_ؤ�C���3��5D���a)C�9���=z*�M�K_~���_N��mb��#�V�W:�H�ϋA�c����9�f�/�8Yɡ��q �y��ijaJ3���,���$B+�ec�$篝��&6zy
��T'�~�SF�>�v� Hs/�5�Gg��y���?��	o��vq!b��д����:A����r�h�'Ԫ%l�Xj5��TC�2`f�1ҽc��'x�K԰�CF3��������T�����`|ZROA0�<���.nQ�"��M�|�~�s b�����W������%j�����6�4����Dɸ�B	aK��j�П��R��H{��>����x*�2�p˗�/_�Y8i���TUu�������7Aӭg�켨RM�ӧ�ʹL5%R��Z.����u*6~���P+E�������|��n��Y�|L����7��b��f�b70@�WQ�W�u�ή�*Pj��~/���#z\�Ϯg���a�T��-[���q܎ƪ	|�蓬s�e5�Z�����]�5����0�,�����(�(� ,\��x#�}�"�a�����	�&[�uK0V�;>�f/,|2�!��X6yx�X1VM�u��-.�OXK��
	�-Zʀ��d�0Bdn�~�2({�.z.Y��@j�����$ϓ��jS򰀓,�ua�qF��N�t4�%��ɇmB�u�YW��:�)�Sd�����p���G!�`��0�oe���Q�`��u���W>��I�B0�ߙ�Șt�0�^ɗFpEYQE��f�4b�z�b��2�p>u:>ĸ���׀zL5{d��g�$ΰ�&���������Цj�bf���M��|!:ь��1磙6G���*���@H�!�fb� B�8�Lӧ�I�=W���� �n,(�v� ��w�P�BM;ODf�58����s��N����M����VP�I*�r0��R�lc�����%g��:��.,g3ma/�09�;�qL���^2�
P(�6Fg��W?��w��:�`Q�/3M�jc3���i�m1g�蝬q���%�� 77O���z
�Õ��r�V� �����Z1p�iJ�Xnτ� �l��`�ৗ�F������G̳ؓ$�4��ZE����˘����ē~�ţf#�R"0�o����w(Z��뮔�s���-���o�E����	����W�P �'Ӛ@���d����ׇ_+
&x�/ȵA&'�@�B=��JWh�$i�­E�ƨ2�#�U�7���������?��`��lr�X��>�LU/)#5��H4�^�ǡ�]F����FJ�|��E�Ur� ��hP���k&��!�$�.������S�Z=�I�ת`��F�h���b�d�Ъx���%Ar#��b|^�.��t��A�	�؏�Q�;�c@|sh/*<�� �Lg���m�����W?b�����$er\�Sܺ��f�O☊V�4���4rt z�h�[<�!!��KC�l��BW���Gv|�9�Q�$媼�b'��_��Ik)��F9
���o���/E.O{��G�f�`_�E��z>I�oq/��HB�����@��F�E�	6�M(�+��`��&��+�Z����3���v�]���zI��U����/��m��v]' I]������u�s��[?��jJ��
,�e���-0��EǴAuUYZ<ؐ�?���p���pgL}Ga��qH2��a��@�r{v��+^���U�$��)/o![���ֱRc����x^��pQ"������ȏ��,H���cǺQ���'RH�t�8�7'|�^3Z��c�v3��"oz��l��\�Q%��/��~��i���a�yP�=�;���b���1�,\��g�_�H:_�|4[�ޝ�60d��a��KP#�F�䃬�*����b����n���n%������
��됓V�Ʉ#J�C��h:�1[����Ή�?�����<°��~�1�Ȧ�����V7<��A�x�=�	���KCc��CD5�0-�%�ė�E���x����44:*�w�.< �R����Xl�|7��CcdɊo�^�?��I.a�HUQ�c�����������TƟ&��N+Ӽ�03�Xm ����\���Bv4�o�a�,äe�ق�;��
$���!/������y+����S����:7�`.9F�,��JSn\��	t�������ߍ����jU�Sl�+eV�O���5�� ��������P��ydW5�ku����!���9�&8�	��R�2_��g���ʺ��'�GԬ�?�_�%�z^�r�~�/t� �n��ie�N[��$&�ϳ��\ƻ���BL����f�I��-���,�6�¥`�HB�/j�޶ߍ�2������Β�H+!�>�+�q|k�`>�(7t|Y������k|+�c#�턃+>NN��"�B@W��a���I!�e�%�G�XSK���.\O��5��G$�I!Z3R�� �{ay��rC��`]]z����0�o�dl��u�u�¥߻��y��Y����Ǡ���P�z)c��r*?�*	2�>@!V�漢�����&�»��X�զ�~��P�d���w�ʇ��m��&����bv�A���dbH|)�	�q�՛����f ����	�k%�!���U�s֑��������0FK��K��Z�d�ъwtuq��	C\;�hA���D�7���ڈ����[Z5f��a�>�y{�@�����s��]d#��.j>��4������9��	�͵.)�D�*9p<�"�B?p	��6��`+�YG����sL��2���`��p����g�[I���`���|6пؚ�8[�z�����0ZT�؈!�e��_�sr�=zD ����0��6�U(Me�@����2K�����no�TA�+��
E����-��ߕo�X:�dj�-Yt[�Z�X���V�:f�q�=�)/t:�[��UϞ%��������6q�ֻ���6.�[�x'TЊ|�Z&Ʀ$)�~�^폿6m'�s�BD����H-�6��ͣ(O^N.l�X$�:��j{L���Ȥ]qӹ�,.��r����.��<��~����&�{h�=��"$T�TN=Ϧa�E6iNٷ�+h]�"�>�ҙwG��u��E�֋H�!�څ�s{�����hu$3R'^$�
�Y3o�]XN�<i:�q9m}��{H�F��*tf�a��S��}��-�;��T���	.��GcS'c���z��xs9�	n.5�`���tV�4l� ���Q&�s���O���+<�q��s(^�� k��i��sM/8��2�av��7�~Ř��}�4�,�b1i��/
	.t�դѧ��1����s�P��X�U�
#~��Ͷ	~V'7����j 4d���魰��]�
"��)xTwS1u0�&���HokR���_�A�
uA��ݒ�ILH��]��<�4
N���)MtE#A\}B�$z��Sa�u��w
RU��NyȆ*��+}^��L�Y��cg
k��u8�/�A��8Y ��pi�����D
����qd2�}̩�4W=�^2#g ��A�����9����!	����D�x��Y�S5��UW����Qq��Bk�2@����l��h�`d�l� F�Q��mD>f�z�Lv[uap��W�٫>4Lޛ�������D���ˈF�<�@ ~�c-[8��+ܷ�>�".�x�`��<梯�@*\�[��5}M\ʩ�?��Hh�b����p���֍^3j��p+.+�@�~�r���iS\�z��a�ڱN�\�X'0<_��V�X�v�X�_�+J�'��MM	3X����$�F.����5h�q$�x�L��M2���cT���g�lG.B����� �dQR�<<Z;oY�,b�!��[8s�ȶɭɺR��&�����8�K���V�UY���)������Aq�X+4��#{0��n�E#!��y��ږ\5�]���!�^t��H28�_���+�(]�'��\�t;/ygGy;��?"_ܼ��Z�e_���eQ�|X���N���'9����Rc�ON������kC'腆?����Jx�ͳm(�}G�󜇖)գ�cuƇ?�01��5����A�h��uh���x(��<_�U����L�A
�#y�ZY�k|����"rcNH�S�-��O�w��F����EѰ��ա����Zg&5����7�F?��������)�&��[P�?�K��yI�R�`�!�'�E�V! �!i�4$�y|�h����6`3�0�s�S �*?�JHz?�-8�$׊xr.H[8���,)��w��a��A�dq�yչ�w�����:ʿ"X��[1Hm�z��#�n�;��ʱ-�>dJWd�H�����{ dOZ�[Np��<�V�]2���y����?�06��y'?�@ �JEu�����l�E!Z�/H�����t\�.n�RyY�޿3���oUa�oL���bmb������5ZDJ�>��+�h<hW��|��v
L ��rz�tDZCzE��k�K\$ʊ��V�=�р���l	�*nh7pGF���� �H�3��h�[h�@G:�#���C�x�r�:��E����7Z���W���0�^d0Q���y��Q)��կ���p ���l�FMo��%����B��N�~i������k�HR�;�p_+H�%��R��j(�����T/���Ȋ ���1��8�1C��w��U���h��y�8��^���82X��DX*������0j��Ay={
D%o�"�ʍ���(9
� �������4J���(����,��:����M��ih�|U�
�`���U�0���<�<�ff�1����|����J�ŖΒ�l3Rf��P�q� ��	(t&�4(<����o�M�ƕ$L63X���#Mdy&�Te�!H�|�ۜlX�ϻ���Zغ�#v�ū���8a/&6��R|(1w)\G���Qb�3��c�v�VlBK���~yB��Z�dy�ї���[4_��&�؜{�wo:�y�\��d�����]�+��[ď�6��n�\`�ͽS`'�Qs�3"rF�G��O*m�4ٕ8{��&�&b�\���F�CU�>���"3@l|���Qm0��T��R_� X��<��dE����y�f����A�;^4��JP	�������^ E��V�I\�i����y�En�:st24����!��I������ŧa���A��0;*�
���@�NQm��.���4]��]kOEr�~�S���s���v�{����揵��;�gX{1����Z1�'��k��C�� ��%� �F^��`�Kqy ���d��o�!��cU��M�P?�������gӁ>��>D9�V ^Z�F��������,{�"3_CwfU�w�[��$Y��Aɞ�����'+�z�rU�'sn��X�)�@�%������g��(pա�
��:���,̩��}�t�\K;�eT��x�,��A�{�h <�Z�=f\��D��tW9�V�v1!��}�J��7`5�Iw�qi~n�����]�Zl��/O_�QO1ۙ����I\8��=����5��&������w,`K_0��2����(�^��_/�1E�L��xx١�Y�T5�|�]U�"�o�M7���˒ *��ï^�>��e���S����=�G^Dw��T�2VS3�_�(;t�|�����_.�N�$Ͼ5~��+^Y�P:I1��u/��|Dl|��H�W�Rӹ1�����%�ʔ�q�~����a��Ʌ#��L�+�D>
f[\y���pB̫���ہ,�\䵴��qv0��7W]�� �F��+'�WJ����<�;������<�e�fk1(,�TL����F"��׀Ĕ'M綽~_��^��A���r�a�E���F�C!��v�$�c�?d}Q)P�M��2�ǋ�h�h���K*����{݊B����E� K�TNRd��׾d��@�w����X3]�{�>���=R� ����@�]gho��tB�E@��P�=g����ǯ&��<��'�K҄�s���?���)�a���G��=l��a���^?��x
�-��PJH 8��tQ������T̀�7�I��[�����Kʳ%��}�dd���h/���ޏ�f2'cq�sC���Gv��i����4�0�߶r^HS�i\��5��Y��e3 �]�[P�4xB���<��*�ɧ�!�Ͳ|��'f���ڕX1?� L.&}?�P�O����q&:���v=��L��s�~�</;��?�c�c�\;>���?�r���ВL��yK9��M���|�v�vH�}�AmdsL	�t4b��Ϝ ���F'��a��펶��#���yif����p$Q��cSP��
��ʦ����$\@�� 	Qz�%���+E'���� e1
��5��ᄷ���B[�*'�VO�J9����1(J�
�3͚qn�M�:�vm����!��uu%c6��}ѥKiz�E�����.��u9@���G��[06\{�� h9E?F]��]M*W�K�w��KE/:��9���dL�6|��X7�3v�c���"��T����N<���k^f�Q�v۲z<�c�t���Ȃ�q��2R1��k�t�^��l����-҆��讔q��b��T8Z\1eCN�tzզ�h��5G&�9�����8E�$�qNAZ�e`+C$L�}��n�NwQO���~�����]?�5�z����`���PD&����/?k��V�6*�� ����!CPeh���veJa3��ϊ`ϕ*Ldɀ|����%o�6;\6y��B�V�fo��G�(8��@�{"CS��������d�8�$8��$�K��$v�2:�=��1��/6�h)��,�Ϝ S��S��`�oI�:��H�C�,Ek�0do�C�(��ݔ��C{����Q����r)�	��t-�Z�W��u{RR�ld�w�.��	r���r$��� HZ����{77�*
��ngH��[�Or��ʹ�1��RsѠ�j�da.��yd91��#����M�7��f[���?I-G�k�����9s���%�#q�o~��Y�柭��Ռ�	��!�Py��!?=+��ԋ�w��N_B�6p�"cgd���D�Y��..�yRXJ��H=�⟘�x+�H�������Akߋ�.�RB���W�aX�X���@&��@��\RG;��].�4gsz,Ka����z�*�="�u�d�}4u��̌��%�_�bI;FI;�p�v�Ocr�������b��m~J��l0�
��P�6�Q#*=K� 
g	ޥ�E��ʽ���^�L�t�����es���}$�?ZJ���:��(�r��p��Ï�I�"�?y���!W-�uu+bs�����^�G����?̗�w1z&o$�}��R|��V�;�g�5I�����`6\�u.�*MB��*��n �'���y��D��_�2�Y *H�R=�T�Q~��!Y�~�љ�84V�i��u�F�j@��N�H8�+v+c���,�m��)�il4��Y���P_m��&�2P�ہ����6����u��X���K1ί	;
���+��e�46;�ي_��H4]�C2��ę���BS"���1F4�B&�t����/m�l��c�G�8��-�P�����:��M�[��X,�dҪ12��7p� �F�wE0+�c	��F߅�kb��
/~�]���*��H��uo�D�7@�,=+��Ĺ:�Ш�^M��d2��a�K}�W��V��&O�&�}ឤdm���ɽ$�k�6�Z��G�V2���@
 ��:�Ŋ	�%�ڮ8G6y8���U�>��[��(|`\q�q���;�ǧlS���C�S-���ց������e��D%��Te01S�A����(��e�Aw��N��ǢY��a��xYZ�mk�͌0� �H.��CO����,���0Z7��� T�>0�=���oHZq�Й�R�s�/c8��o3ۛ������!e�����DC}�ͩ���]2sx{ʾ&�������B�M����t�XdU2�e٩�J�%�@i+�'h�\0;3gu��!���I��4L�D�����>��z�wA�YM�.��믔½�V��q��=�_b��o�F>h�l�c��Ԅ�'�F�R�TA���AI��"�{�#R��*�����lХ�Ep�'�
s�	�o�ڿ]�y�_�Z�'�����וI9���P�K܅���1Y�����1������`W�VR��T�'��ۻ�*@f��&��W񦎢j��	j����g�ἐ�_7O�35��ޭ/�����S���ۓ�Y}FrBn�l��aE\`��v�9��&��h��й=֪
�����otf]N}^5��a�3�pW�!(�^�����{Pa�c~�c�l�=��>�i�>��-)?����47|I���*,*q�ff6�x�c�NG��T������YȀh���=vdL�rƒX�cs9fJ9@q5�FgT�j�;%�Z��P���`���(���-S�(����wIZ�/��u�	_+hr]5>?dqg�~�;�ل�5#���sIlfQ$�<�u@����i�Y��TS�<��"���H�RL�B>m��fM��U�9�����眽�X��<���$��%�eK��z��� � Z����?��6GQ�'���u�ַ�&.�_Ɏ-�%xB��>�l��6A�B�I���y]X7�/O7z".e鈃&�k��O��n���0n�I� _C�EĿ�a�$A~w�ǽ+�ڻ�Xpl�,����߮�=��nN��**n@�1Ooy%���#�kY`:n"����$zR�n?���`��p_l���(ڗV���e<2���;y�Q�o�t=��(���@ʃ^���� �kN��tr�A�>�XH�&Ir�^M@�Zj]����Aw�Ӹgf��@L;8O���5�������Z_��9���
c1U/+���"3�!�P��U&�j�����^�71�}���Z��gqP|O��h��D/"U���?��MV�b�����p��v[Β_�D`���D����/~C��2�����(�6�#���eю9��d�;����"��|V�46W�Q"�� MJ���Pc�t�Ç��(]?I/�P�Ag�
�����=�������ї�Wx6�_`����J7������[�|Y��4|8|]�ҳ�̚�Bt�Q��2X�H��}�Wٿ�:1��G�E�$CZ��L.��e9Śϯ0�RY�_�^fڧo7ළ�X5zI�qɪ���3yw��#QN��T�2`�����H�����ׇ	91�w'��ÐѻX<�x�6�ʠ˚Co�i*2�%i�!�V���X�C��n�P:��VG���%���-9_"�h~�H���#�H��p�I��[d{�#9m
�D�o;�R�z �x!U4�z��D7oୃ�x3�#R�͏(�����:.��'t�@mGz���q�����w�EA� ��M����T��.p|
Ѫ�kx_!E�������n�2.;�J��w���tℱ�����;�En?� ��7PB�ӈ����}�%`�3�t��1���F�{e�ە�z
��^�V�v�|~a��%Oݝ.�� F��?��b"�����e���E�����w��1�-��V��*��[.0q��&�8��HS����"��,�(¿f�UɅ��Lۛ�T�p������M�����dl�ϪZ�y�j2F��'�=bKX���6pn���u�K?�;5��Z�C�%Tp�$3�o[���.h�vxp`��(�Tq	����f�����sZ/��?,���cX����Hܶ�o�	����|��U�Q�dJ� J-��Aه4�	I��τB?���"�ELGak�r��u�5�Z��g��9/�e)뒈"ť!,���yugB\r���sa:�
_�7�_W�.���=d���_����t��<�����gY*K�6���f�m�-F3��P0�8qe�(yX��3x��.�S������?���J*[�#�8�۸r�?��`O}p��[��9-���3�,
),3hRP�<r".^z�^�#�a^T�SL)��y����(m@+�AUA�^d�1�c͉�73�.tS�f
��f�qVw��8K��E�	��Z�*O�Y����2� tF�0Pu�Y����ᾷ>�
T���.�=�]�%>o�X���'I����^�:
��
Ե�8"F�h;w�E8߯��Fl'��;�(_>|�|{�0�Z��q8�"���E�L8�s�Hs�b�$Y,{Tl�%���F�LϏ5H=�1��`p(+001�-7�<�a:Ѱ�����H��C�d�t'��� *�$FWX�&�ȿ�F���BAg����w"�5���֖� ��M�u�=����<yY��K�  !�7k���-y.>Q�hi��'����X�0����}�[p(�,b�c��
�>��d����&�yĊ�Z���H�=!�ʡu1��į��E�s!�T���K��#�uj�L�"-�z���ZoϢ<��N=�nP��r�k�d��1oS���<�f;��#K���x6i�xNxw����O�Ө����h����l��M9^�7T{b`�5�ʵD}:�]bK}�S�
<�04��͹� ���X#��8�Ӻ�-�'��/K'���F�V�P�����cpjj�,�!yu���,r$���]ǚO0�ԑr��|	2p�1�V,D�l���f�{��r�-6k�*�c���8�+J;�f|iw}���h+�;%n�9u��R����4q��F�ްm��":#�ͷF��W=�f�\�t�S�r��m��B�R�7�>�� !�*�)��?@(يd܉r&\>itc�\|�hT�O@��p�.��������*��Z�Ed6-��pܺ��~����+��-j�އ��qF@��{�Q6�΢F�Ɯ��f|ɍY��$�ԛ0�i�S:x�E����v1���K}����@h�"����9,4�oh�H\�a���������Lc���s�i�$l�Ǯt{��"jv�
0g��I~�*ut�+��hO?`�T6U�U��D!�Q�HC���N�Q��,�&ߗA�1`�+~S��m�L��T��G9�<�ۧ���o`�5�}�o��]��Ӵ^/5���d�N���� tR�p.�Vǳ�~�P�$�ͽ�(aP�RL>wgف��C���֬��湺-A�ո�������E�K���{oE��<��9�T���o?6^���N	@�7oL+��ְ{c=��%I��������M��!��
f��Z8(��h�N�̛�u�F1I݃E|�ïw];nx�Tl
���͝pf L�9ǵ�W1���e'UCE/"A;qy3��ؾ�|9��V�~O���[�-9��m��W�"�6�E-z�Hh���Uo��Wj�dV��M�4��Î��6�"ӂ�ғ	A�@S��絛�b1��'���m����(IK�b����G5X�-�^M[�>5�����-sh����� �~n�z�_��[<���C;͚��5����E>��cú��V� ��L�����ZxX�#]BE��4*��$�Z?��słr�\�����G�Z����_�N������y�� ^o���Ċ�9�4�����5����T��@��U���)ո4f�U����G{4�K���X�9Gb	<�A�/$yy���ʱ;���j��=t⥖�G�Q,J鈉�^?C���A�����H�f�}��4R{7 1`ʨ��ik��NB��>Y�g�#?ƚ���<���D+�(���N�"Nh$?O�Y�4�| �F��A������{��Z�as�+�0�*�k����փ���>Z���Bΐ\�i�I�����PU�Ѝi�lV��!H���� ��	D@�z%����D�V:�2��h{XȮ���GYr"�H���c��H���xǌCL��) ���Y��(�sk�̸	�{�ȌN�K�@5CS�N����Z��
�;�#8f>ZTM�Yhl*�A��
�*�!.V�+�1a=d%� ��	�8�J���%dn'�����Ϸ�����!8?��0�W��;6q�S�Wd�B+������ 9{�V��ĭ���(Ď�u��ν����1�L�]�e�2!-Mk��v]Z��0/�=���&޳���]�{��>�I�ھ@�y�0-dG(?�!�¾uܛ�bh1���_���Ps�B).��^6{`��+;������/`j���\�8J|�f�h�;wJrŅ�v�0�;�`����~�E�9�;���������tn��:`� 6��.v�󍀪�}�e;�����1,r��a%�����9,�Z�������t���{3{c)���0N$k���SM�n�_N^�u�o�1$^ ��p�g�X�hy�|����nʋѹc(�i(l�#���w���' ����}���x��6��7��PUӞLg��o��Ҽ��j߆n<���:�[�8�v�Y�*%D>WT��n)����>>�z���^�h�$7bIO����b��x��iƆ�=�k�Q��G,�.�J�>�a�t����-G�k3�?�/m'a��=<�YV��]������Q6݄������U��)�q��o�c#`�y���Kk_Ik��)+ׅ��?���J0��]mP\,-}RH?���g0:���$�5�6�v� ן4��IssQ�J5�Ac�mN�'=�	�*I3�m�O,D��b���%�&}�

P� �\���%ծҴd�1�q�\`��r��q�^ο<����ȭ����'$2�-nѲ�u���d
z��k�����Ĉ��ո '�t�;.���4.+ɚ�~gd�Xb�4����*���}'��f��sMV���4MD��s��e���\8�TR�	 ������fd�V��AM��$���U� �~��?/7sȺ�Ч�D$������l)m�<��Sb�T�;*���L�|s���uh햋ݤ��M��fK;��M?�3�X�ą��r.�<�8���՟B��;���x-��tsܟ:j�FV赏���ɂ�J����uv%�3���R����M^�S�mn,��w�����&����pmd-��1v,a+̹؀����3��,�J�K�5u ���3�+�h�աN�_MIA����j���!�c�F�ʖ�i�(�J��o��Á�'J�������@�#\5]�v���%t����I&��
а��.���>i	�bB���G�C���}_[��G��	�*��B5�+���j"q;R�hOф�4�W���]�"l���m"�{�V5>7AD�*�y��)��H$t�xf�k��A����ps�� �	���+����Y3�#8BO��'�:�9+�O�����y��+2�fF�]L������!K���GZHK��o3�����罹�5K���g�5�W�D6]���Q4�����N��VJ��O�<��1y���&4J�E�e�_����l��B �n'��'���m�P�&�bEu��-��[|<v ��W��[kp���_������-�y.0k쓃�#�)�"�x�|���D+UG�V�#��'B͵NAi�������%�}�;{d�{�R�#�gU;@��9z}�ݸs!�Y����s�C� <��� Z�w�.*�T\b�H������1x�|���z��l�mj�^�q/
1��nm��n�(�oa&xMu���s�/F�����g4�+��~�H�c�j,�ɄL[�H"�֪�/����X蟽�U�
���YY����C��9L�|�ު�D����ʳ�����(2 �.ȺW��`��-��BD�o4�a�V%�NZǼz�ԛ+x��|f����o����p�$,��1�I�R�;ξt�'� ȱk'���?G��d��"ǧ�&sF��Jd%K��4ӽ�B�ճ�At���?졜"A1��臘��%���tb������T#9Ua�Xw4CV�,�聤Gb:d��u�CC��5��3*�i��@��*��*���8h;��M���hɒu9t簉b� ��v�����<f�*n��&�䐌G�$�=l��ǅ�]gUG���mo�<%�� �l>,8��ҁ�9��i4ӎ����E�(VxT��s���X�ŕEUg�`�2A�צ�=�C~TN�b߳�q]��~M)���Ex��*�D���P�b�_ǈeZ�P��5閟Aߛ��|��X��
��ғ��!�T6x��9tHÉ���IRF<+�u���B�Ƌ��E�rܯ.�Y��X�����]��>dy	�� �H)WQ�r&�Xdc��"P�)��';���5y�G��ijѬ;�Z��eoI��8�=��������-��r�\+�&49�4m~h !=ā[Y+R�뿷�]���33ŭY�%�z�x>V���E.�~Wy�B�fF�����y�z�."�\���������ǔ��A�K?��z�x��4���6��K��:�[J��]�jU��6�|a�-�"龇���
1��6��k@r�4�ք���h8��[������Cr/ķR&��@q�bVa���#���6y�ʕ�D��\qZ�Q�����E��� *=$Ak���Hr��h!�����n)�`���{�ȴ��a\��y���JI�:���8dvhAOz��<4�;3ㆩ2�8�k�Z�0�)�0���-}�H�O~Z�"k�z�KΨ�ñ(%�*-�1���H�� 0���eɌ�Y�?-0��'"L�G�}]]�
�
�:�$0���hI+����bm/3���=�{`Dh����/7�R���[���l�������\U+&_դ��ë���rHc�����
Ä���7��(;��򸱧��2���a�r�l)*�b��������q�$���E�w[Kr�m[�ਲ਼d)-��1�hޓ�G��oEA�`�Tˑ�S'	
��x�lY[�~�?�����?���B�ԩ��ʶi �?�#\[e��@�CA���`f��E��7��dDWƧ�E	})���>c�r�*G)��7uN���v��P�զ{����`�R&A�=�V像��]�Ne7�k�R-@ ��e�����X���ܽ@ص���H� |�!�PK�x��ʅ��L?h|��J�����Ս��A�g+���$��
��ч�T��ݖ=��"V���ڢM';F��2�� �MU16�W9������V�3�P����`ZB�����DEo%ş8�?i����vT�p'X�O�u�Q�x�ӳj���r!EQ ��Ѳ}=��  ���Q�s�~ĚQ� ��^���;��{�^�˿�iF�m�F%ɠ`UE���K�G��W��B�;��ق�jK	���4ƚ~�����R�>�4L�)D	�I����5V�&�"V�ƀ�o�~������Q�h�7;P1�f����z��z��|l�
��"`�V�;,l�o�x�3�i�'���N(��V�dR�8�C�J,���=�u�����ZBҵYqH�X߃$н$�P�"�b�&��	���bKjA��6b�c(���٭�űeo򥱦�X��2��I��X�ڭa�ɂ���[�DiJ`厰.0yc����}�I��3YQ�\属]�#LGʇ��QX����(Z�GY��f�sT���q��ʈ5�V��!e� �<�wwKFTؙ��	=�v��Y�	y���(qEń�l��x��ps;S�Z�}d�H�	l��������_~��DSљv��9�6n��>�Yڨjsҗ���!���j�s��C��=��C�Zde��5���6.���ƈ��
S�HێB�� >����e$
c��9x��#�m�us�l+x�����})��ݚ`Ұ|�GP ����� b�%�9]K����D';!˔�����!A�[�^��A?Ix/G�e�o�Ƚo�,��òT����Y��d�b��Թ�;��zrҤ}/LV��Cѿ���C>Q8�H���\M���5nJ��S,O��=^dS�B�=�T�����&�ڨK*}V3ǧ	r5��sbp�fEf�b�t)PA�(���
/��E���?Ø߆�&�Y�0�VX��Zv��nV|`3�_-���ή�ؖ��/���(��˹�A�X�b;K��W�c��hޭ����#�Ø6u��di��O%���N��X��*o�(����Yq�����4z�l����׾��L���#�`Q��E�LSP̺���,����>���g�������ֵ� �F@21�����:k)�TM�'���:*Lȷ_��))��暛�6�c���u���?��&��;jSW]y�v$%��Q�1�I2��N���nA=�/�1s_�m��X	Qp��o��0K|�BF����+PA>MD*cnC�Y�����g�h���~.�t�}a�®3�!���j� �����g����8T��gzF�}�	0~�{��$�C�>�9}#wa	�����g�HRv-�\D�!�&�c(���|%�Cr'3��F���ϛ}�3��S�xAɝ�vRDk�`)#��B�T�J�)q�my#_����I��^,��;=�M��H�q�D\�h�C����tB�%Յ��n�Fu{*�cYN��2�>�!�%ҳf�P�xu��þ�~D+��t�m,��rwJ��>��1)v��3�5�u�n-�WjE�"��m���������Q~!��U�B�k��8���|4��:�CYX�u&����Y�pk��I�<��-�y�n��-��-B{�f�?+ʺ�,���{3	f'9�{H�ލK,�"�ҁZ܁�#���Zl��K���B��<	�UPVe�Z�>6�w��r��!s���5w�}v#e���ߩE�Tw�p���W�cD �||��ѥ��F �(��M�<Y��J��?����Y�C��]\TL��9����FR?vn�&�,DQ.�C !�����P��$�&FK9Yvō����CNQ���Z�t]Ϯ�5w��Y�!���d
1���E7�uJ����� JiJ:���Ҩ�A�������xOd%����ܟ�At�-�)�6j����\s�
o=��1���%��T��L���8�4ɖ���jRҍ�y�7
NK˧�7���U�e4L]*�~f$L��<��R\	��"�K	:�d��Xx���|�����7�i�� ��&GN���{�?��>6��厮D[����h�r��;*��d|_&^��M��T���G������=_���z��xd��.K�A��I�QK�h��o�2�����
�7'flWyj�:t�C�h�PO��
����(sz��	
�\ӎ�wRe<A+��(�� ���,
��&�݁�5�ҫ���q����1 �C6����M9N��iSBZ8��P����V8x� W�M{6��b�f�'k�;/��u�@�0��?9fyj�t="�Gj�{4��Qd ���œ�}��Q�sh��qPX���w��mB�9�Y?�&n�x�*�c4�����w�YJ9w���m.e~x� ���'��{u��y�|��[��y1 ��*���x�Jq7c~h�`."�����M+v�������Ve��m"���ź�	7��L��8�	��m �{�р-wgαNN�wI&�����@Z���f��6�P�n�;ʢ�_}�4�bH�X��Un1�L%0!@�DZ�����{�2$[G���q֕��BK��-=��� ��o5����j9�-\]�mԳ�c��ksl��d0����4��ac����u��%-���P���k��1�x�N���|ǔ{��
��C�Y�b��t�;�x3���8�p��b� �Bm�ap=x�� :��%�B�|4�1)�%����]r��P���ߡ�[.DP��(^N�����w!�2B�|񂊭� ʇ�H����m��83
�jl`�QF+�96��)���x�p�����&_����V�v�ȧ�H�1+aH%'S3�I�ͅjL�S&biN5�2SOD8?Hw!��0��@	$�QjJ��V1]w�+�ǜ}��ѭ��\���/��t1(��mh��U�uUA29�C{.=�1���e?��<*�"���W�m�M9�I�
䂀nt��4�����w@\7�@���Ix��od�����`����x��[�#	�З�n^o��~N�ba�w]�����S\nI�n፨8�.�S\�hM�p���9���[��P1�V��;�*��8��3ք�)c���:�s��E3������07���[�.��b�����/	ZQ���b��U���*���X!}��/�� �����;�}
������p�#7OY���d�0����k�w<�s�f}`��?�����!�.]�3������|8����BI�H�[w�O !�JL��ɒ뎑����/o��r���@wUl�@�wsCaw�j�
�e��d�q�l�E�׵|9��tCQ��Ў���EjK��İ��l�Ԅ�#�nT�J��g���mx;3�U�O��]@ecA	�&SLq)�S�,`X���Ch3��kB�_���z��H_�LR���d�@<� 1:v��F�Oka}�t�+��sB����*�E�g8n/έoܧ��-K{�$d?���qh��6?�o��踐C�p���@�7$��������(������M�R��w0,"�	F+���Vo9F���rs��` S1�sąJ��rGR�>�D��ے�,A�^Y��D՘���E�Q܋�"��ށaʀFW�{&������.��j�DI��%^y��/�
k^@��:Vil�/��f�b8�
�p�2�;H���[���0�����[��h�K9��a���ES/���b;߁��ףp�:�K�F/Ў�$ �Jr�	�VNޙ�}�4��Fp1��A�!�HS/��=��P%P0�����+��*����� ����*q
-�U�;�d�窪��·.����:�B����� ��<̜�L���H�&N�k]�������H��^�kY���b�]r�͇D-P�1��.7��W@Qo�v�a7;�U[a��7��3<���&v߇c�.� ᣢfʃ#�X
c�����D��	���?bu��vm��`�X[:���ؾ��ORO�#j�T����MT�߀� \�g!��C����x�2j��Dbe��1��ymƪ�<tčs��Y6�~X(�P�v[��qsq*Y���G{K�Ls4��zX��%�^�56[4�!m+�&s�M�f��P��3r�;������
�3٭&� a�g߷���+	�i�����R۟�8#G�`i�@��Hu���a-%g�W��|�J� q�S�#��kW��3��J��:���Ur��ufg��vHq@<%�[����֨6�irn��BG�W�Z����$��d�kT�_���M�M�pE��h��4ԬS�Ta�=���<Ig��yk��� �WqR���@���)N�c;�6�א�3�0�]���̋�lxt{C"�En��j�a�":o.г~ת/��J�R�R��>���*`���O�/qOb9j���C�vڥɪ���ؚ���8�7_��,�~���]Ĺ�)���9$�w�O����������H����	f�<[J���v��6y�����̻D?�0��3I�UI������/O&B�����.؇k �d󞣹
�Ugd{�ϣ�(�W@�cbVC�9|H_QbQK����	-���A��k��b����gw v\.#��B� m6�_�XT]bm����p�9e�Si}��s�W����ZSĴ��K�cv���:���E~�A@��va��Ӌ���iΡS�1�`4rDO�!�D�2c�>�s���J���E�p��㿳ko��I#R]3.Z���������w�<�����{R��}<�n�/B���֞-�AH������������g�~n�i�a+\D��֖�L�$o���&9m<��.��;�A����9a9�J��V;)hI���p��	KSm�!��pj�fgT��ANVfe�,�Q���B�!�4�\^�����h���?��G�:oӀ��v���j��|�U`��'G��>�NB�(���*�ב2n_X&40_>�d�xޗ>ep��?(��� �}��� �9߄�q�IZ���������<W��ub���5=HH�t�"C:�����0���2q��/�v��B.��1���.��������	⣋�+�̅���GJ����5�+�4����v%����Iv�W���S�^9��# c,�^e��OD�p}0�y���(3޿��U*��|�B5]n���bpv�՟��r��Q_.��\pj��.������U�Q�Ar �/	a�I%=��p�'��Xm�Y�}&PƽJE�-O�NrƵ_�~�6�1P�K�!���/�X�PD��E�ޚ�4K$�7KNr���Ek}�$���~G�e�)��Q�C+�p���w'_W+�"��a$�m���^?������@����~]{�~{>�f4��)z�jl�fIs ���4 2霷-���܂O�$#i�ߟ���%���ä��:�ᱛvƣ�~�1%~إ�_Q�I�~/�/g�CA�Z�u���#K񁋫"�"����h|��l�閩�"�!c���?K�ݜ�i���+���1��l�@�kf��)�*�kH�3G@OS;��]���7����>�~Fy�a
.�\��f��u-x���OaG�Ժ�0�_�zV����
��}=*���L�:Uwr�@#��ȴ= �xv����¨O�Z�'���]���}�p�p�Y�t�?k�su(6�R�����̀7�2ڥ���h��ʮ1
{��j�2�赩jR w�<e�D�v�Z'r,뚀3j`�w���&Εq͙Yixz
R�z�0�/��dF�G`_�ɔ�\t���R����,�:$}��n7��6o�{���p���o�?��h��~
��+��Sn�x(edp����>����j���%*��(�1<�������'ع���ud	�f�Q���B��� |4�g���yGT��,��Ą/��g��kuJf5Iy��I*2<��͠-M��-�1V��J��'�|�2	Uku,%E��ՔS�S}�V��He���Ԯ�lqs��ȿX(��a�N�A7}K2�k�y�f����O&��}V_����(1�6*jk����=�����XX�%$�2S$�2XLae<�,60ԫ��N��ҰPN�����O9�Sbԭ����4Օ�h}�;��!�_�F��O.qõ=v��Η���TȻ�&��阹V��/���@w%�~!2��P��/�d4)�QXo�JjVV��&���:����E���l��=�����=Qh%(JLղQ�$�ð=�R784�	V{�R���*�;���Ăk�!���Нd����hE��f���p�;��9@���NųA����c�\�̲�{�jDZ5��<��65ɐ�M�Y��Rs5�w����
��9���N�#�3�npp��|Zm=tz{+�z� !�$ Wp��И$I+[�ξ���,]g`�A8f������6���X<"������?O����[SC�"a{'�e�,Hӡ����ʶB�bT3�N�z��C���V
�q�`R����$8�<XIRRU��=3�����TF|��D�}=Ck�mE"�eY�:�ϴ� �	"�a�۳r\�" 4��&��Aء�#���]����"v&Nct@�7�/NoF�8�/�M�z���m����v
����*N���_<8�V���kr����P� `M��\�PҚ��غU��D5NU0/�(��G��hr � ��~Bt���l 7�'tA��X8Xx��տNk��1N�-ɮ�#;l�������1x��֮w�\ff�k�"Q�������K<3S<b������,?L {���g��qua� ޤ��.+�Xk;�NG(c(���ځ���<�59��E)B���j�����_��%.�JBA�&r-^/ǌ�wPY��I��¨���MF�a;�p���O���!r���?C�p2�~#+Q`��鹩1�%)���oay,��J�0�����Zh]Cd&rꮅ��^�S�]瘅�eA$��E�%�Y��`R��!�|�8v�^%���`��fu��MR�	ۅ<No\O��|� M|]R��ȶ(�����e�[	��#P�7���Ul�7�j��S��t��V�q�aϟ[�(G�W��̗5�_�$V|^Zd���N����Z"v&~�@�b_ď����c�R��J�ac����x����|������8i�͏(�Ÿ��7�̧U�eW����+��K��=j�L��&x��5`�Li\6{��&;R�g�����~�Ug�*�����O;�D뒤G3�܂��{Y��{E:$�}ޫ˨���K0�v�^�\���X����kӏq��
vBx]�\��ks~�b��F�0�# ?R��eg�|���*��9��y-��d�UK�.�x�F'1+��
x��5����#��
B���2��w��ȉ�~�񠽫'�G��#��l�
V���e	����tmM��J���e�RN�'��j"ȣ r|;�c��k�d���˂A�Mc<a���$+=>/9��:g+f�o��ʹ�!�R���К�е���'����"�Zv3����=Ҥ���%?�cGq*S�L8����< �6�\��un������+�0Ҷ�I�:8F��
k����G�\�����,c�i�v� P(�~�7��+�Ca�1S���̶���Fs��bQ�v?�\����-R?5��ե�{��	���'Ś����9�Z�%׏m�
���n�X|W�M�Կ	AA��4�̲����Vi"�>�Tk� �B��xZV-G�d���B%�-5�]r�f���g��$����+z�83.-mf�c�� �a��]/�A �YK �f��ZT	)�Ts�e�e���Y�=�k}D4M�w�j�H��}*F�q���"֝?M��ze'10�7ӔQ��Gy�=��&�]��<�7Ϳ)a��%���w�v=\�J����vJi��5��.^�~��$���9�&��r�q�tڽ�˰�;5�܀Q��,NIN��g{���qnx+�
�c\� �8�,dh�7%"��f���oW	V�,�7>�w�p�GxL���5�+�Čd� ��p&s|���A�g��X�ÿW!��exB�W�W�"D�? ��kY���t�j��b��sw�=$o�椦$d�H�̢�ld��gk:3�{8ͱU+:.T9?���%�D�%/nft��+��-���4�����	Cy殯��t}�:�Iv�c��%ET&�B���-{0� gɃR[���l��_��a���lK�;݉�}�ȣ��.���&�^`dy���R�$`�������A�
�Ľ���r�
ZN�h��ע��#���,����o�`#[��ZG�����C�/�P�� g+�]���R�ċu��dj���C"�ۘ}��;Nj!p�Z�{�{�ј4�Z��-C!����f�4{��uæ�]{����xIϒ�&����JL�wΣ��ښ��Q��Ux� S��z1w��^��Sϣ�e� ��h�LD�®5���Z�?�L&��1{�P<V������}�![��Y��4���=������냷��@�ԏ�>��:|�/��5�t ����� �;b( ��R�������&_
'��]g�6�	��v��-��Ka�P 0�	��u����Q��@zJa�`5���ɮ����D3��aIO�p@Xs�h�~|OQyN��m�Ph pO�v�����}\ r��<Na%�u���v�������5�HɖR�R[ļ<aC���ВU����M���
�<A2\Fk�u\�T8�06�>�X:?�Z�����h��t�	�b�E!��V��of�������tOe�>���Y�]D��v��R~LZ�E�����k�ڔs��u*�ѴE�,8{9�VM�f�h�P��'h]?��aB�s�Q����<�����+�ŕ�[��<O�pR0f�LH"SFyZ�*��2{,h�TW3�ȼ)��ayŲ�Ǫ���Ϋm��o�'�-��5��)�9i���������8Zm�K6n��j[�w��C���E>�)���v0 �#�٨_�� .�.e0e��I�̝[b�&g!��ݮ�W:�5���,��y˅×����U.��Yla���5�zR��Qe"s{Cn���_̩6�V\G>-�^�fX�3�:��c��l�n������[�"|�m�]B��	*@�G�P=�+�ٮ�A���@��5���BK/D����3�]��+�8�A�b����*�j:���nfTa�����s�φE٨-��p�]��꧐
�Xc����8R��>���N�"������p,�[���2�3�x�嵅|�*�ߵз�"�x�U��ò�֭YM.mMK'9B\A,�
&����v'۸&�qF�΄�gA%��$�tn��1�/.�N�yu�|�O��H���wZ��c��
����*^&̬%�FB�%"�LM�I�g�X�S�c��E�����{�|L'���>[Bͅ>c��3Az��ߔ�Sd/�S�yI�NPI��0��5�~�Y\��+�?(���.X��)/C9=R(Ke�����P$i�o�9p7[��a��B�S��%����������E
Kn:�޴{Hk^V;��]�u�\�bǢC�Y�&pz/�p�M��z3n���^jI(�|x�
�6A�f�O�Щ��h$�"|�+�d���j���b5���v���%��ӧU0��j�.���&�Q�y��_��� G��E�`/Z֩�p�^@ֳ�ET��A�³� +ިl�MC�Ѩ���/g��u;��wN��2����%�<	��܆sA���C��l��t�Es�Bvy?�w�u�T�.ǎ�D�)�*��k�?�<�����~r����j�a�W�*���M^�\A���G��7Ӓ�^���3�]|����ı	^e)m3O86�wk�8��d�4Gֺ���ûS���k:��I�-T	��,�Q�i1ā@Y�KrQ� �A'˄`�]��z�]I��m;�;�ـ�f?l�i�hx+`+҆�ue<����,c��"����Oo�Ԗ�|p�^1"�ځ�CU�|���vUipu�j����c��0 �:%9c�:C�d�y���\
������	����w=�^Z�.��P�Y�M�]r!߼�zp�W	�˕�E��:�UfX��YL��Xu�r��3�J�"%0y�Z���b���u���ٴ��x�V�(>T�}D���_�#���P��ؚQv�r��V�L
ꐑj�#�re��4l�ψ���zp�_*&�-'_@av���}�=�F��� ֘+�d=\��0�������X1�[�B���x��~Bc=�ր�:g89�e��rd��v MJ0��ht37ÕZ�fC{0^��[��KT�g6�ܕ��������J3	#�[�p�Wy1n��a�Cf0t
���%��0շ�b��h���/N��F����Sb�r�������48B��|�/b艑Bon���2�נu���6�Ү�9��ql�X�����3�& Qui�s1�
���1J���g[�.���ݙ������0�Y��%/&���a�f�8�j����>�P�4
&4x��l�Yf�~"/��L(r� &�䴍}��ߵ����z�K.C�7Ȩ��8��\�F����[��_��(f#l�aO�qU{)�&�U�$��R��u�Y#3f`,|������f`2$^��r�F�vE�r���tq ����S����WVC�N\�q0�/���(W�W��3e��~���Z<���G��y�9�cYN(��/�ɝTj��U��p���]��?��|�WuX�|�)���д���XZmY���o�>���4R�-k��$
���A�:��PQ�GY�t_��k0��#�y$b�G��5 ����-/�6{<5�Fq�8�/L!��w�O�L��)?f�[�����X�3��Xm+�H�E��b�-�$���z�~�V���})�q��8�T^�s0֌��$Z��Pl1�S}/6��ݐ���s�(��#�~�Q�,؜ǺJv�ŷ�t�{!uwTx�*?dJ�K!GpRa�컬SS�w~�b���wm	`4�d�."���O��z���S�׉BI��wud�;��
���h{��\�ᩥ������3,H&�U�Ǟե�(��AG�>;�Q]u���E^aAB
o��sF�*�P�B�{��z�(�M8p�{յ9�|<Ҹt$ٹ+~T�tp�0_�T���p��!I��j}�?�* t_y�����Y��/���Y}�h<H�#���� 3�;�Y?8pւ�h"p7��!�W�R�/�� 2xR̈́�!��Ay��*_���=�]�m���`?�`1^h����W�������8LYZ҅�Ln|������]+���������Y�=��ܔ���X�1�Ym�on����5�_��P�.vd���5���oVu	��՜d��"��c�GL��T!L��˘�+�ZW*W��0�Ķ7X��੭>:�L�NZv�Q�6�`�H�`p�Z��&/��L�{�-�9B����L�!�����y>������2��{�k�~���Л��!�t���'�+sh��~^�6V�
Ɏ(�(�|�2��z��)�5['ƣ^�L� �������:�Cnp?r�� ��+�B4PJ�Ȏ��|�^0e�ٳJe�T����j����C�6�o��zy_)�B�?���E����|!�?������@坦O�/!fzq��2���Sjv�7D11�G�>�g�-1F[ c��Q���?�%]�ٔś��1CE޻����$?�Y6-�0���CВ��f��W��$#�W�$m{�O#d�%q��J�9�.��6�����\���N1?{,��2j���گ�Ɏԋ�D�.]/�� ��Ѝs9ǹ����x���U�Z�Dt��9s���@޺�9	�t��ڱ:Cr&G�D�V�х�RZԙOV�J�dh��\��tnB����1��vp�ړ%�
���v�<�k�M5M�,^�I�����h�=D �ٽ��,mbja�hj��Ɣ�6�fU�u�y��=��@�B�G
Se�i��t"���05p��(@��H�R�(oj�G��0����� DVm8a�;)v��"xO�#4E�܏X��񔃨"u����P2e���\\2��Q@����rU'6q�I�$����l	"�� m���Gp.w	���1K��7e�E��뾼�[L�龍�88�:���p��ژ�`:+�]بI�M�s�%�[G��#��j�iNg�f��gJ��u�ߞ�P�$���1�iC�<��.G,n�r�d��Ȫ�N\f��/ZG�|J�*����F��r,�����'��V=�i�ՒR�m��m^Z���nz;l��w�ƽ75{���
o+���絲)or�`G�[�k����eӤ�� ;��S-�V��6t6������W"�LR�-�r�Xg���M�ޅ1��,�C��� ���*�|J�������f��c�*N���d H�Wf#CUm���3�� �(�{ZY1L��ѐ��+L��5f�X	X�,���h"Aoغ�L����=aI�c�78����[:8['����s�%]ty��H�ۃ�sQT
���;��$}-j�|�.Aw`�$�{=�ސ�d
�5KZ�*5�|�HC&gsN��4�c�K���Ѻ�w�oK�<4Z���?�6����`
H̫qJ�?v~�J+$�1���ig��,��X'����9�ʯ=�3���I�yq�J�Dஶ��@��UZ��.��T��LP��j!�9n�^\��.����C��,cƍXG�2��)tFG�C�Qk2~���^p �~#F�uݠ�g���"m��1X�No�;0��V5��o&y`i�p"�a�нT�[�FpI�M0�����5��*	H�G�� �ʩ��s/s�������4Ny�0�Ω��

	Z�O��K��fn�n�N�S؞t=����$�Op*��ƥ
ɳF ����U�Q��3�J��7�nꌼג��f"�2:*O�Ш�G�k���ˏ��S�В�i�-�*�zo�Dk)�� �
Px�Q���E��"�����pvp;�_����,|���0Y�����# �5�n�!��H0�w�2>�U�,�����8܆��.2�%�|$D�N��Q�'���R=;� ?��44#�>V��ۮ��MFz����m�{�Ţ�Iٜ���+���=�L�-�����p\cz.�rF�L�� ��3��Qϕ��DDxĠ�R4n�Uc�]݄�6A2/�]��Q�L�1���d6�X
���Ըݳ�6�v��3�D��p�������
n�	.�H�Г5�;F#i\4��k1il��Y>��G�\�Y�gg�%w)��٢�d�
��.�Oʾi[��t�P�ϔ�tį�W8��̱~��\��䒈���A�3�j�量������2��))�T�ԓD@;X�2�lw��� ��^�����.ԩ���� �z�Z���H�^24�~4{��t�<�z����tI�rg|�#���;a2bV$���C	6XGvb�/�T��1d]�Q���i"�N�����O��,���Xg
��#u*���>����Jv�w���mw\����C����+b7ʮZJ#�_CY��C����g����UX�U)�� +Y$	o-A׿auo��"��K�Ħpe��Y��N��8�/7�Nr�o�4�匀ʁu���
�܋���� ��
�k��9������h�f����&�ڍ�Ŝ�n�4Tq<Ap=��:òDp*ݎp���`�8"�3�mk�o�dW���em,�Qꐔxi}� ���J�_G�T����6&D/��{��55��?)>'_�66�#lF4tl�A[�	��?���a-�*��j(;b��Lܓ��.�d���w�Xv7FԪ珹�k]��x�n�z��(,�@�̈r �?����ڌ����I)?�D�]?Pq0��H�S�3z��v���&���v�	3��*�$ukR��Ak��A�dǳGv�!V{�0���r�ʟ�/�gt�pa��t����{�!w�d-����h8�IQ������HfG,+P�)�n�w�=�P��e����W���J�"D�Ə���ǅ�)�F�&o�m8���i�o��o�Qs]�y�К!�� Zo��I?�7H~-r�c����Qq߾\!n^�E�ڏ<2z��J��c�f��j-jl)7�=���MJ]�Ƹ3�am'�����P0�䲖_0�(���ཾ�p�ud�Sm��V��[�Dx�v<(=v��67w�Y�Л�����]X�%�����~ _`�>j�����u��1{��)-�}pR���u4s���%�*�@�m��H|�����A��]��
�����D��O��� M]��/[6�T�<��YcpX�ۜ��T�&��;���P�vX`#�����a��zq�|��+)�2M�'$�qc��ئ_za�c'�-�yϋ�y����!�i�G˽�.-�@�j-���r)�br�D�y�\��}���8�"^ƭD�}�ch��2�nR���8��ё4~��]θ\k�[��¯��|螊��p�iW«�Hpk%�
Uu���Fk���di���`<���1��'�������4�aQ��>3���%���Kdݓ&�$��JV�l_����a�A�w`kfoCX3�y��0�K;܃�9�H.��_�4\���̾}�� ~C�V�;����u���O.�Ƞ���/>�f����3��{��[Fr� �b�#қ����R�×�u5�@w�3&}�g�C8�z��uϲm��Խ�[{+�\+2��� ��31�w��D!�"���Q���j͋1�%��t�&���a�M!>H+������H~��J).�AC��k�D�¯�jAT���4L�tNz��r$ ��Ir�,:?YU�,���=�p��ν{���S�������`��C�27&�ı���}s"h<v���{�F���\��~%RM	ӕ(�3	�^/����x��Gk�q��ϔ��~��@m ��$dR\7:�ъ "��,2�h?��+�6UD�:���<�{�� ��y�n�4<�i>�#[�}0��Uu�#�]�)?����ѯkO��i" cD�'�������ؾp�Ng�$�"����LB�9)���3{��ș���9P;Z=J��մ�	�y�i���cc՛��$��"���mulN9�*�w�UG��@D9�Ck�d%�

���� �pg8.�Q$�RN@���j-uVh(r����PM�#��_z�����?��Y��:��qP�Xe���l�*!���RV�<V3th��r;y�)doѐ~��b�m�K���5�/�{�}��Tژ���t����JY�Rs!"�;!���\	2H�� "P#�O�Ϸ����(�f �mp�����.�V3�]��T��v�f/8BB�Z �}�	X��}c:"B��b��lG��v��{T�h�녲�v��ksg�ɛ�Ip=�"�l�������xc�ǩ�� ��}b@1B����N�q�'�j������� V�-u��'z��,gս��O0��|�5�#��N�q�����U^�{�9���R�{Xu�c�W���5],t�ƪ��i�*0L�ז�K��W�T�u4��˲�+�1���0���I�p'��]��6�R�4~�=,�RaSu�Py��u�[ 
���v�`��:p����m��p�˭i�/&e 1���w����_b'� V�Xz��#��½E?���-�S���Aq�]�X��Ice0�����2D	�N��
���/Bۙ�08{'�ЋHڸI��^+���V��qq73����*�s�a�U�-�,�� ���[l�?\�FXj �dj�/%L9�쐪�������S�0eD�Tޛ��:�Qv-h1Ν�l�_I�p�
��x.��l�%�2�0~~�jU yj8q��F��t�,��]j�	�N�w��LVd��-O|�C7����F��,�x1��yu��r���t����Ԅ��e�:�}����M+�ys�a���.ʅS0��NJ �i�t�+� I���wܥ�������q���X�ab"��!
v_)U�Y�2*��d����Ҹ���즘�˵�Rͻ0�A�q�M��i�Jg6���HN��O@H���nԟx��0*�n��v�q�[w�{��'���^��b�>v�]L5����ʙmI�$m�y9�|�0�(\�H}Os˖bsM���Zܵ�����I#ٲ�&"G�Y��npK�俕r����!{.�(�勚�SٿZ�V�c��6���Yc�~�g�ۅ��g �b�I��r��x�Ɗ�T���4R��9=t	����l���|����e�"�+��
9 R����j)Tf�A9�YH Tq�i����zf�^ ґG��d���d�V=�/v��S��Ηz�����5�P;@Ouf<;"t_�����X���x�����g�\����-��,X�FeW|�8��f���.��UՔb�j���+�*Ǿ�M0��F~Q�9I/����1�~]��p��~Ԇ~������9=u�xQ9�@���i���U��g���1f�A!bx�N����B�F��:�=��c'�&醈�e��EǇ[�s�i�c&�.(��{�G1^JD��cA�\x�zᡦ�!��j�33f�~��s�`	Weh	��˔�3��ZbC�ZT�g���l%0��n�2��e<8<
�AqZ���� �j���E� D�}�ކs���9�o4�N�8�P�Q��z�&�5y��I"$"�+r�ܵ�}MN@'ڧ�-�m��S�$5Y	*�Z�P��[E�q��S���>���хm嶃b�G�����N��MxS��e��k���D>�Q���*�R�1�oqR���aԎ����d����� v�sX�*�:��-4dB�ܡ��뇺z�ˬIB6V��<&c�t̠�V3��d%�5���-�dFB���U��?����P,��~�U\t�|v)��uh�Q�w��%4��^C{��!,����N�t��3�9|gHE�`���
4��Y�x�6T���Ls���0�*���c�\�[.��oͰQR��&z�s/99	�f�w��A�g���N���ЮR(�W����d�����+��ŗ��*Rx�����E�K���B=�y��ѹXB�+�B�Ab��k�6U��o��� ����_�@��LZ2�)��?��hw�n��X�"��M
�=J�ީo��JTù�Gt�'`(��ݻ��!��D[Eȉ=?��2���iښ����Poh�理�'ī�7uho��8�S�S�]^��/M#4���.A�c��zc�>0g+� j~{*\�ZC�B�Y)��+f�s<��Zj��!����;H�Q�Z��c�����K�!p�J�����km��ìKg��q�s����U�0�5dm��FS��oᒘ;Y����F#��u�2�	�����L�����%Ic�pG�d�Iڒ�m���V%/b��>��5�ɳ�B�Y�fG��B*M�v�p�^��꡾Ŧ��f�.}:m��Ss����[1�����~��$&�)Y�+��������Y�V���8�.�Մ_f����0�k� ��@z�m!�z�v��J{'`�K�[C�I^0���&�T3tQџ']<L͏�c��W�������z����m_�5�����n��ɻlK���5��v��&�(��eDp�9U�\��s��iq����W�$$����W���@
<>�3Q�Z�bו4��8����(�7#�	"s8�OS�
��p��\!�Rc��ȿ�����é=Gn�R)�z��ʋ�GN���;�R�$;�3�	��dC��G�4�j��<���,MƸ�S���&��0�-�s�=0,H\�]�e��!������� �P�����+B�X�p������T�o㝼�5>PG�R
�4�qLu��E��fKph��Ӛ��/���ɂ��`���d�(��B�o�OlHsE������
/�8�=:���gJ� ���a������@�o	�4�]($��y�%�7���`�
T\<�Ѵ�Ӎ#<%���v�x�6q5�����i�#��^�sW�U�qFe���,�����:���H}�插^:��D���k��8���2��5����۵A�J+oi8�rly��x��kv~�xu~9���H�el�\�w
!pdRl�[�{FH%��)yH�{|�����|GV��X0ְN�_�Mb���l�t��-�%[�����F1!M֔�n%�؁�\����k������%ڠ�7���O���O����?L"�S)�W��b� �"Ɛ>D
���¸
}�%on��}�s�����.IpY]-N�H�g���;�d�::��%���Ϩ`
���g]C��0�}o1�E �q�]�V�eպ+rh��&��Ν���/-;��a�"���NW
�gNg{)
Q䂧;hz!�B6%w���1�]���M@�)�]�ٕ��E\��7���^L�Z�����Imo�c���5��o�+{1��s	�o�h�b�,9iĿ�<Tr���- ���L����̕��/�O�߲`C,�rSͶ����KU䓽ً��vL��-R�b�Q�B��Kݰ�V���U�0�42���c�c��4��GΏ�_�S6L��/J��
r�j�V�_�M$V8(g��.y$�c�z�`5m�,b��?�eW�	D
�{*%b�����N�p2�u�ȱB�u�`�W#�è��HX"G Ӱ�2�q0�y��i0|�nѦ/��L�M��M���_,��@�`eQ���Z��ߔEe�:�8��b��lj������<�;F
�xQ"�0��QSUX6�Ć�O����M��ן�%�,����iwFo�i̷����U���A8|�V���u,�wkHڿ�܃��& �P��Չg�XvS�8���]���M�!nj�k$$�G���8]��~�qoĕ�p`[��\�F2?%�l[�ҋj��D�<�����vm}�$�d���rξ�Rhc5M�.>��!gHmS5��2rM�|�sw�j�6Ņ
&;�눠�Ȥ́QM\{�a��۴�7�4Ξ:�����I\l�Ѩb�]ǘ����N���ѳ�"��^��I�`T ��$?9����C��JB�ތ�+�!m������~H� ���A�$�ȴiU����\�r�d?DND@�mZ��1ke����4��'��Ü�씈n���M�h�J���O�1~Cp�?����B�
|����G2ve
)���9���,ݢh�r�&�Q�9���Ƨ���^t4�`�T]$�s��U�������_�P<Ş�m��:x��φ�,�55�._����1�hu�-���_7g�4z�6J|�zv��\6� �U�i
��F؉ٗ��P�#�vSDo%�n��A�l���^<g$�q�嬒�~߶�lP�*��Hְ�
��G+��bnlhc���aA0*�
]�:�����j�2��Aϸ�ZI���]i���Zg#Y�|�^v��s��0��G�E{�<�;=�wV�殦��E�V\����ʈP�}�b�Ȑ����E��1��8����.��ޭ�T�#UI�L��]^H���0"O��5_f�3�2��:(/t7�����7������x� �#>.���fzǣC�UY�r�3��r'�@����%t�B�le˛�M?�I��N�xz��sc�����z��״K4D|�=8�	a!���.��jk�p� t��=m�K�Ļ�����TO��S�y��K�bt��a^�H�V]q�U��YwflfT�Ɍ����w@���p�&o?y�{h�|=����,���_�:��(�{���okV~�際XqN�F�u�2��c F�nd�*V~۪E?��Dm@t�M �/�$S4A@V�A���O|���b���x�G��<!�e�t�T/�CG�'8�qI���w�%��b|/�qvS�,���s>QŸV�_E�3g
�'Ri&�M|.����I�d��M1�K� ,{�d�y9���{�i�.wAj���$W3K����._&���2���<�y+����O����m+<��?\'�䅝�Y��E>9���H;$���5e����$��$lE�*(`���dH�{$���њ����Ov�}_��Sx��� �`u�����X�+��R3���xp>�,��JR����Ԭ����8�(��B!���	�Q�'$k���8G�XY�}V��m��Sk�ñt!ب~3�J�������A���&�>,�,j	@4��tG�Z-ҫ��
�G\8c��f�3�QE����"R�L%ݰ�{�rXѢc�_1��n�O���#� ^>�N,^Xiڸ�N�Ͽg�����oY�+�S(��z*�ncx^���뾗��9�����1��������we�U�'�eDk����vs���w[��`"��8�O�r2B�jUZ��{��i&Ȋ���	6In�;�]t�֙]�r9�xD�b~�Ϥ�M���c��jH���x�z��j(Jĳw	���3 I�	uc����gv����*�м?��S��d\gF��)9���y�Pc���O8�-�Rrf�Z��;?w�nVاO!E����'3a�����8R]#`(���k�U-}��9��率�ɒD���	%��)�UC�cyv�o�+
Ǔ�qM���GL����O��^vy�(i?�d��j� g�ܭ���2���^��֓'G��=aʒ���%�VGS�YT�~Z�W�1�)n��3�&�Ʃ��6-�OF�*>%�xO�Ǡd���b{	��r�M��^!��U�dA�B�k�G��a�ԃH���@��:@�UH3gĩ��,���%�S����~�l�e�v��M(� �CA��AU�,}k�	m�a��}�`�V����r�����>BR}ݒz'M�f�-��0�k��V���$�/E_�g܈�4�e��b��+Te-��)<�FQ�[SLO��-��XJA�E�����髿�o㩢`::�WFR�(������:9鼋ή-đz]�A����/M�S��@���V0�ޙ��*����㚎ٗ(+�cκ*���.󅶦�)���=���R�u�-����31#�'�Z7x޿��TCO}7^ij`�B����%T	���t���0�g�Ai'���2�hhn���ЩRr�>:"���r@���Yqm���f����8tk�����+Zd�8���VAH��Ӣ��(W%h3)Q��T�7Ѷ�t��8zz��o�\ڤ��r� Y�>��0M�ٹ�B
G]h\а�cm{�P���	e�d��(��ى&����Wb�잉Y� cC�g��� ��2p[ �S�i�m�4�6��^�����3�a�G��?�f�LB�aJI�}O�2����))�[��35Y`Ԣ���{!`�j㊡�t
�:@`�
{�������	��Gs@� <�j`Ĥ��KA�׫�@��$�u��p�˹��u�2��t��{�
8���]��!��BN
X�C�}Y!�8����ў���R	\T$�N�c����^ �z�-D1̜p�d��2R-v�Ys�'�L�a��,eg�7�i.��\�e�Z���NL�t��U��&8�f8���eau.!��`�fO�������>��a�@�
g.�[Ⴒ���@[���6�ȋ�*��	�<����f���AK�����P��fZ��㰋p�����{=N �u�ꐚ]TN>��CG�o)���5DF�i��gw��%2�dGX���`�@����<
��݌��6�\s�F���}�a������h4�`jd���K]��+�Q�&U 1�W
<�H�Wk��@�uC�S]Rz��0�.��!�be����tm��8��#�00NL�_�d�?��h'@���E�����z�ּ/�g7`��Y>�AM*ݒ�y�ZS��;�]쌏�qGH<6A�����R�[`4�n�:9hj\�������^�X'L!���(k퉩���#�D���Y����"c��W��k������B���?���=y,���Wr���;w�d� h�[j��Q��b����Y��aZ���]�m"=��#P������^o��"�+u)�Pӯ���g!��>����K����5WqV����d��q$?|1�(.9&v���1Ä�f�KI[d��T�482�ǉ�䕌w��0K�q�y���M��fW����y�5ύR��0IxZ�n�5��{��]L��J��\
#y>'X�����I�8弖��*^�Q+�@�>�{m�ڻ��R�ev�ۇ��u����ќ~3�C뒼A��H�(7@�#&��!�m�9$;�d�K)ar]t�w����y��K,T�Q8�U(�/Նm,�^"�N&	ٱ�(}��$�-��SWG�8ˁ�_��Z��I	ׅ�� vt*Ŝ�V;�:0����i^ER��|G�+k��s���45�4׊w��@(sԄ%)���0f���<� �ظ᫁q�{�"@o��$s�IW�D�5M� �#'1�_����衎�M�r�s����hEFS�5[��緰p@OAs�ef�����:M�E���ע�%/�G���zi���Xd�$�)�4�q��N'�+��Ob"V��R��`*|�iA�2X�B��3.^?��_8���~'��г߈C\�<�@��A�U�K��O�Z�Y�`&��3����,䲋W.E�ZJl(�m��5$m�`"���}�Y^k�'��k�CXBɆ��J��Դ����^A���.\��֘H+#/����ҥ��;r��M\a��s6�Ȧ�[��MZl�d�Yת=rx0�"�U��#xk�`U&`��q��;��Ji��%���������@��7Dv�e�ݺ/�(�"b�R�z�^�Ǫ�ɟ(�>4��P>Mm|��,��+(���W�'�z�����J��  ɰ��_y��X�H�o�UO5������8j>�:�&߆}�X�$�T	'���x1u?�s�)a���;i�A��\2⨒�	+�����=0����}��L���r��D�w&`��w������Q=�����=����ש�5� "t�J��^�Ahg����M�a\\�pX[0:�0c�C�T9�q���NJ�Ӟ�zh,��dQ�1R���m��~C��ddY���U݅�փ��y��J�R��V���ee���$���<�0���A�SV��ka����O���h�j?R�1�%A)	s��Yl���ڌQ�Ok��ϟ�ۂ i���������׉ ">'��\tm9�<<ۄ_G�9�-X"Խ�@��h���	NR���W�;-I$�!隚ꗼ%Q��g^�T��tLB�']g�h}[��G��Ɋh���#o�3�C��|6����_�^�����u=Zfn��s�~/s�c+Gx����n`t��T��B]�5��ӗ���=R(l���8V���S;9���/OÐR+�!�)wM�$qp���a��0%� ��	�,N�E(r�P�nwе�>p+�bz�?�x�X�R��g�j�f�M�LX�< M�-1�t�lL��9 	b.��-Ǥ����~FH�J�te�U\v�܅hO Ɂvb�� gɗ���'\���Wg��`i�~��Ӏ@T��]�G^2�<�Dq:�r�:W�c�9�|��B�~���椀���fp��5:���k|]ד$�Ə��s��Ye5�|�/��� ��PX�x�����r��5v�f�{S�1��>�]�kB���^n���~�,�)4��7���ɦ~ZB�Yz(�2{�$�j��`:��K��������!�����`UA؉����W�yR���U�,&��m�<#�vY�s� �[��z`���WT�Ap�w_��	��}�	�k�Ku����O>�{PT�8�;ц��t��Ƌx��g,�{����S����7xOF�����8�[� ���}<N�C�f�����&vfȴ�"�Y���}*k�x1e\��A{��/ߛ�Cl|�k�ō_膈(���Q���a=�i���(x۶�_�^7��2�h������:�����	V��-��?��2r���Q-��h���Mx���/�g̀wD/�H~�r�Ě�L���x5���.l�<>EB���Y.�4L�nO�=CI���So7�}�)v����1��uA-��(I���R�Hݒ_��	��~�����*�6��K?���cs7؅�F|����L�&����AR�R���h���bA0>~U��$���>��W��N�\��lsg��'tmG�O��I7��#;��1u5��m��Di��Fƿ��;��{�J\{̧1�iĻ �3rX)��Ъ0?t�lw+�sJ��$*�z<��	�%�hi���>thv� E	�j�Lb�'E�� �ZےU	����Ax��]:��}v���薚�<���o���̥�Lp�V��m�ܘ��(�(2��͚�W�I7�Fz�(������iNo�o�:�Ab�·?n/PY,�K����/�]q]Q9��]��Nױ���W���8�^��d6����KBz�$�)C�-ȝ6�tsްJ��j�ƹ �*���6��0����3#�� ��*�khپz>7�v��[-��ܹ|[�F�x?��`��$wUs,Y5�j_����(s��Ӧ!�,��ɿ����f���*��8����^���c&�������:��0��zlV��n���p��sĺ�`'�j��A&Ն�1�5$�âD��uU�{�J���5�=m�ٙ�Ub{����!��{�!��л���f�q��	�FV�6D�)�0�4V$IR�E�07-\m���m�6�ē��.e��:�,˘�gd���я䌸��H��g})CZJL���0i���Il�_�"���%��3�(e�l5��5��(7?�ā��g����>�̟	�Ō��5dK��{	�8�p�:�w���E�Q�瞲.eX�I�E���Fco�E���*R��N\��5��&��Q�N!Q���"�Ӻ�q4��N:�bs�3�8s?�Nb�,z�1��ҍ狓U�� >���_2x���I����� ٖ�㡷�g���&�=B�M5=3&B]Hl-�-�J��`��;�ՊyJZU�y�f�F���pG�=����/�����rUˈLճ�g���������F���&J��5��[�n���{�}��:��+����bP�!�(l�r3Ɇ�X;��t�i�<�qއ�fʰʶs��u���-U�1��,�����ݪ� �b� 6t~
��&Ky��7e�h?���Y�j����&���ݳ�� $������ʔ�7��8������4�uY-`��Ar�{���wS㑴�~e�{���|��AG�N�L[�a~@^��FY����Y>��O�]��a@�������ݮ��'��#?3��a!���F��3����ѳ>�*iue��Tؔ%�_~���N���+ԫ�1L���	A��n�EK���0�.D.	����	ܘ`@qA�CCܩ�DM�s_����=F���N�EF�Fl¸bɝ�p�-F
 T�p���Q|�����(,�nP����j����¬�^\q�(���o@�@KՐ���1ya�;4`��.���Ֆ��a�ҕ��[a���� V����d���I,;�@�9?�ԯP�0�
9��8��k� ��� m]���d;�C}�,!�õwk�t�M�Z�T��t���j��z��R8��W[G�hv˪��%����6CoD��%kB��g�e�V�a)�1����lꌣ�b�"��5e3EPWۊ�%�÷�j,,���Y�r��M�t�U���F1�iƩH��i������>��!
/Ϋ�9��Y��PK��f�ɔ6�����	b?|�����ƨv�.�򔻔k����lK��ރy:�.`
�ӕ���?De���VGܤ�|��U�Hb�y���	Y�w+p�;tV�o��lYSܿ��@{	���,n	�>��Y��I�_����k����/=���CJ���Y.� �l�G�!ȯ {�oo��@-�,�FA9�	�I�4����q]&s��-,��.o灰^SjU�[�E'��aq��&Ds
I���Y�j���Pd[�P�ʵg:�;iJR��e��@+;������̗5S,4M£�QT�S|:L�Y	�9>�L�1���9W�ό4A�g��o��r�"�mD�SZVZ{(?�(Y9���fR$�:M� ��OFڲ�d�CQ�F������ݽ.٘����ƨ�oK~H&ˊ���� $:xR�S^7W�}*�t���3�7x`CS��.2O	 %&�e��F;��d�s���(��{�1,�]�{(�;��W�{ө�t�5��d푯����9jo@.������}���l�P*l啰����c��0x|t��o)�j�c��5�MA�GA ��q8��m�S��4��n��G��v��o��̋�`�+#����|tޅ��Q��}YB��H��6��5���ܘ�X'G�1�~V[�@��AX.�m�+�M"H@��D�T"[��{���{j�@��׾�R-PJ�9�ƺ�<�xu�� ��[�")Q!�Ȼ=]ζ|�`�'Pl^em�a�|$��V�r�
�k0[��7�9��E�&�V���^�<(�l�����6���RGS�P���+�q�w���r�w��X:.RT����b��@��#
���n�8hKY�e�Y�G�X�w�K;
XYz*���;~(���`|

����:n^Ef�Lr�#�E�S�'깸��3�6�疁/O-����$����n�`�l�T˸��L�~O�Wf$Z�nHe�]�k8�%�`�����U &vi�=�J�u����	p,,8rG�/[��͌m���������vZC� ��N��X(���/L�_m���c�n=��|C4	�c��o�;�g���J�|��[s���ϘWtʞL���[E�~%k\�}�KQ�2�!p4�n�K6�v5��������%g��9�φ�J��HWTZY�GM�����L.&e�;q�o��I=�'�25�5�gd,����R�	���!�5IS7��Bm���Za��IRu��ŉp��V�׹�U��~�� jPq2�������01����!t�'�2};#�Q�#��7)�l	�� 4]SL�@��] O��$S<�IO�7O ?� ��d�{����Y%Tw���#���hU@m}�@��qw�o[�r�g�L�dgHu,��trd$�P��9-��Ͼ�n�L���wX.���K�(���?�g�h��8��C������KCkM�@fHV2�q��R���nԿ�5��,7�J9s,z �@�%jE ��>��9=Ũ�"NFf|B�~$5gWR<ϸ�8�t�ӻbhL���rQH�5�p���fTkd �Zc�O:���hE�aS/�6��J:�����0`�6�
��-��]��7���G�}]Ì��������ǒw��KL������>«���Y����-���J�{H�]
;�V
����aCŏ�QSQ3"�H�}'沐z�{v��ڣnG����q)ެ�}�=��E������Xf�Q����IJ��� �%y�hjqZ�R¿���"�F	c�x��q��p���	��o��$+�ޗ��D��Ӵ��#�5�@r�Q����G�q�y�Tw���;`ؽ��5Q��v�k�	�i��\Pdy�w-0~.e/�P�)���Z��&��K�4��f1b������]�c�˘�,�d\��G�<�=�K���"���ɘ��,�K�w�M�E߱(O��V����܈n �0�19���g1����A���K��e9ŝН����)9�`�``^���y������i�\� �2��$���@Q�d="+OHA��q'7�{i4��1H�M����l���+L(�����f)�w֔\~O���z�B��ǻ��E.�|��� �7�΀U4�$(����L�q�(���8�q�L�I�FЪ��X��(-7����T8[�b͕�$ Q�6�8��|�H��7��cB���Ǻ����t�=v=��d2�CF;� §��%Q��Kݑ�) �R�Y��N �:4�|����B�i�5��?�.0cs��Z�rh@//�	���b��U4���f�$`�h���v���S��z��D����Ik�g�=#Z$���l#&�\alHu/˓j�B9b�Y�/��^Q�/EN�"���{}� ����'�������1"2���2h��HI�C�X$�(��Mi��b��R ��	u9��3��i�\3o�v�ᵜ�,��˟�n���Ywǿ ��e�nOZ����.��x_�U0�W��^���'��(�QY�*#hVnD�bK��}hO��L��i���F�P��F��c�k҈��EN29���//�S@6��;m|y���G	I�	uoƊ_�{(j���'�W4��,�OX��/^z�I����+p)�k��5*�(�u��5���_���U[��z�t�pu��bIH�
r��$=����F�X���x3(8�46��a�y�G^�{�߈ُ�,w24<B��Ӝ�<��'+�_+Veqo8nd-�%�sv��j��F'j�=�5��]�s��r��}i#�ů	G3�<�a�2�V�V��o�ُ��/�o��A��+k�&��3����lv�\~'������E%���DZ��(M� n���.����1��1���E�=c��R�+��[�E�_����Dr;��hr�ך1��Cf�f�һ�����G����Y��=�z�|��tS �ё�	��[dF���/,�ԾP=V��l�"A���j��rؒ"2�C�X��π��K�m֡�P�C�Sa�� �b���T��%�M��/L4�p�րIYP�������}%@�/9)�/��=%/��Yc'���6�J�r�oE}��$�س�KoII5�^��������N	"�OL�ٲ~m������CO+��H���{��ߊTy��ޞ�[�YFR�p9[��-�S���v=m������J5�!㇁ţ)Cb a����X�Z��ǘ;
��N�auv�w��O����Y�Y0����|���������o/mb���}�oj'!h>��:
a�G�)���ڌ�Է�*��N���y����@ai.�ww�	�I]��D��Jx*:�I~D�@�ߖ�s(�Ӎ �q���Y8=aV���<Nk�����p�K�`�>�É?t 9�XߦC{��@<�ba�����hnח�Uۘ!s29��&��ѷb@1�a�Y�_���Ƭ��P����닫�?=��⻴*���z�[��P�j�m��G�|T���]�i�90���{�u�B��3K�ۻ����n����&���lР��c�G������GP3L&Ú�=\��kΓ��ǜP������,nRc�ե�L^���+/��^U���*?��U�J|���)�PZ��u�d�if�d��B�F,���o�L9趢j|	)19��r�e�F~آt7�p4��-�1�}��]C�&��V���љ�x��,�r[����	V�~y;��K�������L��]A�T$��l9,/��T!d.��vv٢S}21�SQ�J�'H=���9W1�Ax�>!�P��5�%7Ցq���*���;5P�|���N�T>�w�7;�{s�[Ϧ�t�hq5�Cf8|_3���g�P�x�����z�}K���Pw%Z_��X�#���!F(W��Z���XxHQ�0�J,:��ۅF��(�?,�_$>�d��G�i���D[!cww�R�b>�e�).YW�U��%�~��zI�YVy�V�ETP[���v���E.���\��th�u;�����a��EI���5nҳ5T�=sU���-E��Q$u�Wh:vt�v��>��8Q�Hc��Q|��$)v�a��p������t66�`��^����j�z��Y�!�?�f>��<�����u�l���`Çk=��>˒-��M���p��x��\�����l���1ճ�`oj��\���TW� �)�l�µ�����
�+��ŷ�al�0��|J����[Ƿ�Z{�?z0B�zE�s����5��Ys�����"$�H�G��O��ϘGb8�jv��ŉ� n���^e�\���W$�Nim�1�C����� �b��Q��v��������}`�J��+��o�-3���m���`҄f!^�A�`{�Prk%�/��� 51zH��l�kmr�U��/4�Ե�A���>����%(s��˹�[b>�:�u4�����9g!�8m0fZ&�kI1 BD�/�g�}�4�-൬~%��*<%�6�U3�&�M	�3/��7u�[��~�P�	%��r��,(s�N�� �O7��R��������݋X��L_�/^Fx�G�k���ۂ!É��G�c�Dm$\����+��kB���� 
���[�"\�'��lW���Y���3��XƲ�V���禞�l�"-��v��Ʋ��>o�h�Y����a��~�pd���E$����4�c���^���VQA&ى
lɍ�V=%�c��~���M���~:�ܽmc��C�tc�6ʢYi(b��>�C{a�?�fނЃFKG�n�-^����B��=Ӱ�Y����"�:��Xt�!�_�aT��q�y�����5��<QB�����$�:YRw!#�s �[��<�u�iԧ�8��f�G_�G�d��蜲�ĉ�kh�!�`}B��C�w����Q�[�Ѯ��6��=�|�
L3qu�i�WI~��ݶ��9���,���>8�Xa�3asn�&à��1.�Ŭ�������Q���LM��a�1���-�ŭ}ޭ���z�7.,;<pnk��q97ԧ�K}��{�懩}ZF��t����jQ�i��6T!]XG��et�6��4�7I��1낍�^V�M�c��	��>�`�#��+9��D{ғ����bNG⣼[�9t0�?e�ϖ���A����������,�3�T~IG�Y(���W��H����8/��8ˠ߆Q�4�n��A7[�W4�s�O�(G6�T�����\s��ڡ��ư.��ӌrN ����=��[�w�L �"�EB[�&ZI�!���|�7���GH>;f�f�〲?�8ݭ[4B�7���`�bt-����_p��767"g��AzM�� ���{ݩ��o|�Z���e��u"�Y�2�� ���K@	i'LυY�~���-?��Ň}i��=�K6�a�xf�Ff;Ц�au�yO���!1F��f.���/����o�P����"8�"{�s���@c<+���?������ �Y��UA��=�/4k�����@H8�����-$��E��_�!��C���Y��5 ��e�ߴ�%��U�*n�G���;(�"�N��n"6��p�.[�H�+<%[���0i8*����n��C��i�k�*�����&��LQ.Uy�P�Z�U�bCh��8�����p�ᒢ�c(+��-�Q�Lh�	�����y�(��i��D�݀���$�]D�È��E���]RO���O�3�M���S����U`��w���[���;��Lr����1l��E��2���`�t�)dC?�=�:wI��]�fM�Yx��Mb�V�s������a�ZP�s`��`(U��.k*��.!d���U:�{�0s���$�s?UV�7cxXM6;I�1"��_�ڻ/%E�H��TV@�����������b�|���Uh�/�Y�K^�j����i�h��o���z��Ian<�}s��������9t�pB����H2�@�'��wk�D�P�ѯh����E��D�{�K��K[�rpw�q��H�l�Q�e��|�Q��g-���(�����ŭU�^G;d� Mڏ�.X��.�sD�_R���n�g��klᴚ�cӗ��J�1��$�.��U��	G�+�rz>Gn)�TӥN_�$�~�m9�[�F��8^���şq�Mc�l��ޛ�k����tM��_E�
�_b� �vo�8��*�kvԬ��V>���Kt�'��i,��p�4v����2a�+�U!6�c.��D�r��C�Jײ�ㄗ��MƯ�l�?�(y�69�9|�P��p��
+��3������Tzҫ.F+��w��A�ɢ𭔒R�O��#��o'��HF���kq��3�=��l`��ɱ7���$���Ȳ�J"�s�$���d�iEL���\����/���5ϳF�����O�'�$H�r������P�fI�
�j���҄/Ȼ�A%g�߷�7LS<h��U��cv����������g�K�<���'�Z��1W.W�'9�7��4G�m�9ҿm��e��1���Q��󞶹���3�T,�T�W�w�������2��,�(c��F���}TG]s��V������+S#�%�5� F���obL �rɁ�� ��m0���tP�B��z�V`O��������N�8�j�-����b%=)���@�c�V�b�_�X���m�4[gP�wp2����[ͧĖkB����_�gp�������X���_1���
�}�O��nok���6	Q��<P3
�����B��5̫Ŗ������&���R�ۅ^�;1�\B9龔��c� ��oe{���l�*G�ĕT��>
�Rݓ���Txa�8�"5B�~,N�?#�J"���v��9�VH�?�R�A��&���+�$��qb�H$�7��e��&�EF�d�Ȗ�`��/��j̤@�L��!5�,��39�����0΂'��{����q��'�U��ܥs�7�6�E�>�����RL9'��N;)����f�?����߹��e;رZ�3��`�b��Hd\���m+x�}�N�(���;��F�ͧ}���u^�z�x���f���آi���z��VAϨ'z�#&��#��2�b�ڕ<:�9ְ��i�3���� 1'�����z��z����=�%0��z�~=�)I5<�iH��^u� ���.�D2}Y����	T�^�U`�x�����C����P'U�a��c}e��	{�u��8���E����R�^$:���Cj�c�p�}���V%�#��}8д�{>��y�70|"�ݸC9�y}-�$7q�l?{�|��d��e��(B��A`ks���6bS�����IxO���>�2?Bn�oH*��������ˋ����n�{S��)��!�<^ٻ�����]���Je�iT�߫��}6|���n��8�F�:��d��j)�@\���r��hf�,4Q�o�b�?��9�c���
ׇ708��Z�G܋�)/\�7�{��}�L����s��b�&MڇBҠ� &�
��|[�Ɠ�P�!�7�m��cl����
X���W�$3iB��p֡�ET����hނh�H񒉣|x����0��������W]��k{���	嘎�s����P[�rBOR�_��vvcTR<lSx"4�F[9�70��~{o���a��˓�&&���S���s�T�8꠆�m�n�6�)��_������������w�#�Rv���J͚H�3�˷{.�}�:��&id�!��ࠍ@��HN�Q˪C{�#V�$���ʪ?T����L��:a�ʕ-�Bi�Lt��d���K�t��4`������=��}qW&Y��A�``(QO�g��1�2x���Y�*�f�>������;��x"���1�Z���Tf(��&�W��C뉉�u�}z{����_��HQ�k,$�
e�\K�����q��ڇH�2+�s(�Eb�Q* ��>�<$8�����'�=n���B=�o�ۜB����,!N���Dk�p�T]�h���s�^f��{x뜺�8 .��A���R�41�axX���y{,v�k^f�A�4T�ΖS�����Sy���d��,��N�[͑��|�}ٹ/���nIc��p	�?�i�"��5r�r��:�|̺��f��Y�lNvL�ٛ	K� �[�>�>���� +S੪�xk�|C�Ơt>2^��u��t���d��F2z惈��(l�ٹ��Q����")���wY�j����sE�����ΰ�1���7�o�V뙇��N�6e>��pNѓ=�E06ҟfQJ�	�;�mz{qa;��̹b���T�[_�kw,L��� @���ww.��h����Ӛ�g���-�y����f�C�3 �0 �Z�n8e�߀3��d؎�y�ѵ'�&Q�&��>)HAjD���j2��~Qg!������qt�e�A@���0��m�V.6�t�h��b:��}D�����4=��s�<���!���3��AL�ҤF���=�֪�B���| �����2�wیw�,~}w\�ɏ�Z0���SثGہQ���7�4��-xG�4�-���52�ȫy�Ԟ���'�<fI�G����4�]�B���C}��b� ��BW9@���j�^�eut��T5��W�"$��BWB�0���y�T�}�o�	��k�K�M�M��y���n6�����=��̓��	�kCph%ZE~�S}t.��8[���O���ż�i<�P,�WD&� 48(�N��������ḆG �vP�߈�d-���G	��椓��S�Z�~���^k��5׍[�M��*�Q�,��϶Y����R�r���=2��\���ȑ9s��|����y��dJ!��iD�&M�j�
�i�Q���d-�
�IM��L��gIBF=[<�S�װNL$�*i�4ix;u'iO-�~X-%c__ oV�tl�m�1��X^; ]��6C薰�v��z���>��9w�q&��o�1$(rb�'͋Q�u��o��Si�ݷ��x�>�!f��?���h8����	 Gv~�p��wm($��w؞N���o_��S��W�Q��1�)�W�G�+,}�8�T*|�*F�DV	8�d�?fj&��j�����NS� ����:G��YNƣ��B񼒗,�-��87L|y���s"�2�O��J9?n���{D�P�dC>D�FG�7S�޴#���ͳ�H�a���}1�F�ӵ�J�5��B;�K�^��+�����.�	Q��c ��U�8kS�j���f<��K�`���*��=�J�[4���CM�Ҿ�mBs �/��)�Q��Ƈ���?7��b��g����T�L�"�P�����J=i� >��#�6��W?�mK��=�'#� ��h� �֎N�	��bP�?��Z"�ӭ�RǪ0Q���`JuL�_�K3 �$�D#2a�&NU�F���K$?�5���B5�*^O<Aʚ��|rx\o�#���^v��+8S�+Lq�'U�+yQ0��	k�c���T5.ʍI�o�"��[x޻N� �M�(�%�H!�� �Zv*{넺�K^��t�^�`Խ�@����<+v��T���h���&��+�3n�()P�+����^u�U���.�m51���b����
`KѥXK:\KMs���L�*� �j،K�@<�E�E�J!c�f�	g�{|��n}��/l�W0I����y����������%�=��[E_�zT�(�4�NL|q#�G���@���6�p��@��C�ݐdBZ��S>�|�I
+r�HGIF<�v���TPF�lr�F<��PWs�[V}��A��<*�1M+�w��rO-%#J���۔H���}E�ߨ*H��M6��)��6� ��"s�	M�\��4p����'�0��	; (L��}���*�jA���`B:�:1`�<
�ay��|M"P���U��~W�<��2[M:��׌6�8P{p^��9Ȧ|Ð6���RH,,�zt����fD���cV%��>s�X�8��[4J:w�O%�<<�hQ���˃R�{Fc�,Լ��[!��e�W�..H�N�{T,�6ђHj��n�_��a¨�������"�����ꁊ#h�+��ѣ,B��Ju3�=�c3�̦&�ɭ�	�d�pz)p�O���������ݐh�O�܇?̎�s��Eo�9$&���Y��5��B���n/�?u{�^�@I ��j�ǆoh��'$���%\���;�{vS�����1)4,���wC�YW�<."qz����o��bӞk4N�B0�^� W�@gt�y	�m7X(/�[�Yz.�,���]x��V�������H��r+ ���X/3�)�T��
M�������P��K�5�fcW���<K�y��ǭ��O��?���o�h��k�
�­���L䀜McfX��_������Sw�5lY������O3���� �hջ�_�$_u�>�V�G�Ѳ��N!�">��c5jҢb��k�e�Fe�«k�zӽL[	_/���i�<�0̐���\ut	��Vt�8���L�x��@�S�L+�{㻉��$�O�o����F���3�m�����oQ+��:��Mӯ`&�Nj�bhb���6ޝ�v$Z.��H���'�j������n��w��e�h{uB-"V�h�!ڥA�vU�^N����bx��F�~������׭�,���\}x�Q�����wi5�%��H��nQ��$�:N렙ڰ��'��IU��R�̞�3���X��C�������Q��F���j�R$Lhr4/�O�j!��~�����7�h�K+`�AsY�5�"��s{-/�}A��w(M�kb�T�E�jan����Yȟ�s�h2���GXb@���G�q�sU��x�.r\�U'Rc,�]����\0D���Ws	�?����{#���Ұ��*o'[�(p*_��g1Vy�0��eY�Jv^R.'W*l�c�'����ؼ�L�F���P����Sb��cV��d����.4m�e%�-�*>
�0ћa��f����@�IG��)��M��Y������lA�(T*��"(�c'��E_@���{S�k��I��Kz�ݠv S�6k����h��NO���O��3�l���E�\�� ���D�G���q̝���F����8�_SP��Ri�'�k�F_�[[`��w�=9SRޣc�W��:�W�h\���+8��M���4��.t�<9nJ�����g]�7�)�i$/�l��S�t�4��ȩF0fL��zLs��%d~V�O�%�)��(m�����:��S��"��[7H�q,�`��v��k�j�!�͸���ֿ�<�h��%cȔ���R 	��*7H�?�,�L�D���"�}�e~h��Q:aG��h�_諺, ����DR@+}����8xo~�3�ku�4�m-;L��$�q��b'K���h!�:I;�����?
?]���w�\��eζoݳ'Sk�6!�3	��'����)j��L�t1�OF�j6���$
 m1B� ���2���1n#�#ǔ��|���d��Z�h��}FC:YBܟ���+�ă:ZtY�W�°��x��r��4��/E(�2G�mj����v~�FF��d�sX�u�_O>����讂�cHrС��8l��8�[2�������Ěj04�q�u��ґ}��NC9���cn׬c>\+4��VA��N�����#q9��q �}%�aY3��F�cY*i�d�:q������^Rb�-��crth���*y�l�w��5�9Ӿ�t7ʪ�)g�5��f��1S�{#=Wى���C����О��� L:���@�8�j^eA>�w�{�ǐ$wө���-e�F�<|.�0C��-��4���q2�r;Q�:~<�E�"i�$�x:���p����b����s�4�A�?��;�g)zB��a��zBc��(!\�FB��<xԃ���#�M;����;��Q��u�>���;([�n����^p~�ۜY5�&��$��8�����2D#�V����`�N$�or%��'�-�	�.���!2S�Py��d�ɔ��-KL��e!��G������1Ŭ\|#�����(-e N�x�ѹ%0�aO��ú{o}��a�+�`��-�&���LG�v"�gdry����2����+� �� �3[m�ks�E��ѭ��J������r�0�p��lM�B�[�,8��yB�N�pZ��T������`�A����Up���~�@�g�l�	8��F�Kڞ�Y�@���j�����v�C��yo���M�C�#S���"ܟ�.��K��"�}��U k��=� S���B� &�6#d���+Vrg֐��j�/SΡ�L���(Q*w�.A�\�胐g��l�xMfES�8̍A�e�������Y�lϕ�X-��G{�s{���za�T_��"�Fc�}	>�G\�.Y7�2҈BZ�WQ�[>�rJ�*�Z�}E���yѯ{`�:��0��P�F�����FV�5�<��u��9U�����I�x��E�?�jM�ڨqhc�đ��OD%��%,���3)-�<k�-��2�
J�@Ļ6�����ߞ���.�I��x�F0�f�ά�G8Yۅ�k�A����Fi�R�ԧ���	]�i%L~��N�B���c��t�ۇ�u�Β�p&�|݁cdh2���1�!��ڊ���ҙg���h=�g�1�����|���%]��� M	�͗�1mx�i���)�y�,X2���|H��V�`�t}0�%��y�/8�:b�� �[F�Z]�9��f��M9>��X|N?P;̪=�T�ی�Q�И��-��;1��ϐ#��Y�[@���"�Kd����w��� ,��"�Ň����t��.�/���\dg�g�8삘�=�Ǳ�
 '���m�h�`�z�<�����$xx����"����<Ÿ�ݮ�O|��F�#m��XlL�\�]mH>����h`��H1Qq�fx߸xh�!+�%q�xhù�e���7U��^��D�v.����W��e�ҙ �B!�1,(-�jʍ&*�w�,���+�����j�l���N�B&[5��	~�a����I,�X3^Z�����z`tu���po�5�ׇ�+�t���H����[����