// DE1_SoC_QSYS.v

// Generated using ACDS version 13.1 178 at 2014.05.16.15:21:44

`timescale 1 ps / 1 ps
module DE1_SoC_QSYS (
		output wire        out_port_from_the_i2c_scl,                 //    i2c_scl_external_connection.export
		inout  wire        bidir_port_to_and_from_the_i2c_sda,        //    i2c_sda_external_connection.export
		output wire        out_port_from_the_td_reset_n,              // td_reset_n_external_connection.export
		input  wire        clk_50,                                    //                  clk_50_clk_in.clk
		input  wire [1:0]  in_port_to_the_td_status,                  //  td_status_external_connection.export
		input  wire        reset_n,                                   //            clk_50_clk_in_reset.reset_n
		input  wire        vid_clk_to_the_alt_vip_cti_0,              //    alt_vip_cti_0_clocked_video.vid_clk
		input  wire [7:0]  vid_data_to_the_alt_vip_cti_0,             //                               .vid_data
		output wire        overflow_from_the_alt_vip_cti_0,           //                               .overflow
		input  wire        vid_datavalid_to_the_alt_vip_cti_0,        //                               .vid_datavalid
		input  wire        vid_locked_to_the_alt_vip_cti_0,           //                               .vid_locked
		output wire [12:0] zs_addr_from_the_sdram,                    //                     sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                      //                               .ba
		output wire        zs_cas_n_from_the_sdram,                   //                               .cas_n
		output wire        zs_cke_from_the_sdram,                     //                               .cke
		output wire        zs_cs_n_from_the_sdram,                    //                               .cs_n
		inout  wire [15:0] zs_dq_to_and_from_the_sdram,               //                               .dq
		output wire [1:0]  zs_dqm_from_the_sdram,                     //                               .dqm
		output wire        zs_ras_n_from_the_sdram,                   //                               .ras_n
		output wire        zs_we_n_from_the_sdram,                    //                               .we_n
		output wire        pll_0_locked_export,                       //                   pll_0_locked.export
		output wire        clk_sdram_clk,                             //                      clk_sdram.clk
		output wire        clk_vga_clk,                               //                        clk_vga.clk
		output wire [47:0] seg7_conduit_end_export,                   //               seg7_conduit_end.export
		output wire [9:0]  ledr_external_connection_export,           //       ledr_external_connection.export
		input  wire [3:0]  key_external_connection_export,            //        key_external_connection.export
		input  wire [9:0]  sw_external_connection_export,             //         sw_external_connection.export
		input  wire        spi_0_external_MISO,                       //                 spi_0_external.MISO
		output wire        spi_0_external_MOSI,                       //                               .MOSI
		output wire        spi_0_external_SCLK,                       //                               .SCLK
		output wire        spi_0_external_SS_n,                       //                               .SS_n
		output wire        audio_conduit_end_XCK,                     //              audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                  //                               .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                  //                               .ADCLRC
		output wire        audio_conduit_end_DACDAT,                  //                               .DACDAT
		input  wire        audio_conduit_end_DACLRC,                  //                               .DACLRC
		input  wire        audio_conduit_end_BCLK,                    //                               .BCLK
		input  wire        uart_external_connection_rxd,              //       uart_external_connection.rxd
		output wire        uart_external_connection_txd,              //                               .txd
		output wire        pll_audio_locked_export,                   //               pll_audio_locked.export
		output wire [14:0] memory_mem_a,                              //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                               .mem_ba
		output wire        memory_mem_ck,                             //                               .mem_ck
		output wire        memory_mem_ck_n,                           //                               .mem_ck_n
		output wire        memory_mem_cke,                            //                               .mem_cke
		output wire        memory_mem_cs_n,                           //                               .mem_cs_n
		output wire        memory_mem_ras_n,                          //                               .mem_ras_n
		output wire        memory_mem_cas_n,                          //                               .mem_cas_n
		output wire        memory_mem_we_n,                           //                               .mem_we_n
		output wire        memory_mem_reset_n,                        //                               .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                               .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                               .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                               .mem_dqs_n
		output wire        memory_mem_odt,                            //                               .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                               .mem_dm
		input  wire        memory_oct_rzqin,                          //                               .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,           //                         hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,             //                               .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,             //                               .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,             //                               .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,             //                               .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,             //                               .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,             //                               .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,              //                               .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,           //                               .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,           //                               .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,           //                               .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,             //                               .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,             //                               .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,             //                               .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,               //                               .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,               //                               .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,               //                               .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,               //                               .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,               //                               .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,               //                               .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,               //                               .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                //                               .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                //                               .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,               //                               .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                //                               .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                //                               .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                //                               .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                //                               .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                //                               .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                //                               .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                //                               .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                //                               .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                //                               .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                //                               .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,               //                               .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,               //                               .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,               //                               .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,               //                               .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,              //                               .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,             //                               .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,             //                               .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,              //                               .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,               //                               .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,               //                               .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,               //                               .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,               //                               .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,               //                               .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,               //                               .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,            //                               .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,            //                               .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,            //                               .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,            //                               .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,            //                               .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,            //                               .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,            //                               .hps_io_gpio_inst_GPIO61
		output wire        hps_0_h2f_reset_reset_n,                   //                hps_0_h2f_reset.reset_n
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //    alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                               .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                               .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                               .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                               .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                               .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                               .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                               .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                               .vid_v
		input  wire        ir_rx_conduit_end_export                   //              ir_rx_conduit_end.export
	);

	wire          alt_vip_cti_0_dout_endofpacket;                                // alt_vip_cti_0:is_eop -> alt_vip_cpr_0:din0_endofpacket
	wire          alt_vip_cti_0_dout_valid;                                      // alt_vip_cti_0:is_valid -> alt_vip_cpr_0:din0_valid
	wire          alt_vip_cti_0_dout_startofpacket;                              // alt_vip_cti_0:is_sop -> alt_vip_cpr_0:din0_startofpacket
	wire    [7:0] alt_vip_cti_0_dout_data;                                       // alt_vip_cti_0:is_data -> alt_vip_cpr_0:din0_data
	wire          alt_vip_cti_0_dout_ready;                                      // alt_vip_cpr_0:din0_ready -> alt_vip_cti_0:is_ready
	wire          alt_vip_cpr_0_dout0_endofpacket;                               // alt_vip_cpr_0:dout0_endofpacket -> alt_vip_dil_0:din_endofpacket
	wire          alt_vip_cpr_0_dout0_valid;                                     // alt_vip_cpr_0:dout0_valid -> alt_vip_dil_0:din_valid
	wire          alt_vip_cpr_0_dout0_startofpacket;                             // alt_vip_cpr_0:dout0_startofpacket -> alt_vip_dil_0:din_startofpacket
	wire   [15:0] alt_vip_cpr_0_dout0_data;                                      // alt_vip_cpr_0:dout0_data -> alt_vip_dil_0:din_data
	wire          alt_vip_cpr_0_dout0_ready;                                     // alt_vip_dil_0:din_ready -> alt_vip_cpr_0:dout0_ready
	wire          alt_vip_clip_0_dout_endofpacket;                               // alt_vip_clip_0:dout_endofpacket -> alt_vip_cl_scl_0:din_endofpacket
	wire          alt_vip_clip_0_dout_valid;                                     // alt_vip_clip_0:dout_valid -> alt_vip_cl_scl_0:din_valid
	wire          alt_vip_clip_0_dout_startofpacket;                             // alt_vip_clip_0:dout_startofpacket -> alt_vip_cl_scl_0:din_startofpacket
	wire   [23:0] alt_vip_clip_0_dout_data;                                      // alt_vip_clip_0:dout_data -> alt_vip_cl_scl_0:din_data
	wire          alt_vip_clip_0_dout_ready;                                     // alt_vip_cl_scl_0:din_ready -> alt_vip_clip_0:dout_ready
	wire          alt_vip_crs_0_dout_endofpacket;                                // alt_vip_crs_0:dout_endofpacket -> alt_vip_csc_0:din_endofpacket
	wire          alt_vip_crs_0_dout_valid;                                      // alt_vip_crs_0:dout_valid -> alt_vip_csc_0:din_valid
	wire          alt_vip_crs_0_dout_startofpacket;                              // alt_vip_crs_0:dout_startofpacket -> alt_vip_csc_0:din_startofpacket
	wire   [23:0] alt_vip_crs_0_dout_data;                                       // alt_vip_crs_0:dout_data -> alt_vip_csc_0:din_data
	wire          alt_vip_crs_0_dout_ready;                                      // alt_vip_csc_0:din_ready -> alt_vip_crs_0:dout_ready
	wire          alt_vip_csc_0_dout_endofpacket;                                // alt_vip_csc_0:dout_endofpacket -> alt_vip_clip_0:din_endofpacket
	wire          alt_vip_csc_0_dout_valid;                                      // alt_vip_csc_0:dout_valid -> alt_vip_clip_0:din_valid
	wire          alt_vip_csc_0_dout_startofpacket;                              // alt_vip_csc_0:dout_startofpacket -> alt_vip_clip_0:din_startofpacket
	wire   [23:0] alt_vip_csc_0_dout_data;                                       // alt_vip_csc_0:dout_data -> alt_vip_clip_0:din_data
	wire          alt_vip_csc_0_dout_ready;                                      // alt_vip_clip_0:din_ready -> alt_vip_csc_0:dout_ready
	wire          pll_sys_outclk2_clk;                                           // pll_sys:outclk_2 -> [clock_crossing_io_slow:m0_clk, i2c_scl:clk, i2c_sda:clk, irq_synchronizer:receiver_clk, key:clk, ledr:clk, mm_interconnect_0:pll_sys_outclk2_clk, mm_interconnect_2:pll_sys_outclk2_clk, rst_controller:clk, seg7:s_clk, sw:clk, sysid:clock, td_reset_n:clk, td_status:clk, timer:clk]
	wire          pll_sys_outclk0_clk;                                           // pll_sys:outclk_0 -> [alt_vip_cl_scl_0:main_clock, alt_vip_clip_0:clock, alt_vip_cpr_0:clock, alt_vip_cpr_1:clock, alt_vip_cpr_2:clock, alt_vip_crs_0:clock, alt_vip_csc_0:clock, alt_vip_cti_0:is_clk, alt_vip_dil_0:clock, alt_vip_itc_0:is_clk, alt_vip_mix_0:clock, alt_vip_vfb_0:clock, alt_vip_vfr_0:clock, alt_vip_vfr_0:master_clock, clock_crossing_io_slow:s0_clk, cpu:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_clock_crossing_bridge_1:s0_clk, mm_interconnect_0:pll_sys_outclk0_clk, mm_interconnect_1:pll_sys_outclk0_clk, mm_interconnect_4:pll_sys_outclk0_clk, onchip_memory2:clk, rst_controller_001:clk, rst_controller_002:clk, sdram:clk, timer_stamp:clk, uart:clk]
	wire          pll_audio_outclk0_clk;                                         // pll_audio:outclk_0 -> [audio:avs_s1_clk, mm_interconnect_0:pll_audio_outclk0_clk, rst_controller_005:clk]
	wire          pll_sys_outclk4_clk;                                           // pll_sys:outclk_4 -> [irq_synchronizer_001:receiver_clk, mm_clock_crossing_bridge_1:m0_clk, mm_interconnect_3:pll_sys_outclk4_clk, rst_controller_004:clk, spi_0:clk]
	wire          alt_vip_dil_0_dout_endofpacket;                                // alt_vip_dil_0:dout_endofpacket -> alt_vip_crs_0:din_endofpacket
	wire          alt_vip_dil_0_dout_valid;                                      // alt_vip_dil_0:dout_valid -> alt_vip_crs_0:din_valid
	wire          alt_vip_dil_0_dout_startofpacket;                              // alt_vip_dil_0:dout_startofpacket -> alt_vip_crs_0:din_startofpacket
	wire   [15:0] alt_vip_dil_0_dout_data;                                       // alt_vip_dil_0:dout_data -> alt_vip_crs_0:din_data
	wire          alt_vip_dil_0_dout_ready;                                      // alt_vip_crs_0:din_ready -> alt_vip_dil_0:dout_ready
	wire          alt_vip_cl_scl_0_dout_endofpacket;                             // alt_vip_cl_scl_0:dout_endofpacket -> alt_vip_vfb_0:din_endofpacket
	wire          alt_vip_cl_scl_0_dout_valid;                                   // alt_vip_cl_scl_0:dout_valid -> alt_vip_vfb_0:din_valid
	wire          alt_vip_cl_scl_0_dout_startofpacket;                           // alt_vip_cl_scl_0:dout_startofpacket -> alt_vip_vfb_0:din_startofpacket
	wire   [23:0] alt_vip_cl_scl_0_dout_data;                                    // alt_vip_cl_scl_0:dout_data -> alt_vip_vfb_0:din_data
	wire          alt_vip_cl_scl_0_dout_ready;                                   // alt_vip_vfb_0:din_ready -> alt_vip_cl_scl_0:dout_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;             // alt_vip_vfr_0:dout_endofpacket -> alt_vip_cpr_1:din0_endofpacket
	wire          alt_vip_vfr_0_avalon_streaming_source_valid;                   // alt_vip_vfr_0:dout_valid -> alt_vip_cpr_1:din0_valid
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;           // alt_vip_vfr_0:dout_startofpacket -> alt_vip_cpr_1:din0_startofpacket
	wire   [31:0] alt_vip_vfr_0_avalon_streaming_source_data;                    // alt_vip_vfr_0:dout_data -> alt_vip_cpr_1:din0_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;                   // alt_vip_cpr_1:din0_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_mix_0_dout_endofpacket;                                // alt_vip_mix_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          alt_vip_mix_0_dout_valid;                                      // alt_vip_mix_0:dout_valid -> alt_vip_itc_0:is_valid
	wire          alt_vip_mix_0_dout_startofpacket;                              // alt_vip_mix_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire   [23:0] alt_vip_mix_0_dout_data;                                       // alt_vip_mix_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_mix_0_dout_ready;                                      // alt_vip_itc_0:is_ready -> alt_vip_mix_0:dout_ready
	wire          alt_vip_vfb_0_dout_endofpacket;                                // alt_vip_vfb_0:dout_endofpacket -> alt_vip_cpr_2:din0_endofpacket
	wire          alt_vip_vfb_0_dout_valid;                                      // alt_vip_vfb_0:dout_valid -> alt_vip_cpr_2:din0_valid
	wire          alt_vip_vfb_0_dout_startofpacket;                              // alt_vip_vfb_0:dout_startofpacket -> alt_vip_cpr_2:din0_startofpacket
	wire   [23:0] alt_vip_vfb_0_dout_data;                                       // alt_vip_vfb_0:dout_data -> alt_vip_cpr_2:din0_data
	wire          alt_vip_vfb_0_dout_ready;                                      // alt_vip_cpr_2:din0_ready -> alt_vip_vfb_0:dout_ready
	wire          alt_vip_cpr_1_dout0_endofpacket;                               // alt_vip_cpr_1:dout0_endofpacket -> alt_vip_mix_0:din_0_endofpacket
	wire          alt_vip_cpr_1_dout0_valid;                                     // alt_vip_cpr_1:dout0_valid -> alt_vip_mix_0:din_0_valid
	wire          alt_vip_cpr_1_dout0_startofpacket;                             // alt_vip_cpr_1:dout0_startofpacket -> alt_vip_mix_0:din_0_startofpacket
	wire   [23:0] alt_vip_cpr_1_dout0_data;                                      // alt_vip_cpr_1:dout0_data -> alt_vip_mix_0:din_0_data
	wire          alt_vip_cpr_1_dout0_ready;                                     // alt_vip_mix_0:din_0_ready -> alt_vip_cpr_1:dout0_ready
	wire          alt_vip_cpr_2_dout0_endofpacket;                               // alt_vip_cpr_2:dout0_endofpacket -> alt_vip_mix_0:din_1_endofpacket
	wire          alt_vip_cpr_2_dout0_valid;                                     // alt_vip_cpr_2:dout0_valid -> alt_vip_mix_0:din_1_valid
	wire          alt_vip_cpr_2_dout0_startofpacket;                             // alt_vip_cpr_2:dout0_startofpacket -> alt_vip_mix_0:din_1_startofpacket
	wire   [23:0] alt_vip_cpr_2_dout0_data;                                      // alt_vip_cpr_2:dout0_data -> alt_vip_mix_0:din_1_data
	wire          alt_vip_cpr_2_dout0_ready;                                     // alt_vip_mix_0:din_1_ready -> alt_vip_cpr_2:dout0_ready
	wire   [31:0] mm_interconnect_0_ir_rx_avalon_slave_writedata;                // mm_interconnect_0:ir_rx_avalon_slave_writedata -> ir_rx:s_writedata
	wire    [0:0] mm_interconnect_0_ir_rx_avalon_slave_address;                  // mm_interconnect_0:ir_rx_avalon_slave_address -> ir_rx:s_address
	wire          mm_interconnect_0_ir_rx_avalon_slave_chipselect;               // mm_interconnect_0:ir_rx_avalon_slave_chipselect -> ir_rx:s_cs_n
	wire          mm_interconnect_0_ir_rx_avalon_slave_write;                    // mm_interconnect_0:ir_rx_avalon_slave_write -> ir_rx:s_write
	wire          mm_interconnect_0_ir_rx_avalon_slave_read;                     // mm_interconnect_0:ir_rx_avalon_slave_read -> ir_rx:s_read
	wire   [31:0] mm_interconnect_0_ir_rx_avalon_slave_readdata;                 // ir_rx:s_readdata -> mm_interconnect_0:ir_rx_avalon_slave_readdata
	wire   [31:0] mm_interconnect_0_sw_s1_writedata;                             // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire    [1:0] mm_interconnect_0_sw_s1_address;                               // mm_interconnect_0:sw_s1_address -> sw:address
	wire          mm_interconnect_0_sw_s1_chipselect;                            // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire          mm_interconnect_0_sw_s1_write;                                 // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire   [31:0] mm_interconnect_0_sw_s1_readdata;                              // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_writedata;                // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire    [2:0] mm_interconnect_0_audio_avalon_slave_address;                  // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire          mm_interconnect_0_audio_avalon_slave_write;                    // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire          mm_interconnect_0_audio_avalon_slave_read;                     // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_readdata;                 // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire   [31:0] mm_interconnect_0_ledr_s1_writedata;                           // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire    [1:0] mm_interconnect_0_ledr_s1_address;                             // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire          mm_interconnect_0_ledr_s1_chipselect;                          // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire          mm_interconnect_0_ledr_s1_write;                               // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire   [31:0] mm_interconnect_0_ledr_s1_readdata;                            // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [15:0] mm_interconnect_0_alt_vip_cti_0_control_writedata;             // mm_interconnect_0:alt_vip_cti_0_control_writedata -> alt_vip_cti_0:av_writedata
	wire    [3:0] mm_interconnect_0_alt_vip_cti_0_control_address;               // mm_interconnect_0:alt_vip_cti_0_control_address -> alt_vip_cti_0:av_address
	wire          mm_interconnect_0_alt_vip_cti_0_control_write;                 // mm_interconnect_0:alt_vip_cti_0_control_write -> alt_vip_cti_0:av_write
	wire          mm_interconnect_0_alt_vip_cti_0_control_read;                  // mm_interconnect_0:alt_vip_cti_0_control_read -> alt_vip_cti_0:av_read
	wire   [15:0] mm_interconnect_0_alt_vip_cti_0_control_readdata;              // alt_vip_cti_0:av_readdata -> mm_interconnect_0:alt_vip_cti_0_control_readdata
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                 // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire   [15:0] mm_interconnect_0_onchip_memory2_s1_address;                   // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire          mm_interconnect_0_onchip_memory2_s1_chipselect;                // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire          mm_interconnect_0_onchip_memory2_s1_clken;                     // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire          mm_interconnect_0_onchip_memory2_s1_write;                     // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                  // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire    [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire   [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata;        // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire    [4:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address;          // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire          mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write;            // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire          mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read;             // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire   [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata;         // alt_vip_vfr_0:slave_readdata -> mm_interconnect_0:alt_vip_vfr_0_avalon_slave_readdata
	wire   [15:0] mm_interconnect_0_uart_s1_writedata;                           // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire    [2:0] mm_interconnect_0_uart_s1_address;                             // mm_interconnect_0:uart_s1_address -> uart:address
	wire          mm_interconnect_0_uart_s1_chipselect;                          // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire          mm_interconnect_0_uart_s1_write;                               // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire          mm_interconnect_0_uart_s1_read;                                // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire   [15:0] mm_interconnect_0_uart_s1_readdata;                            // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire          mm_interconnect_0_uart_s1_begintransfer;                       // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire   [15:0] mm_interconnect_0_alt_vip_mix_0_control_writedata;             // mm_interconnect_0:alt_vip_mix_0_control_writedata -> alt_vip_mix_0:control_av_writedata
	wire    [5:0] mm_interconnect_0_alt_vip_mix_0_control_address;               // mm_interconnect_0:alt_vip_mix_0_control_address -> alt_vip_mix_0:control_av_address
	wire          mm_interconnect_0_alt_vip_mix_0_control_chipselect;            // mm_interconnect_0:alt_vip_mix_0_control_chipselect -> alt_vip_mix_0:control_av_chipselect
	wire          mm_interconnect_0_alt_vip_mix_0_control_write;                 // mm_interconnect_0:alt_vip_mix_0_control_write -> alt_vip_mix_0:control_av_write
	wire   [15:0] mm_interconnect_0_alt_vip_mix_0_control_readdata;              // alt_vip_mix_0:control_av_readdata -> mm_interconnect_0:alt_vip_mix_0_control_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire   [15:0] mm_interconnect_0_timer_stamp_s1_writedata;                    // mm_interconnect_0:timer_stamp_s1_writedata -> timer_stamp:writedata
	wire    [2:0] mm_interconnect_0_timer_stamp_s1_address;                      // mm_interconnect_0:timer_stamp_s1_address -> timer_stamp:address
	wire          mm_interconnect_0_timer_stamp_s1_chipselect;                   // mm_interconnect_0:timer_stamp_s1_chipselect -> timer_stamp:chipselect
	wire          mm_interconnect_0_timer_stamp_s1_write;                        // mm_interconnect_0:timer_stamp_s1_write -> timer_stamp:write_n
	wire   [15:0] mm_interconnect_0_timer_stamp_s1_readdata;                     // timer_stamp:readdata -> mm_interconnect_0:timer_stamp_s1_readdata
	wire    [7:0] mm_interconnect_0_seg7_avalon_slave_writedata;                 // mm_interconnect_0:seg7_avalon_slave_writedata -> seg7:s_writedata
	wire    [2:0] mm_interconnect_0_seg7_avalon_slave_address;                   // mm_interconnect_0:seg7_avalon_slave_address -> seg7:s_address
	wire          mm_interconnect_0_seg7_avalon_slave_write;                     // mm_interconnect_0:seg7_avalon_slave_write -> seg7:s_write
	wire          mm_interconnect_0_seg7_avalon_slave_read;                      // mm_interconnect_0:seg7_avalon_slave_read -> seg7:s_read
	wire    [7:0] mm_interconnect_0_seg7_avalon_slave_readdata;                  // seg7:s_readdata -> mm_interconnect_0:seg7_avalon_slave_readdata
	wire   [31:0] mm_interconnect_0_key_s1_writedata;                            // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire    [1:0] mm_interconnect_0_key_s1_address;                              // mm_interconnect_0:key_s1_address -> key:address
	wire          mm_interconnect_0_key_s1_chipselect;                           // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire          mm_interconnect_0_key_s1_write;                                // mm_interconnect_0:key_s1_write -> key:write_n
	wire   [31:0] mm_interconnect_0_key_s1_readdata;                             // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire          mm_interconnect_0_cpu_jtag_debug_module_waitrequest;           // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire   [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;             // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;               // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire          mm_interconnect_0_cpu_jtag_debug_module_write;                 // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire          mm_interconnect_0_cpu_jtag_debug_module_read;                  // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;              // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire          mm_interconnect_0_cpu_jtag_debug_module_debugaccess;           // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;            // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire          hps_0_h2f_lw_axi_master_awvalid;                               // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                               // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire          hps_0_h2f_lw_axi_master_arready;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                  // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire          hps_0_h2f_lw_axi_master_rready;                                // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire          hps_0_h2f_lw_axi_master_bready;                                // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire          hps_0_h2f_lw_axi_master_arvalid;                               // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                 // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire          hps_0_h2f_lw_axi_master_awready;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                  // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire          hps_0_h2f_lw_axi_master_bvalid;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                   // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                               // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                 // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_rvalid;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                 // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_wready;                                // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                               // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                               // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                 // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_wvalid;                                // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire          hps_0_h2f_lw_axi_master_wlast;                                 // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire          hps_0_h2f_lw_axi_master_rlast;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          cpu_instruction_master_waitrequest;                            // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire   [19:0] cpu_instruction_master_address;                                // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire          cpu_instruction_master_read;                                   // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire   [31:0] cpu_instruction_master_readdata;                               // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                          // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire          mm_interconnect_0_clock_crossing_io_slow_s0_waitrequest;       // clock_crossing_io_slow:s0_waitrequest -> mm_interconnect_0:clock_crossing_io_slow_s0_waitrequest
	wire    [0:0] mm_interconnect_0_clock_crossing_io_slow_s0_burstcount;        // mm_interconnect_0:clock_crossing_io_slow_s0_burstcount -> clock_crossing_io_slow:s0_burstcount
	wire   [31:0] mm_interconnect_0_clock_crossing_io_slow_s0_writedata;         // mm_interconnect_0:clock_crossing_io_slow_s0_writedata -> clock_crossing_io_slow:s0_writedata
	wire    [8:0] mm_interconnect_0_clock_crossing_io_slow_s0_address;           // mm_interconnect_0:clock_crossing_io_slow_s0_address -> clock_crossing_io_slow:s0_address
	wire          mm_interconnect_0_clock_crossing_io_slow_s0_write;             // mm_interconnect_0:clock_crossing_io_slow_s0_write -> clock_crossing_io_slow:s0_write
	wire          mm_interconnect_0_clock_crossing_io_slow_s0_read;              // mm_interconnect_0:clock_crossing_io_slow_s0_read -> clock_crossing_io_slow:s0_read
	wire   [31:0] mm_interconnect_0_clock_crossing_io_slow_s0_readdata;          // clock_crossing_io_slow:s0_readdata -> mm_interconnect_0:clock_crossing_io_slow_s0_readdata
	wire          mm_interconnect_0_clock_crossing_io_slow_s0_debugaccess;       // mm_interconnect_0:clock_crossing_io_slow_s0_debugaccess -> clock_crossing_io_slow:s0_debugaccess
	wire          mm_interconnect_0_clock_crossing_io_slow_s0_readdatavalid;     // clock_crossing_io_slow:s0_readdatavalid -> mm_interconnect_0:clock_crossing_io_slow_s0_readdatavalid
	wire    [3:0] mm_interconnect_0_clock_crossing_io_slow_s0_byteenable;        // mm_interconnect_0:clock_crossing_io_slow_s0_byteenable -> clock_crossing_io_slow:s0_byteenable
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest;   // mm_clock_crossing_bridge_1:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_waitrequest
	wire    [0:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_burstcount -> mm_clock_crossing_bridge_1:s0_burstcount
	wire   [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_writedata -> mm_clock_crossing_bridge_1:s0_writedata
	wire    [8:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_address -> mm_clock_crossing_bridge_1:s0_address
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_write -> mm_clock_crossing_bridge_1:s0_write
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_read -> mm_clock_crossing_bridge_1:s0_read
	wire   [31:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata;      // mm_clock_crossing_bridge_1:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdata
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_debugaccess -> mm_clock_crossing_bridge_1:s0_debugaccess
	wire          mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid; // mm_clock_crossing_bridge_1:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_1_s0_readdatavalid
	wire    [3:0] mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_1_s0_byteenable -> mm_clock_crossing_bridge_1:s0_byteenable
	wire          cpu_data_master_waitrequest;                                   // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                     // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire   [25:0] cpu_data_master_address;                                       // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire          cpu_data_master_write;                                         // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire          cpu_data_master_read;                                          // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire   [31:0] cpu_data_master_readdata;                                      // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                   // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire          cpu_data_master_readdatavalid;                                 // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                    // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire    [2:0] alt_vip_vfb_0_write_master_burstcount;                         // alt_vip_vfb_0:write_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_write_master_burstcount
	wire          alt_vip_vfb_0_write_master_waitrequest;                        // mm_interconnect_1:alt_vip_vfb_0_write_master_waitrequest -> alt_vip_vfb_0:write_master_av_waitrequest
	wire   [31:0] alt_vip_vfb_0_write_master_writedata;                          // alt_vip_vfb_0:write_master_av_writedata -> mm_interconnect_1:alt_vip_vfb_0_write_master_writedata
	wire   [31:0] alt_vip_vfb_0_write_master_address;                            // alt_vip_vfb_0:write_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_write_master_address
	wire          alt_vip_vfb_0_write_master_write;                              // alt_vip_vfb_0:write_master_av_write -> mm_interconnect_1:alt_vip_vfb_0_write_master_write
	wire          mm_interconnect_1_sdram_s1_waitrequest;                        // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire   [15:0] mm_interconnect_1_sdram_s1_writedata;                          // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire   [24:0] mm_interconnect_1_sdram_s1_address;                            // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_1_sdram_s1_chipselect;                         // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire          mm_interconnect_1_sdram_s1_write;                              // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire          mm_interconnect_1_sdram_s1_read;                               // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire   [15:0] mm_interconnect_1_sdram_s1_readdata;                           // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire          mm_interconnect_1_sdram_s1_readdatavalid;                      // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire    [1:0] mm_interconnect_1_sdram_s1_byteenable;                         // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire    [2:0] alt_vip_vfb_0_read_master_burstcount;                          // alt_vip_vfb_0:read_master_av_burstcount -> mm_interconnect_1:alt_vip_vfb_0_read_master_burstcount
	wire          alt_vip_vfb_0_read_master_waitrequest;                         // mm_interconnect_1:alt_vip_vfb_0_read_master_waitrequest -> alt_vip_vfb_0:read_master_av_waitrequest
	wire   [31:0] alt_vip_vfb_0_read_master_address;                             // alt_vip_vfb_0:read_master_av_address -> mm_interconnect_1:alt_vip_vfb_0_read_master_address
	wire          alt_vip_vfb_0_read_master_read;                                // alt_vip_vfb_0:read_master_av_read -> mm_interconnect_1:alt_vip_vfb_0_read_master_read
	wire   [31:0] alt_vip_vfb_0_read_master_readdata;                            // mm_interconnect_1:alt_vip_vfb_0_read_master_readdata -> alt_vip_vfb_0:read_master_av_readdata
	wire          alt_vip_vfb_0_read_master_readdatavalid;                       // mm_interconnect_1:alt_vip_vfb_0_read_master_readdatavalid -> alt_vip_vfb_0:read_master_av_readdatavalid
	wire   [31:0] mm_interconnect_2_td_reset_n_s1_writedata;                     // mm_interconnect_2:td_reset_n_s1_writedata -> td_reset_n:writedata
	wire    [1:0] mm_interconnect_2_td_reset_n_s1_address;                       // mm_interconnect_2:td_reset_n_s1_address -> td_reset_n:address
	wire          mm_interconnect_2_td_reset_n_s1_chipselect;                    // mm_interconnect_2:td_reset_n_s1_chipselect -> td_reset_n:chipselect
	wire          mm_interconnect_2_td_reset_n_s1_write;                         // mm_interconnect_2:td_reset_n_s1_write -> td_reset_n:write_n
	wire   [31:0] mm_interconnect_2_td_reset_n_s1_readdata;                      // td_reset_n:readdata -> mm_interconnect_2:td_reset_n_s1_readdata
	wire   [31:0] mm_interconnect_2_i2c_scl_s1_writedata;                        // mm_interconnect_2:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire    [1:0] mm_interconnect_2_i2c_scl_s1_address;                          // mm_interconnect_2:i2c_scl_s1_address -> i2c_scl:address
	wire          mm_interconnect_2_i2c_scl_s1_chipselect;                       // mm_interconnect_2:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire          mm_interconnect_2_i2c_scl_s1_write;                            // mm_interconnect_2:i2c_scl_s1_write -> i2c_scl:write_n
	wire   [31:0] mm_interconnect_2_i2c_scl_s1_readdata;                         // i2c_scl:readdata -> mm_interconnect_2:i2c_scl_s1_readdata
	wire    [1:0] mm_interconnect_2_td_status_s1_address;                        // mm_interconnect_2:td_status_s1_address -> td_status:address
	wire   [31:0] mm_interconnect_2_td_status_s1_readdata;                       // td_status:readdata -> mm_interconnect_2:td_status_s1_readdata
	wire   [31:0] mm_interconnect_2_i2c_sda_s1_writedata;                        // mm_interconnect_2:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire    [1:0] mm_interconnect_2_i2c_sda_s1_address;                          // mm_interconnect_2:i2c_sda_s1_address -> i2c_sda:address
	wire          mm_interconnect_2_i2c_sda_s1_chipselect;                       // mm_interconnect_2:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire          mm_interconnect_2_i2c_sda_s1_write;                            // mm_interconnect_2:i2c_sda_s1_write -> i2c_sda:write_n
	wire   [31:0] mm_interconnect_2_i2c_sda_s1_readdata;                         // i2c_sda:readdata -> mm_interconnect_2:i2c_sda_s1_readdata
	wire   [15:0] mm_interconnect_2_timer_s1_writedata;                          // mm_interconnect_2:timer_s1_writedata -> timer:writedata
	wire    [2:0] mm_interconnect_2_timer_s1_address;                            // mm_interconnect_2:timer_s1_address -> timer:address
	wire          mm_interconnect_2_timer_s1_chipselect;                         // mm_interconnect_2:timer_s1_chipselect -> timer:chipselect
	wire          mm_interconnect_2_timer_s1_write;                              // mm_interconnect_2:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_2_timer_s1_readdata;                           // timer:readdata -> mm_interconnect_2:timer_s1_readdata
	wire    [0:0] mm_interconnect_2_sysid_control_slave_address;                 // mm_interconnect_2:sysid_control_slave_address -> sysid:address
	wire   [31:0] mm_interconnect_2_sysid_control_slave_readdata;                // sysid:readdata -> mm_interconnect_2:sysid_control_slave_readdata
	wire    [0:0] clock_crossing_io_slow_m0_burstcount;                          // clock_crossing_io_slow:m0_burstcount -> mm_interconnect_2:clock_crossing_io_slow_m0_burstcount
	wire          clock_crossing_io_slow_m0_waitrequest;                         // mm_interconnect_2:clock_crossing_io_slow_m0_waitrequest -> clock_crossing_io_slow:m0_waitrequest
	wire    [8:0] clock_crossing_io_slow_m0_address;                             // clock_crossing_io_slow:m0_address -> mm_interconnect_2:clock_crossing_io_slow_m0_address
	wire   [31:0] clock_crossing_io_slow_m0_writedata;                           // clock_crossing_io_slow:m0_writedata -> mm_interconnect_2:clock_crossing_io_slow_m0_writedata
	wire          clock_crossing_io_slow_m0_write;                               // clock_crossing_io_slow:m0_write -> mm_interconnect_2:clock_crossing_io_slow_m0_write
	wire          clock_crossing_io_slow_m0_read;                                // clock_crossing_io_slow:m0_read -> mm_interconnect_2:clock_crossing_io_slow_m0_read
	wire   [31:0] clock_crossing_io_slow_m0_readdata;                            // mm_interconnect_2:clock_crossing_io_slow_m0_readdata -> clock_crossing_io_slow:m0_readdata
	wire          clock_crossing_io_slow_m0_debugaccess;                         // clock_crossing_io_slow:m0_debugaccess -> mm_interconnect_2:clock_crossing_io_slow_m0_debugaccess
	wire    [3:0] clock_crossing_io_slow_m0_byteenable;                          // clock_crossing_io_slow:m0_byteenable -> mm_interconnect_2:clock_crossing_io_slow_m0_byteenable
	wire          clock_crossing_io_slow_m0_readdatavalid;                       // mm_interconnect_2:clock_crossing_io_slow_m0_readdatavalid -> clock_crossing_io_slow:m0_readdatavalid
	wire    [0:0] mm_clock_crossing_bridge_1_m0_burstcount;                      // mm_clock_crossing_bridge_1:m0_burstcount -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_burstcount
	wire          mm_clock_crossing_bridge_1_m0_waitrequest;                     // mm_interconnect_3:mm_clock_crossing_bridge_1_m0_waitrequest -> mm_clock_crossing_bridge_1:m0_waitrequest
	wire    [8:0] mm_clock_crossing_bridge_1_m0_address;                         // mm_clock_crossing_bridge_1:m0_address -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_address
	wire   [31:0] mm_clock_crossing_bridge_1_m0_writedata;                       // mm_clock_crossing_bridge_1:m0_writedata -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_writedata
	wire          mm_clock_crossing_bridge_1_m0_write;                           // mm_clock_crossing_bridge_1:m0_write -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_write
	wire          mm_clock_crossing_bridge_1_m0_read;                            // mm_clock_crossing_bridge_1:m0_read -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_read
	wire   [31:0] mm_clock_crossing_bridge_1_m0_readdata;                        // mm_interconnect_3:mm_clock_crossing_bridge_1_m0_readdata -> mm_clock_crossing_bridge_1:m0_readdata
	wire          mm_clock_crossing_bridge_1_m0_debugaccess;                     // mm_clock_crossing_bridge_1:m0_debugaccess -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_debugaccess
	wire    [3:0] mm_clock_crossing_bridge_1_m0_byteenable;                      // mm_clock_crossing_bridge_1:m0_byteenable -> mm_interconnect_3:mm_clock_crossing_bridge_1_m0_byteenable
	wire          mm_clock_crossing_bridge_1_m0_readdatavalid;                   // mm_interconnect_3:mm_clock_crossing_bridge_1_m0_readdatavalid -> mm_clock_crossing_bridge_1:m0_readdatavalid
	wire   [15:0] mm_interconnect_3_spi_0_spi_control_port_writedata;            // mm_interconnect_3:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire    [2:0] mm_interconnect_3_spi_0_spi_control_port_address;              // mm_interconnect_3:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire          mm_interconnect_3_spi_0_spi_control_port_chipselect;           // mm_interconnect_3:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire          mm_interconnect_3_spi_0_spi_control_port_write;                // mm_interconnect_3:spi_0_spi_control_port_write -> spi_0:write_n
	wire          mm_interconnect_3_spi_0_spi_control_port_read;                 // mm_interconnect_3:spi_0_spi_control_port_read -> spi_0:read_n
	wire   [15:0] mm_interconnect_3_spi_0_spi_control_port_readdata;             // spi_0:data_to_cpu -> mm_interconnect_3:spi_0_spi_control_port_readdata
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_awvalid;                 // mm_interconnect_4:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_arsize;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_arlock;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_awcache;                 // mm_interconnect_4:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_arready;                 // hps_0:f2h_ARREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_arready
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_arid;                    // mm_interconnect_4:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rready;                  // mm_interconnect_4:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_bready;                  // mm_interconnect_4:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_awsize;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_awprot;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_arvalid;                 // mm_interconnect_4:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [2:0] mm_interconnect_4_hps_0_f2h_axi_slave_arprot;                  // mm_interconnect_4:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_bid;                     // hps_0:f2h_BID -> mm_interconnect_4:hps_0_f2h_axi_slave_bid
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_arlen;                   // mm_interconnect_4:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_awready;                 // hps_0:f2h_AWREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_awready
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_awid;                    // mm_interconnect_4:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_bvalid;                  // hps_0:f2h_BVALID -> mm_interconnect_4:hps_0_f2h_axi_slave_bvalid
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_wid;                     // mm_interconnect_4:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_awlock;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_awburst;                 // mm_interconnect_4:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_bresp;                   // hps_0:f2h_BRESP -> mm_interconnect_4:hps_0_f2h_axi_slave_bresp
	wire    [4:0] mm_interconnect_4_hps_0_f2h_axi_slave_aruser;                  // mm_interconnect_4:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire    [4:0] mm_interconnect_4_hps_0_f2h_axi_slave_awuser;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire   [15:0] mm_interconnect_4_hps_0_f2h_axi_slave_wstrb;                   // mm_interconnect_4:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rvalid;                  // hps_0:f2h_RVALID -> mm_interconnect_4:hps_0_f2h_axi_slave_rvalid
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_arburst;                 // mm_interconnect_4:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire  [127:0] mm_interconnect_4_hps_0_f2h_axi_slave_wdata;                   // mm_interconnect_4:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wready;                  // hps_0:f2h_WREADY -> mm_interconnect_4:hps_0_f2h_axi_slave_wready
	wire  [127:0] mm_interconnect_4_hps_0_f2h_axi_slave_rdata;                   // hps_0:f2h_RDATA -> mm_interconnect_4:hps_0_f2h_axi_slave_rdata
	wire   [31:0] mm_interconnect_4_hps_0_f2h_axi_slave_araddr;                  // mm_interconnect_4:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_arcache;                 // mm_interconnect_4:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire    [3:0] mm_interconnect_4_hps_0_f2h_axi_slave_awlen;                   // mm_interconnect_4:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [31:0] mm_interconnect_4_hps_0_f2h_axi_slave_awaddr;                  // mm_interconnect_4:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [7:0] mm_interconnect_4_hps_0_f2h_axi_slave_rid;                     // hps_0:f2h_RID -> mm_interconnect_4:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wvalid;                  // mm_interconnect_4:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire    [1:0] mm_interconnect_4_hps_0_f2h_axi_slave_rresp;                   // hps_0:f2h_RRESP -> mm_interconnect_4:hps_0_f2h_axi_slave_rresp
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_wlast;                   // mm_interconnect_4:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire          mm_interconnect_4_hps_0_f2h_axi_slave_rlast;                   // hps_0:f2h_RLAST -> mm_interconnect_4:hps_0_f2h_axi_slave_rlast
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                       // mm_interconnect_4:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire    [5:0] alt_vip_vfr_0_avalon_master_burstcount;                        // alt_vip_vfr_0:master_burstcount -> mm_interconnect_4:alt_vip_vfr_0_avalon_master_burstcount
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                           // alt_vip_vfr_0:master_address -> mm_interconnect_4:alt_vip_vfr_0_avalon_master_address
	wire          alt_vip_vfr_0_avalon_master_read;                              // alt_vip_vfr_0:master_read -> mm_interconnect_4:alt_vip_vfr_0_avalon_master_read
	wire  [127:0] alt_vip_vfr_0_avalon_master_readdata;                          // mm_interconnect_4:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;                     // mm_interconnect_4:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire          irq_mapper_receiver1_irq;                                      // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                      // uart:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver4_irq;                                      // timer_stamp:irq -> irq_mapper:receiver4_irq
	wire   [31:0] cpu_d_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:d_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                            // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                            // irq_mapper_002:sender_irq -> hps_0:f2h_irq_p1
	wire          irq_mapper_receiver0_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                 // timer:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver3_irq;                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                             // spi_0:irq -> irq_synchronizer_001:receiver_irq
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [clock_crossing_io_slow:m0_reset, i2c_scl:reset_n, i2c_sda:reset_n, irq_synchronizer:receiver_reset, key:reset_n, ledr:reset_n, mm_interconnect_0:ledr_reset_reset_bridge_in_reset_reset, mm_interconnect_2:clock_crossing_io_slow_m0_reset_reset_bridge_in_reset_reset, seg7:s_reset, sw:reset_n, sysid:reset_n, td_reset_n:reset_n, td_status:reset_n, timer:reset_n]
	wire          rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:onchip_memory2_reset1_reset_bridge_in_reset_reset, onchip_memory2:reset]
	wire          rst_controller_001_reset_out_reset_req;                        // rst_controller_001:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire          cpu_jtag_debug_module_reset_reset;                             // cpu:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	wire          rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [alt_vip_cl_scl_0:main_reset, alt_vip_clip_0:reset, alt_vip_cpr_0:reset, alt_vip_cpr_1:reset, alt_vip_cpr_2:reset, alt_vip_crs_0:reset, alt_vip_csc_0:reset, alt_vip_cti_0:rst, alt_vip_dil_0:reset, alt_vip_itc_0:rst, alt_vip_mix_0:reset, alt_vip_vfb_0:reset, alt_vip_vfr_0:master_reset, alt_vip_vfr_0:reset, clock_crossing_io_slow:s0_reset, cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_clock_crossing_bridge_1:s0_reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:alt_vip_vfb_0_reset_reset_bridge_in_reset_reset, mm_interconnect_4:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, sdram:reset_n, timer_stamp:reset_n, uart:reset_n]
	wire          rst_controller_002_reset_out_reset_req;                        // rst_controller_002:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_003_reset_out_reset;                            // rst_controller_003:reset_out -> [ir_rx:reset_n, mm_interconnect_0:ir_rx_clock_sink_reset_reset_bridge_in_reset_reset, pll_audio:rst, pll_sys:rst]
	wire          rst_controller_004_reset_out_reset;                            // rst_controller_004:reset_out -> [irq_synchronizer_001:receiver_reset, mm_clock_crossing_bridge_1:m0_reset, mm_interconnect_3:mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset, spi_0:reset_n]
	wire          rst_controller_005_reset_out_reset;                            // rst_controller_005:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_clock_sink_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_006_reset_out_reset;                            // rst_controller_006:reset_out -> [mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_4:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	DE1_SoC_QSYS_timer timer (
		.clk        (pll_sys_outclk2_clk),                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_2_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_2_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_2_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_2_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_2_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	DE1_SoC_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (pll_sys_outclk0_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)          //       .reset_req
	);

	DE1_SoC_QSYS_sdram sdram (
		.clk            (pll_sys_outclk0_clk),                      //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                   //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                     //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                  //      .export
		.zs_cke         (zs_cke_from_the_sdram),                    //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                   //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),              //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                    //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                  //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                    //      .export
	);

	DE1_SoC_QSYS_i2c_scl i2c_scl (
		.clk        (pll_sys_outclk2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_i2c_scl)                // external_connection.export
	);

	DE1_SoC_QSYS_i2c_sda i2c_sda (
		.clk        (pll_sys_outclk2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_i2c_sda)       // external_connection.export
	);

	DE1_SoC_QSYS_jtag_uart jtag_uart (
		.clk            (pll_sys_outclk0_clk),                                       //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	alt_vipcti131_Vid2IS #(
		.BPS                           (8),
		.NUMBER_OF_COLOUR_PLANES       (2),
		.COLOUR_PLANES_ARE_IN_PARALLEL (0),
		.SYNC_TO                       (0),
		.USE_EMBEDDED_SYNCS            (1),
		.ADD_DATA_ENABLE_SIGNAL        (0),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.USE_STD                       (0),
		.STD_WIDTH                     (1),
		.GENERATE_ANC                  (0),
		.INTERLACED                    (1),
		.H_ACTIVE_PIXELS_F0            (720),
		.V_ACTIVE_LINES_F0             (288),
		.V_ACTIVE_LINES_F1             (288),
		.FIFO_DEPTH                    (1440),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (1),
		.GENERATE_SYNC                 (0)
	) alt_vip_cti_0 (
		.is_clk            (pll_sys_outclk0_clk),                               //        is_clk_rst.clk
		.rst               (rst_controller_002_reset_out_reset),                //  is_clk_rst_reset.reset
		.av_address        (mm_interconnect_0_alt_vip_cti_0_control_address),   //           control.address
		.av_read           (mm_interconnect_0_alt_vip_cti_0_control_read),      //                  .read
		.av_readdata       (mm_interconnect_0_alt_vip_cti_0_control_readdata),  //                  .readdata
		.av_write          (mm_interconnect_0_alt_vip_cti_0_control_write),     //                  .write
		.av_writedata      (mm_interconnect_0_alt_vip_cti_0_control_writedata), //                  .writedata
		.status_update_int (),                                                  // status_update_irq.irq
		.is_data           (alt_vip_cti_0_dout_data),                           //              dout.data
		.is_valid          (alt_vip_cti_0_dout_valid),                          //                  .valid
		.is_ready          (alt_vip_cti_0_dout_ready),                          //                  .ready
		.is_sop            (alt_vip_cti_0_dout_startofpacket),                  //                  .startofpacket
		.is_eop            (alt_vip_cti_0_dout_endofpacket),                    //                  .endofpacket
		.vid_clk           (vid_clk_to_the_alt_vip_cti_0),                      //     clocked_video.export
		.vid_data          (vid_data_to_the_alt_vip_cti_0),                     //                  .export
		.overflow          (overflow_from_the_alt_vip_cti_0),                   //                  .export
		.vid_datavalid     (vid_datavalid_to_the_alt_vip_cti_0),                //                  .export
		.vid_locked        (vid_locked_to_the_alt_vip_cti_0)                    //                  .export
	);

	DE1_SoC_QSYS_alt_vip_cpr_0 alt_vip_cpr_0 (
		.clock               (pll_sys_outclk0_clk),                // clock.clk
		.reset               (rst_controller_002_reset_out_reset), // reset.reset
		.din0_ready          (alt_vip_cti_0_dout_ready),           //  din0.ready
		.din0_valid          (alt_vip_cti_0_dout_valid),           //      .valid
		.din0_data           (alt_vip_cti_0_dout_data),            //      .data
		.din0_startofpacket  (alt_vip_cti_0_dout_startofpacket),   //      .startofpacket
		.din0_endofpacket    (alt_vip_cti_0_dout_endofpacket),     //      .endofpacket
		.dout0_ready         (alt_vip_cpr_0_dout0_ready),          // dout0.ready
		.dout0_valid         (alt_vip_cpr_0_dout0_valid),          //      .valid
		.dout0_data          (alt_vip_cpr_0_dout0_data),           //      .data
		.dout0_startofpacket (alt_vip_cpr_0_dout0_startofpacket),  //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_0_dout0_endofpacket)     //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_dil_0 alt_vip_dil_0 (
		.clock              (pll_sys_outclk0_clk),                // clock.clk
		.reset              (rst_controller_002_reset_out_reset), // reset.reset
		.din_ready          (alt_vip_cpr_0_dout0_ready),          //   din.ready
		.din_valid          (alt_vip_cpr_0_dout0_valid),          //      .valid
		.din_data           (alt_vip_cpr_0_dout0_data),           //      .data
		.din_startofpacket  (alt_vip_cpr_0_dout0_startofpacket),  //      .startofpacket
		.din_endofpacket    (alt_vip_cpr_0_dout0_endofpacket),    //      .endofpacket
		.dout_ready         (alt_vip_dil_0_dout_ready),           //  dout.ready
		.dout_valid         (alt_vip_dil_0_dout_valid),           //      .valid
		.dout_data          (alt_vip_dil_0_dout_data),            //      .data
		.dout_startofpacket (alt_vip_dil_0_dout_startofpacket),   //      .startofpacket
		.dout_endofpacket   (alt_vip_dil_0_dout_endofpacket)      //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_crs_0 alt_vip_crs_0 (
		.clock              (pll_sys_outclk0_clk),                // clock.clk
		.reset              (rst_controller_002_reset_out_reset), // reset.reset
		.din_ready          (alt_vip_dil_0_dout_ready),           //   din.ready
		.din_valid          (alt_vip_dil_0_dout_valid),           //      .valid
		.din_data           (alt_vip_dil_0_dout_data),            //      .data
		.din_startofpacket  (alt_vip_dil_0_dout_startofpacket),   //      .startofpacket
		.din_endofpacket    (alt_vip_dil_0_dout_endofpacket),     //      .endofpacket
		.dout_ready         (alt_vip_crs_0_dout_ready),           //  dout.ready
		.dout_valid         (alt_vip_crs_0_dout_valid),           //      .valid
		.dout_data          (alt_vip_crs_0_dout_data),            //      .data
		.dout_startofpacket (alt_vip_crs_0_dout_startofpacket),   //      .startofpacket
		.dout_endofpacket   (alt_vip_crs_0_dout_endofpacket)      //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_csc_0 alt_vip_csc_0 (
		.clock              (pll_sys_outclk0_clk),                // clock.clk
		.reset              (rst_controller_002_reset_out_reset), // reset.reset
		.din_ready          (alt_vip_crs_0_dout_ready),           //   din.ready
		.din_valid          (alt_vip_crs_0_dout_valid),           //      .valid
		.din_data           (alt_vip_crs_0_dout_data),            //      .data
		.din_startofpacket  (alt_vip_crs_0_dout_startofpacket),   //      .startofpacket
		.din_endofpacket    (alt_vip_crs_0_dout_endofpacket),     //      .endofpacket
		.dout_ready         (alt_vip_csc_0_dout_ready),           //  dout.ready
		.dout_valid         (alt_vip_csc_0_dout_valid),           //      .valid
		.dout_data          (alt_vip_csc_0_dout_data),            //      .data
		.dout_startofpacket (alt_vip_csc_0_dout_startofpacket),   //      .startofpacket
		.dout_endofpacket   (alt_vip_csc_0_dout_endofpacket)      //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_clip_0 alt_vip_clip_0 (
		.clock              (pll_sys_outclk0_clk),                // clock.clk
		.reset              (rst_controller_002_reset_out_reset), // reset.reset
		.din_ready          (alt_vip_csc_0_dout_ready),           //   din.ready
		.din_valid          (alt_vip_csc_0_dout_valid),           //      .valid
		.din_data           (alt_vip_csc_0_dout_data),            //      .data
		.din_startofpacket  (alt_vip_csc_0_dout_startofpacket),   //      .startofpacket
		.din_endofpacket    (alt_vip_csc_0_dout_endofpacket),     //      .endofpacket
		.dout_ready         (alt_vip_clip_0_dout_ready),          //  dout.ready
		.dout_valid         (alt_vip_clip_0_dout_valid),          //      .valid
		.dout_data          (alt_vip_clip_0_dout_data),           //      .data
		.dout_startofpacket (alt_vip_clip_0_dout_startofpacket),  //      .startofpacket
		.dout_endofpacket   (alt_vip_clip_0_dout_endofpacket)     //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_vfb_0 alt_vip_vfb_0 (
		.clock                        (pll_sys_outclk0_clk),                     //        clock.clk
		.reset                        (rst_controller_002_reset_out_reset),      //        reset.reset
		.din_ready                    (alt_vip_cl_scl_0_dout_ready),             //          din.ready
		.din_valid                    (alt_vip_cl_scl_0_dout_valid),             //             .valid
		.din_data                     (alt_vip_cl_scl_0_dout_data),              //             .data
		.din_startofpacket            (alt_vip_cl_scl_0_dout_startofpacket),     //             .startofpacket
		.din_endofpacket              (alt_vip_cl_scl_0_dout_endofpacket),       //             .endofpacket
		.dout_ready                   (alt_vip_vfb_0_dout_ready),                //         dout.ready
		.dout_valid                   (alt_vip_vfb_0_dout_valid),                //             .valid
		.dout_data                    (alt_vip_vfb_0_dout_data),                 //             .data
		.dout_startofpacket           (alt_vip_vfb_0_dout_startofpacket),        //             .startofpacket
		.dout_endofpacket             (alt_vip_vfb_0_dout_endofpacket),          //             .endofpacket
		.read_master_av_address       (alt_vip_vfb_0_read_master_address),       //  read_master.address
		.read_master_av_read          (alt_vip_vfb_0_read_master_read),          //             .read
		.read_master_av_waitrequest   (alt_vip_vfb_0_read_master_waitrequest),   //             .waitrequest
		.read_master_av_readdatavalid (alt_vip_vfb_0_read_master_readdatavalid), //             .readdatavalid
		.read_master_av_readdata      (alt_vip_vfb_0_read_master_readdata),      //             .readdata
		.read_master_av_burstcount    (alt_vip_vfb_0_read_master_burstcount),    //             .burstcount
		.write_master_av_address      (alt_vip_vfb_0_write_master_address),      // write_master.address
		.write_master_av_write        (alt_vip_vfb_0_write_master_write),        //             .write
		.write_master_av_writedata    (alt_vip_vfb_0_write_master_writedata),    //             .writedata
		.write_master_av_waitrequest  (alt_vip_vfb_0_write_master_waitrequest),  //             .waitrequest
		.write_master_av_burstcount   (alt_vip_vfb_0_write_master_burstcount)    //             .burstcount
	);

	DE1_SoC_QSYS_td_status td_status (
		.clk      (pll_sys_outclk2_clk),                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_2_td_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_2_td_status_s1_readdata), //                    .readdata
		.in_port  (in_port_to_the_td_status)                 // external_connection.export
	);

	DE1_SoC_QSYS_i2c_scl td_reset_n (
		.clk        (pll_sys_outclk2_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_2_td_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_td_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_td_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_td_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_td_reset_n_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_td_reset_n)                // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (256),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) clock_crossing_io_slow (
		.m0_clk           (pll_sys_outclk2_clk),                                       //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (pll_sys_outclk0_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                        // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_clock_crossing_io_slow_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_clock_crossing_io_slow_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_clock_crossing_io_slow_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_clock_crossing_io_slow_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_clock_crossing_io_slow_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_clock_crossing_io_slow_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_clock_crossing_io_slow_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_clock_crossing_io_slow_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_clock_crossing_io_slow_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_clock_crossing_io_slow_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_io_slow_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_io_slow_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_io_slow_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_io_slow_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_io_slow_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_io_slow_m0_address),                         //         .address
		.m0_write         (clock_crossing_io_slow_m0_write),                           //         .write
		.m0_read          (clock_crossing_io_slow_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_io_slow_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_io_slow_m0_debugaccess)                      //         .debugaccess
	);

	DE1_SoC_QSYS_cpu cpu (
		.clk                                   (pll_sys_outclk0_clk),                                 //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	DE1_SoC_QSYS_sysid sysid (
		.clock    (pll_sys_outclk2_clk),                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_control_slave_address)   //              .address
	);

	DE1_SoC_QSYS_alt_vip_cl_scl_0 #(
		.SYMBOLS_IN_SEQ      (1),
		.SYMBOLS_IN_PAR      (3),
		.BITS_PER_SYMBOL     (8),
		.EXTRA_PIPELINING    (0),
		.IS_422              (0),
		.NO_BLANKING         (1),
		.MAX_IN_WIDTH        (640),
		.MAX_IN_HEIGHT       (480),
		.MAX_OUT_WIDTH       (270),
		.MAX_OUT_HEIGHT      (200),
		.RUNTIME_CONTROL     (0),
		.ALWAYS_DOWNSCALE    (1),
		.ALGORITHM_NAME      ("POLYPHASE"),
		.DEFAULT_EDGE_THRESH (7),
		.DEFAULT_UPPER_BLUR  (15),
		.DEFAULT_LOWER_BLUR  (0),
		.ENABLE_FIR          (0),
		.ARE_IDENTICAL       (1),
		.V_TAPS              (8),
		.V_PHASES            (16),
		.H_TAPS              (8),
		.H_PHASES            (16),
		.V_SIGNED            (1),
		.V_INTEGER_BITS      (1),
		.V_FRACTION_BITS     (7),
		.H_SIGNED            (1),
		.H_INTEGER_BITS      (1),
		.H_FRACTION_BITS     (7),
		.PRESERVE_BITS       (0),
		.LOAD_AT_RUNTIME     (0),
		.V_BANKS             (1),
		.V_SYMMETRIC         (0),
		.V_FUNCTION          ("LANCZOS_2"),
		.V_COEFF_FILE        ("<enter file name (including full path)>"),
		.H_BANKS             (1),
		.H_SYMMETRIC         (0),
		.H_FUNCTION          ("LANCZOS_2"),
		.H_COEFF_FILE        ("<enter file name (including full path)>"),
		.IS_420              (0)
	) alt_vip_cl_scl_0 (
		.main_clock         (pll_sys_outclk0_clk),                 // main_clock.clk
		.main_reset         (rst_controller_002_reset_out_reset),  // main_reset.reset
		.din_data           (alt_vip_clip_0_dout_data),            //        din.data
		.din_valid          (alt_vip_clip_0_dout_valid),           //           .valid
		.din_startofpacket  (alt_vip_clip_0_dout_startofpacket),   //           .startofpacket
		.din_endofpacket    (alt_vip_clip_0_dout_endofpacket),     //           .endofpacket
		.din_ready          (alt_vip_clip_0_dout_ready),           //           .ready
		.dout_data          (alt_vip_cl_scl_0_dout_data),          //       dout.data
		.dout_valid         (alt_vip_cl_scl_0_dout_valid),         //           .valid
		.dout_startofpacket (alt_vip_cl_scl_0_dout_startofpacket), //           .startofpacket
		.dout_endofpacket   (alt_vip_cl_scl_0_dout_endofpacket),   //           .endofpacket
		.dout_ready         (alt_vip_cl_scl_0_dout_ready)          //           .ready
	);

	DE1_SoC_QSYS_pll_sys pll_sys (
		.refclk   (clk_50),                             //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (pll_sys_outclk0_clk),                // outclk0.clk
		.outclk_1 (clk_sdram_clk),                      // outclk1.clk
		.outclk_2 (pll_sys_outclk2_clk),                // outclk2.clk
		.outclk_3 (clk_vga_clk),                        // outclk3.clk
		.outclk_4 (pll_sys_outclk4_clk),                // outclk4.clk
		.locked   (pll_0_locked_export)                 //  locked.export
	);

	SEG7_IF #(
		.SEG7_NUM       (6),
		.ADDR_WIDTH     (3),
		.DEFAULT_ACTIVE (1),
		.LOW_ACTIVE     (1)
	) seg7 (
		.s_address   (mm_interconnect_0_seg7_avalon_slave_address),   //     avalon_slave.address
		.s_read      (mm_interconnect_0_seg7_avalon_slave_read),      //                 .read
		.s_readdata  (mm_interconnect_0_seg7_avalon_slave_readdata),  //                 .readdata
		.s_write     (mm_interconnect_0_seg7_avalon_slave_write),     //                 .write
		.s_writedata (mm_interconnect_0_seg7_avalon_slave_writedata), //                 .writedata
		.SEG7        (seg7_conduit_end_export),                       //      conduit_end.export
		.s_clk       (pll_sys_outclk2_clk),                           //       clock_sink.clk
		.s_reset     (rst_controller_reset_out_reset)                 // clock_sink_reset.reset
	);

	DE1_SoC_QSYS_sw sw (
		.clk        (pll_sys_outclk2_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        ()                                    //                 irq.irq
	);

	DE1_SoC_QSYS_key key (
		.clk        (pll_sys_outclk2_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        ()                                     //                 irq.irq
	);

	DE1_SoC_QSYS_ledr ledr (
		.clk        (pll_sys_outclk2_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)       // external_connection.export
	);

	DE1_SoC_QSYS_spi_0 spi_0 (
		.clk           (pll_sys_outclk4_clk),                                 //              clk.clk
		.reset_n       (~rst_controller_004_reset_out_reset),                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_3_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_3_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_3_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_3_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_3_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_3_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_001_receiver_irq),                   //              irq.irq
		.MISO          (spi_0_external_MISO),                                 //         external.export
		.MOSI          (spi_0_external_MOSI),                                 //                 .export
		.SCLK          (spi_0_external_SCLK),                                 //                 .export
		.SS_n          (spi_0_external_SS_n)                                  //                 .export
	);

	AUDIO_IF audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (pll_audio_outclk0_clk),                          //       clock_sink.clk
		.avs_s1_reset         (rst_controller_005_reset_out_reset),             // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	DE1_SoC_QSYS_pll_audio pll_audio (
		.refclk   (clk_50),                             //  refclk.clk
		.rst      (rst_controller_003_reset_out_reset), //   reset.reset
		.outclk_0 (pll_audio_outclk0_clk),              // outclk0.clk
		.locked   (pll_audio_locked_export)             //  locked.export
	);

	DE1_SoC_QSYS_uart uart (
		.clk           (pll_sys_outclk0_clk),                     //                 clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_external_connection_rxd),            // external_connection.export
		.txd           (uart_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	DE1_SoC_QSYS_timer_stamp timer_stamp (
		.clk        (pll_sys_outclk0_clk),                         //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_stamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_stamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_stamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_stamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_stamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                     //   irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) mm_clock_crossing_bridge_1 (
		.m0_clk           (pll_sys_outclk4_clk),                                           //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (pll_sys_outclk0_clk),                                           //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_1_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_1_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_1_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_1_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_1_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_1_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_1_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_1_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_1_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_1_m0_debugaccess)                      //         .debugaccess
	);

	DE1_SoC_QSYS_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                  //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),               //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                 //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                 //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                 //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                 //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                 //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                 //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                  //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),               //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),               //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),               //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                 //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                 //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                 //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                   //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                   //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                   //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                   //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                   //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                   //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                   //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                    //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                    //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                    //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                    //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                    //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                    //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                    //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                    //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                    //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                   //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                   //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                   //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                   //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                  //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                 //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                 //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                  //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                   //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                   //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                   //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                   //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                   //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_50),                                        //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                              //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                              //                  .awaddr
		.h2f_AWLEN                (),                                              //                  .awlen
		.h2f_AWSIZE               (),                                              //                  .awsize
		.h2f_AWBURST              (),                                              //                  .awburst
		.h2f_AWLOCK               (),                                              //                  .awlock
		.h2f_AWCACHE              (),                                              //                  .awcache
		.h2f_AWPROT               (),                                              //                  .awprot
		.h2f_AWVALID              (),                                              //                  .awvalid
		.h2f_AWREADY              (),                                              //                  .awready
		.h2f_WID                  (),                                              //                  .wid
		.h2f_WDATA                (),                                              //                  .wdata
		.h2f_WSTRB                (),                                              //                  .wstrb
		.h2f_WLAST                (),                                              //                  .wlast
		.h2f_WVALID               (),                                              //                  .wvalid
		.h2f_WREADY               (),                                              //                  .wready
		.h2f_BID                  (),                                              //                  .bid
		.h2f_BRESP                (),                                              //                  .bresp
		.h2f_BVALID               (),                                              //                  .bvalid
		.h2f_BREADY               (),                                              //                  .bready
		.h2f_ARID                 (),                                              //                  .arid
		.h2f_ARADDR               (),                                              //                  .araddr
		.h2f_ARLEN                (),                                              //                  .arlen
		.h2f_ARSIZE               (),                                              //                  .arsize
		.h2f_ARBURST              (),                                              //                  .arburst
		.h2f_ARLOCK               (),                                              //                  .arlock
		.h2f_ARCACHE              (),                                              //                  .arcache
		.h2f_ARPROT               (),                                              //                  .arprot
		.h2f_ARVALID              (),                                              //                  .arvalid
		.h2f_ARREADY              (),                                              //                  .arready
		.h2f_RID                  (),                                              //                  .rid
		.h2f_RDATA                (),                                              //                  .rdata
		.h2f_RRESP                (),                                              //                  .rresp
		.h2f_RLAST                (),                                              //                  .rlast
		.h2f_RVALID               (),                                              //                  .rvalid
		.h2f_RREADY               (),                                              //                  .rready
		.f2h_axi_clk              (clk_50),                                        //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_4_hps_0_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_4_hps_0_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_4_hps_0_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_4_hps_0_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_4_hps_0_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_4_hps_0_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_4_hps_0_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_4_hps_0_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_4_hps_0_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_4_hps_0_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_4_hps_0_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_4_hps_0_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_4_hps_0_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_4_hps_0_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_4_hps_0_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_4_hps_0_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_4_hps_0_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_4_hps_0_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_4_hps_0_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_4_hps_0_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_4_hps_0_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_4_hps_0_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_4_hps_0_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_4_hps_0_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_4_hps_0_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_4_hps_0_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_4_hps_0_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_4_hps_0_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_4_hps_0_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_4_hps_0_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_4_hps_0_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_4_hps_0_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_4_hps_0_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_4_hps_0_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_4_hps_0_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_4_hps_0_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_4_hps_0_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_4_hps_0_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (clk_50),                                        //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (1024),
		.MAX_IMAGE_HEIGHT               (768),
		.MEM_PORT_WIDTH                 (128),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_0 (
		.clock                (pll_sys_outclk0_clk),                                    //             clock_reset.clk
		.reset                (rst_controller_002_reset_out_reset),                     //       clock_reset_reset.reset
		.master_clock         (pll_sys_outclk0_clk),                                    //            clock_master.clk
		.master_reset         (rst_controller_002_reset_out_reset),                     //      clock_master_reset.reset
		.slave_address        (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1024),
		.V_ACTIVE_LINES                (768),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (10240),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (10239),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (24),
		.H_BACK_PORCH                  (160),
		.V_SYNC_LENGTH                 (6),
		.V_FRONT_PORCH                 (3),
		.V_BACK_PORCH                  (29),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_sys_outclk0_clk),                       //       is_clk_rst.clk
		.rst           (rst_controller_002_reset_out_reset),        // is_clk_rst_reset.reset
		.is_data       (alt_vip_mix_0_dout_data),                   //              din.data
		.is_valid      (alt_vip_mix_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_mix_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_mix_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_mix_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	DE1_SoC_QSYS_alt_vip_cpr_1 alt_vip_cpr_1 (
		.clock               (pll_sys_outclk0_clk),                                 // clock.clk
		.reset               (rst_controller_002_reset_out_reset),                  // reset.reset
		.din0_ready          (alt_vip_vfr_0_avalon_streaming_source_ready),         //  din0.ready
		.din0_valid          (alt_vip_vfr_0_avalon_streaming_source_valid),         //      .valid
		.din0_data           (alt_vip_vfr_0_avalon_streaming_source_data),          //      .data
		.din0_startofpacket  (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //      .startofpacket
		.din0_endofpacket    (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //      .endofpacket
		.dout0_ready         (alt_vip_cpr_1_dout0_ready),                           // dout0.ready
		.dout0_valid         (alt_vip_cpr_1_dout0_valid),                           //      .valid
		.dout0_data          (alt_vip_cpr_1_dout0_data),                            //      .data
		.dout0_startofpacket (alt_vip_cpr_1_dout0_startofpacket),                   //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_1_dout0_endofpacket)                      //      .endofpacket
	);

	DE1_SoC_QSYS_alt_vip_mix_0 alt_vip_mix_0 (
		.clock                 (pll_sys_outclk0_clk),                                //   clock.clk
		.reset                 (rst_controller_002_reset_out_reset),                 //   reset.reset
		.din_0_ready           (alt_vip_cpr_1_dout0_ready),                          //   din_0.ready
		.din_0_valid           (alt_vip_cpr_1_dout0_valid),                          //        .valid
		.din_0_data            (alt_vip_cpr_1_dout0_data),                           //        .data
		.din_0_startofpacket   (alt_vip_cpr_1_dout0_startofpacket),                  //        .startofpacket
		.din_0_endofpacket     (alt_vip_cpr_1_dout0_endofpacket),                    //        .endofpacket
		.din_1_ready           (alt_vip_cpr_2_dout0_ready),                          //   din_1.ready
		.din_1_valid           (alt_vip_cpr_2_dout0_valid),                          //        .valid
		.din_1_data            (alt_vip_cpr_2_dout0_data),                           //        .data
		.din_1_startofpacket   (alt_vip_cpr_2_dout0_startofpacket),                  //        .startofpacket
		.din_1_endofpacket     (alt_vip_cpr_2_dout0_endofpacket),                    //        .endofpacket
		.dout_ready            (alt_vip_mix_0_dout_ready),                           //    dout.ready
		.dout_valid            (alt_vip_mix_0_dout_valid),                           //        .valid
		.dout_data             (alt_vip_mix_0_dout_data),                            //        .data
		.dout_startofpacket    (alt_vip_mix_0_dout_startofpacket),                   //        .startofpacket
		.dout_endofpacket      (alt_vip_mix_0_dout_endofpacket),                     //        .endofpacket
		.control_av_chipselect (mm_interconnect_0_alt_vip_mix_0_control_chipselect), // control.chipselect
		.control_av_write      (mm_interconnect_0_alt_vip_mix_0_control_write),      //        .write
		.control_av_address    (mm_interconnect_0_alt_vip_mix_0_control_address),    //        .address
		.control_av_writedata  (mm_interconnect_0_alt_vip_mix_0_control_writedata),  //        .writedata
		.control_av_readdata   (mm_interconnect_0_alt_vip_mix_0_control_readdata)    //        .readdata
	);

	DE1_SoC_QSYS_alt_vip_cpr_2 alt_vip_cpr_2 (
		.clock               (pll_sys_outclk0_clk),                // clock.clk
		.reset               (rst_controller_002_reset_out_reset), // reset.reset
		.din0_ready          (alt_vip_vfb_0_dout_ready),           //  din0.ready
		.din0_valid          (alt_vip_vfb_0_dout_valid),           //      .valid
		.din0_data           (alt_vip_vfb_0_dout_data),            //      .data
		.din0_startofpacket  (alt_vip_vfb_0_dout_startofpacket),   //      .startofpacket
		.din0_endofpacket    (alt_vip_vfb_0_dout_endofpacket),     //      .endofpacket
		.dout0_ready         (alt_vip_cpr_2_dout0_ready),          // dout0.ready
		.dout0_valid         (alt_vip_cpr_2_dout0_valid),          //      .valid
		.dout0_data          (alt_vip_cpr_2_dout0_data),           //      .data
		.dout0_startofpacket (alt_vip_cpr_2_dout0_startofpacket),  //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_2_dout0_endofpacket)     //      .endofpacket
	);

	TERASIC_IR_RX_FIFO ir_rx (
		.s_read      (mm_interconnect_0_ir_rx_avalon_slave_read),        //     avalon_slave.read
		.s_cs_n      (~mm_interconnect_0_ir_rx_avalon_slave_chipselect), //                 .chipselect_n
		.s_readdata  (mm_interconnect_0_ir_rx_avalon_slave_readdata),    //                 .readdata
		.s_write     (mm_interconnect_0_ir_rx_avalon_slave_write),       //                 .write
		.s_writedata (mm_interconnect_0_ir_rx_avalon_slave_writedata),   //                 .writedata
		.s_address   (mm_interconnect_0_ir_rx_avalon_slave_address),     //                 .address
		.clk         (clk_50),                                           //       clock_sink.clk
		.reset_n     (~rst_controller_003_reset_out_reset),              // clock_sink_reset.reset_n
		.ir          (ir_rx_conduit_end_export),                         //      conduit_end.export
		.irq         ()                                                  // interrupt_sender.irq
	);

	DE1_SoC_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                  //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                 //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                               //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                               //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                               //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                               //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                   //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                 //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                 //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                 //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                   //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                 //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                  //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                 //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                               //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                               //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                               //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                               //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                   //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                 //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                 //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                 //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                //                                                              .rready
		.clk_50_clk_clk                                                      (clk_50),                                                        //                                                    clk_50_clk.clk
		.pll_audio_outclk0_clk                                               (pll_audio_outclk0_clk),                                         //                                             pll_audio_outclk0.clk
		.pll_sys_outclk0_clk                                                 (pll_sys_outclk0_clk),                                           //                                               pll_sys_outclk0.clk
		.pll_sys_outclk2_clk                                                 (pll_sys_outclk2_clk),                                           //                                               pll_sys_outclk2.clk
		.audio_clock_sink_reset_reset_bridge_in_reset_reset                  (rst_controller_005_reset_out_reset),                            //                  audio_clock_sink_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                             (rst_controller_002_reset_out_reset),                            //                             cpu_reset_n_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                            // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.ir_rx_clock_sink_reset_reset_bridge_in_reset_reset                  (rst_controller_003_reset_out_reset),                            //                  ir_rx_clock_sink_reset_reset_bridge_in_reset.reset
		.ledr_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                                //                              ledr_reset_reset_bridge_in_reset.reset
		.onchip_memory2_reset1_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                            //                   onchip_memory2_reset1_reset_bridge_in_reset.reset
		.cpu_data_master_address                                             (cpu_data_master_address),                                       //                                               cpu_data_master.address
		.cpu_data_master_waitrequest                                         (cpu_data_master_waitrequest),                                   //                                                              .waitrequest
		.cpu_data_master_byteenable                                          (cpu_data_master_byteenable),                                    //                                                              .byteenable
		.cpu_data_master_read                                                (cpu_data_master_read),                                          //                                                              .read
		.cpu_data_master_readdata                                            (cpu_data_master_readdata),                                      //                                                              .readdata
		.cpu_data_master_readdatavalid                                       (cpu_data_master_readdatavalid),                                 //                                                              .readdatavalid
		.cpu_data_master_write                                               (cpu_data_master_write),                                         //                                                              .write
		.cpu_data_master_writedata                                           (cpu_data_master_writedata),                                     //                                                              .writedata
		.cpu_data_master_debugaccess                                         (cpu_data_master_debugaccess),                                   //                                                              .debugaccess
		.cpu_instruction_master_address                                      (cpu_instruction_master_address),                                //                                        cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                                  (cpu_instruction_master_waitrequest),                            //                                                              .waitrequest
		.cpu_instruction_master_read                                         (cpu_instruction_master_read),                                   //                                                              .read
		.cpu_instruction_master_readdata                                     (cpu_instruction_master_readdata),                               //                                                              .readdata
		.cpu_instruction_master_readdatavalid                                (cpu_instruction_master_readdatavalid),                          //                                                              .readdatavalid
		.alt_vip_cti_0_control_address                                       (mm_interconnect_0_alt_vip_cti_0_control_address),               //                                         alt_vip_cti_0_control.address
		.alt_vip_cti_0_control_write                                         (mm_interconnect_0_alt_vip_cti_0_control_write),                 //                                                              .write
		.alt_vip_cti_0_control_read                                          (mm_interconnect_0_alt_vip_cti_0_control_read),                  //                                                              .read
		.alt_vip_cti_0_control_readdata                                      (mm_interconnect_0_alt_vip_cti_0_control_readdata),              //                                                              .readdata
		.alt_vip_cti_0_control_writedata                                     (mm_interconnect_0_alt_vip_cti_0_control_writedata),             //                                                              .writedata
		.alt_vip_mix_0_control_address                                       (mm_interconnect_0_alt_vip_mix_0_control_address),               //                                         alt_vip_mix_0_control.address
		.alt_vip_mix_0_control_write                                         (mm_interconnect_0_alt_vip_mix_0_control_write),                 //                                                              .write
		.alt_vip_mix_0_control_readdata                                      (mm_interconnect_0_alt_vip_mix_0_control_readdata),              //                                                              .readdata
		.alt_vip_mix_0_control_writedata                                     (mm_interconnect_0_alt_vip_mix_0_control_writedata),             //                                                              .writedata
		.alt_vip_mix_0_control_chipselect                                    (mm_interconnect_0_alt_vip_mix_0_control_chipselect),            //                                                              .chipselect
		.alt_vip_vfr_0_avalon_slave_address                                  (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),          //                                    alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                                    (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),            //                                                              .write
		.alt_vip_vfr_0_avalon_slave_read                                     (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),             //                                                              .read
		.alt_vip_vfr_0_avalon_slave_readdata                                 (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),         //                                                              .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                                (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata),        //                                                              .writedata
		.audio_avalon_slave_address                                          (mm_interconnect_0_audio_avalon_slave_address),                  //                                            audio_avalon_slave.address
		.audio_avalon_slave_write                                            (mm_interconnect_0_audio_avalon_slave_write),                    //                                                              .write
		.audio_avalon_slave_read                                             (mm_interconnect_0_audio_avalon_slave_read),                     //                                                              .read
		.audio_avalon_slave_readdata                                         (mm_interconnect_0_audio_avalon_slave_readdata),                 //                                                              .readdata
		.audio_avalon_slave_writedata                                        (mm_interconnect_0_audio_avalon_slave_writedata),                //                                                              .writedata
		.clock_crossing_io_slow_s0_address                                   (mm_interconnect_0_clock_crossing_io_slow_s0_address),           //                                     clock_crossing_io_slow_s0.address
		.clock_crossing_io_slow_s0_write                                     (mm_interconnect_0_clock_crossing_io_slow_s0_write),             //                                                              .write
		.clock_crossing_io_slow_s0_read                                      (mm_interconnect_0_clock_crossing_io_slow_s0_read),              //                                                              .read
		.clock_crossing_io_slow_s0_readdata                                  (mm_interconnect_0_clock_crossing_io_slow_s0_readdata),          //                                                              .readdata
		.clock_crossing_io_slow_s0_writedata                                 (mm_interconnect_0_clock_crossing_io_slow_s0_writedata),         //                                                              .writedata
		.clock_crossing_io_slow_s0_burstcount                                (mm_interconnect_0_clock_crossing_io_slow_s0_burstcount),        //                                                              .burstcount
		.clock_crossing_io_slow_s0_byteenable                                (mm_interconnect_0_clock_crossing_io_slow_s0_byteenable),        //                                                              .byteenable
		.clock_crossing_io_slow_s0_readdatavalid                             (mm_interconnect_0_clock_crossing_io_slow_s0_readdatavalid),     //                                                              .readdatavalid
		.clock_crossing_io_slow_s0_waitrequest                               (mm_interconnect_0_clock_crossing_io_slow_s0_waitrequest),       //                                                              .waitrequest
		.clock_crossing_io_slow_s0_debugaccess                               (mm_interconnect_0_clock_crossing_io_slow_s0_debugaccess),       //                                                              .debugaccess
		.cpu_jtag_debug_module_address                                       (mm_interconnect_0_cpu_jtag_debug_module_address),               //                                         cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                         (mm_interconnect_0_cpu_jtag_debug_module_write),                 //                                                              .write
		.cpu_jtag_debug_module_read                                          (mm_interconnect_0_cpu_jtag_debug_module_read),                  //                                                              .read
		.cpu_jtag_debug_module_readdata                                      (mm_interconnect_0_cpu_jtag_debug_module_readdata),              //                                                              .readdata
		.cpu_jtag_debug_module_writedata                                     (mm_interconnect_0_cpu_jtag_debug_module_writedata),             //                                                              .writedata
		.cpu_jtag_debug_module_byteenable                                    (mm_interconnect_0_cpu_jtag_debug_module_byteenable),            //                                                              .byteenable
		.cpu_jtag_debug_module_waitrequest                                   (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),           //                                                              .waitrequest
		.cpu_jtag_debug_module_debugaccess                                   (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),           //                                                              .debugaccess
		.ir_rx_avalon_slave_address                                          (mm_interconnect_0_ir_rx_avalon_slave_address),                  //                                            ir_rx_avalon_slave.address
		.ir_rx_avalon_slave_write                                            (mm_interconnect_0_ir_rx_avalon_slave_write),                    //                                                              .write
		.ir_rx_avalon_slave_read                                             (mm_interconnect_0_ir_rx_avalon_slave_read),                     //                                                              .read
		.ir_rx_avalon_slave_readdata                                         (mm_interconnect_0_ir_rx_avalon_slave_readdata),                 //                                                              .readdata
		.ir_rx_avalon_slave_writedata                                        (mm_interconnect_0_ir_rx_avalon_slave_writedata),                //                                                              .writedata
		.ir_rx_avalon_slave_chipselect                                       (mm_interconnect_0_ir_rx_avalon_slave_chipselect),               //                                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                                              .write
		.jtag_uart_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                                              .chipselect
		.key_s1_address                                                      (mm_interconnect_0_key_s1_address),                              //                                                        key_s1.address
		.key_s1_write                                                        (mm_interconnect_0_key_s1_write),                                //                                                              .write
		.key_s1_readdata                                                     (mm_interconnect_0_key_s1_readdata),                             //                                                              .readdata
		.key_s1_writedata                                                    (mm_interconnect_0_key_s1_writedata),                            //                                                              .writedata
		.key_s1_chipselect                                                   (mm_interconnect_0_key_s1_chipselect),                           //                                                              .chipselect
		.ledr_s1_address                                                     (mm_interconnect_0_ledr_s1_address),                             //                                                       ledr_s1.address
		.ledr_s1_write                                                       (mm_interconnect_0_ledr_s1_write),                               //                                                              .write
		.ledr_s1_readdata                                                    (mm_interconnect_0_ledr_s1_readdata),                            //                                                              .readdata
		.ledr_s1_writedata                                                   (mm_interconnect_0_ledr_s1_writedata),                           //                                                              .writedata
		.ledr_s1_chipselect                                                  (mm_interconnect_0_ledr_s1_chipselect),                          //                                                              .chipselect
		.mm_clock_crossing_bridge_1_s0_address                               (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_address),       //                                 mm_clock_crossing_bridge_1_s0.address
		.mm_clock_crossing_bridge_1_s0_write                                 (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_write),         //                                                              .write
		.mm_clock_crossing_bridge_1_s0_read                                  (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_read),          //                                                              .read
		.mm_clock_crossing_bridge_1_s0_readdata                              (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdata),      //                                                              .readdata
		.mm_clock_crossing_bridge_1_s0_writedata                             (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_writedata),     //                                                              .writedata
		.mm_clock_crossing_bridge_1_s0_burstcount                            (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_burstcount),    //                                                              .burstcount
		.mm_clock_crossing_bridge_1_s0_byteenable                            (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_byteenable),    //                                                              .byteenable
		.mm_clock_crossing_bridge_1_s0_readdatavalid                         (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_readdatavalid), //                                                              .readdatavalid
		.mm_clock_crossing_bridge_1_s0_waitrequest                           (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_waitrequest),   //                                                              .waitrequest
		.mm_clock_crossing_bridge_1_s0_debugaccess                           (mm_interconnect_0_mm_clock_crossing_bridge_1_s0_debugaccess),   //                                                              .debugaccess
		.onchip_memory2_s1_address                                           (mm_interconnect_0_onchip_memory2_s1_address),                   //                                             onchip_memory2_s1.address
		.onchip_memory2_s1_write                                             (mm_interconnect_0_onchip_memory2_s1_write),                     //                                                              .write
		.onchip_memory2_s1_readdata                                          (mm_interconnect_0_onchip_memory2_s1_readdata),                  //                                                              .readdata
		.onchip_memory2_s1_writedata                                         (mm_interconnect_0_onchip_memory2_s1_writedata),                 //                                                              .writedata
		.onchip_memory2_s1_byteenable                                        (mm_interconnect_0_onchip_memory2_s1_byteenable),                //                                                              .byteenable
		.onchip_memory2_s1_chipselect                                        (mm_interconnect_0_onchip_memory2_s1_chipselect),                //                                                              .chipselect
		.onchip_memory2_s1_clken                                             (mm_interconnect_0_onchip_memory2_s1_clken),                     //                                                              .clken
		.seg7_avalon_slave_address                                           (mm_interconnect_0_seg7_avalon_slave_address),                   //                                             seg7_avalon_slave.address
		.seg7_avalon_slave_write                                             (mm_interconnect_0_seg7_avalon_slave_write),                     //                                                              .write
		.seg7_avalon_slave_read                                              (mm_interconnect_0_seg7_avalon_slave_read),                      //                                                              .read
		.seg7_avalon_slave_readdata                                          (mm_interconnect_0_seg7_avalon_slave_readdata),                  //                                                              .readdata
		.seg7_avalon_slave_writedata                                         (mm_interconnect_0_seg7_avalon_slave_writedata),                 //                                                              .writedata
		.sw_s1_address                                                       (mm_interconnect_0_sw_s1_address),                               //                                                         sw_s1.address
		.sw_s1_write                                                         (mm_interconnect_0_sw_s1_write),                                 //                                                              .write
		.sw_s1_readdata                                                      (mm_interconnect_0_sw_s1_readdata),                              //                                                              .readdata
		.sw_s1_writedata                                                     (mm_interconnect_0_sw_s1_writedata),                             //                                                              .writedata
		.sw_s1_chipselect                                                    (mm_interconnect_0_sw_s1_chipselect),                            //                                                              .chipselect
		.timer_stamp_s1_address                                              (mm_interconnect_0_timer_stamp_s1_address),                      //                                                timer_stamp_s1.address
		.timer_stamp_s1_write                                                (mm_interconnect_0_timer_stamp_s1_write),                        //                                                              .write
		.timer_stamp_s1_readdata                                             (mm_interconnect_0_timer_stamp_s1_readdata),                     //                                                              .readdata
		.timer_stamp_s1_writedata                                            (mm_interconnect_0_timer_stamp_s1_writedata),                    //                                                              .writedata
		.timer_stamp_s1_chipselect                                           (mm_interconnect_0_timer_stamp_s1_chipselect),                   //                                                              .chipselect
		.uart_s1_address                                                     (mm_interconnect_0_uart_s1_address),                             //                                                       uart_s1.address
		.uart_s1_write                                                       (mm_interconnect_0_uart_s1_write),                               //                                                              .write
		.uart_s1_read                                                        (mm_interconnect_0_uart_s1_read),                                //                                                              .read
		.uart_s1_readdata                                                    (mm_interconnect_0_uart_s1_readdata),                            //                                                              .readdata
		.uart_s1_writedata                                                   (mm_interconnect_0_uart_s1_writedata),                           //                                                              .writedata
		.uart_s1_begintransfer                                               (mm_interconnect_0_uart_s1_begintransfer),                       //                                                              .begintransfer
		.uart_s1_chipselect                                                  (mm_interconnect_0_uart_s1_chipselect)                           //                                                              .chipselect
	);

	DE1_SoC_QSYS_mm_interconnect_1 mm_interconnect_1 (
		.pll_sys_outclk0_clk                             (pll_sys_outclk0_clk),                      //                           pll_sys_outclk0.clk
		.alt_vip_vfb_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),       // alt_vip_vfb_0_reset_reset_bridge_in_reset.reset
		.alt_vip_vfb_0_read_master_address               (alt_vip_vfb_0_read_master_address),        //                 alt_vip_vfb_0_read_master.address
		.alt_vip_vfb_0_read_master_waitrequest           (alt_vip_vfb_0_read_master_waitrequest),    //                                          .waitrequest
		.alt_vip_vfb_0_read_master_burstcount            (alt_vip_vfb_0_read_master_burstcount),     //                                          .burstcount
		.alt_vip_vfb_0_read_master_read                  (alt_vip_vfb_0_read_master_read),           //                                          .read
		.alt_vip_vfb_0_read_master_readdata              (alt_vip_vfb_0_read_master_readdata),       //                                          .readdata
		.alt_vip_vfb_0_read_master_readdatavalid         (alt_vip_vfb_0_read_master_readdatavalid),  //                                          .readdatavalid
		.alt_vip_vfb_0_write_master_address              (alt_vip_vfb_0_write_master_address),       //                alt_vip_vfb_0_write_master.address
		.alt_vip_vfb_0_write_master_waitrequest          (alt_vip_vfb_0_write_master_waitrequest),   //                                          .waitrequest
		.alt_vip_vfb_0_write_master_burstcount           (alt_vip_vfb_0_write_master_burstcount),    //                                          .burstcount
		.alt_vip_vfb_0_write_master_write                (alt_vip_vfb_0_write_master_write),         //                                          .write
		.alt_vip_vfb_0_write_master_writedata            (alt_vip_vfb_0_write_master_writedata),     //                                          .writedata
		.sdram_s1_address                                (mm_interconnect_1_sdram_s1_address),       //                                  sdram_s1.address
		.sdram_s1_write                                  (mm_interconnect_1_sdram_s1_write),         //                                          .write
		.sdram_s1_read                                   (mm_interconnect_1_sdram_s1_read),          //                                          .read
		.sdram_s1_readdata                               (mm_interconnect_1_sdram_s1_readdata),      //                                          .readdata
		.sdram_s1_writedata                              (mm_interconnect_1_sdram_s1_writedata),     //                                          .writedata
		.sdram_s1_byteenable                             (mm_interconnect_1_sdram_s1_byteenable),    //                                          .byteenable
		.sdram_s1_readdatavalid                          (mm_interconnect_1_sdram_s1_readdatavalid), //                                          .readdatavalid
		.sdram_s1_waitrequest                            (mm_interconnect_1_sdram_s1_waitrequest),   //                                          .waitrequest
		.sdram_s1_chipselect                             (mm_interconnect_1_sdram_s1_chipselect)     //                                          .chipselect
	);

	DE1_SoC_QSYS_mm_interconnect_2 mm_interconnect_2 (
		.pll_sys_outclk2_clk                                         (pll_sys_outclk2_clk),                            //                                       pll_sys_outclk2.clk
		.clock_crossing_io_slow_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // clock_crossing_io_slow_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_io_slow_m0_address                           (clock_crossing_io_slow_m0_address),              //                             clock_crossing_io_slow_m0.address
		.clock_crossing_io_slow_m0_waitrequest                       (clock_crossing_io_slow_m0_waitrequest),          //                                                      .waitrequest
		.clock_crossing_io_slow_m0_burstcount                        (clock_crossing_io_slow_m0_burstcount),           //                                                      .burstcount
		.clock_crossing_io_slow_m0_byteenable                        (clock_crossing_io_slow_m0_byteenable),           //                                                      .byteenable
		.clock_crossing_io_slow_m0_read                              (clock_crossing_io_slow_m0_read),                 //                                                      .read
		.clock_crossing_io_slow_m0_readdata                          (clock_crossing_io_slow_m0_readdata),             //                                                      .readdata
		.clock_crossing_io_slow_m0_readdatavalid                     (clock_crossing_io_slow_m0_readdatavalid),        //                                                      .readdatavalid
		.clock_crossing_io_slow_m0_write                             (clock_crossing_io_slow_m0_write),                //                                                      .write
		.clock_crossing_io_slow_m0_writedata                         (clock_crossing_io_slow_m0_writedata),            //                                                      .writedata
		.clock_crossing_io_slow_m0_debugaccess                       (clock_crossing_io_slow_m0_debugaccess),          //                                                      .debugaccess
		.i2c_scl_s1_address                                          (mm_interconnect_2_i2c_scl_s1_address),           //                                            i2c_scl_s1.address
		.i2c_scl_s1_write                                            (mm_interconnect_2_i2c_scl_s1_write),             //                                                      .write
		.i2c_scl_s1_readdata                                         (mm_interconnect_2_i2c_scl_s1_readdata),          //                                                      .readdata
		.i2c_scl_s1_writedata                                        (mm_interconnect_2_i2c_scl_s1_writedata),         //                                                      .writedata
		.i2c_scl_s1_chipselect                                       (mm_interconnect_2_i2c_scl_s1_chipselect),        //                                                      .chipselect
		.i2c_sda_s1_address                                          (mm_interconnect_2_i2c_sda_s1_address),           //                                            i2c_sda_s1.address
		.i2c_sda_s1_write                                            (mm_interconnect_2_i2c_sda_s1_write),             //                                                      .write
		.i2c_sda_s1_readdata                                         (mm_interconnect_2_i2c_sda_s1_readdata),          //                                                      .readdata
		.i2c_sda_s1_writedata                                        (mm_interconnect_2_i2c_sda_s1_writedata),         //                                                      .writedata
		.i2c_sda_s1_chipselect                                       (mm_interconnect_2_i2c_sda_s1_chipselect),        //                                                      .chipselect
		.sysid_control_slave_address                                 (mm_interconnect_2_sysid_control_slave_address),  //                                   sysid_control_slave.address
		.sysid_control_slave_readdata                                (mm_interconnect_2_sysid_control_slave_readdata), //                                                      .readdata
		.td_reset_n_s1_address                                       (mm_interconnect_2_td_reset_n_s1_address),        //                                         td_reset_n_s1.address
		.td_reset_n_s1_write                                         (mm_interconnect_2_td_reset_n_s1_write),          //                                                      .write
		.td_reset_n_s1_readdata                                      (mm_interconnect_2_td_reset_n_s1_readdata),       //                                                      .readdata
		.td_reset_n_s1_writedata                                     (mm_interconnect_2_td_reset_n_s1_writedata),      //                                                      .writedata
		.td_reset_n_s1_chipselect                                    (mm_interconnect_2_td_reset_n_s1_chipselect),     //                                                      .chipselect
		.td_status_s1_address                                        (mm_interconnect_2_td_status_s1_address),         //                                          td_status_s1.address
		.td_status_s1_readdata                                       (mm_interconnect_2_td_status_s1_readdata),        //                                                      .readdata
		.timer_s1_address                                            (mm_interconnect_2_timer_s1_address),             //                                              timer_s1.address
		.timer_s1_write                                              (mm_interconnect_2_timer_s1_write),               //                                                      .write
		.timer_s1_readdata                                           (mm_interconnect_2_timer_s1_readdata),            //                                                      .readdata
		.timer_s1_writedata                                          (mm_interconnect_2_timer_s1_writedata),           //                                                      .writedata
		.timer_s1_chipselect                                         (mm_interconnect_2_timer_s1_chipselect)           //                                                      .chipselect
	);

	DE1_SoC_QSYS_mm_interconnect_3 mm_interconnect_3 (
		.pll_sys_outclk4_clk                                             (pll_sys_outclk4_clk),                                 //                                           pll_sys_outclk4.clk
		.mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                  // mm_clock_crossing_bridge_1_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_1_m0_address                           (mm_clock_crossing_bridge_1_m0_address),               //                             mm_clock_crossing_bridge_1_m0.address
		.mm_clock_crossing_bridge_1_m0_waitrequest                       (mm_clock_crossing_bridge_1_m0_waitrequest),           //                                                          .waitrequest
		.mm_clock_crossing_bridge_1_m0_burstcount                        (mm_clock_crossing_bridge_1_m0_burstcount),            //                                                          .burstcount
		.mm_clock_crossing_bridge_1_m0_byteenable                        (mm_clock_crossing_bridge_1_m0_byteenable),            //                                                          .byteenable
		.mm_clock_crossing_bridge_1_m0_read                              (mm_clock_crossing_bridge_1_m0_read),                  //                                                          .read
		.mm_clock_crossing_bridge_1_m0_readdata                          (mm_clock_crossing_bridge_1_m0_readdata),              //                                                          .readdata
		.mm_clock_crossing_bridge_1_m0_readdatavalid                     (mm_clock_crossing_bridge_1_m0_readdatavalid),         //                                                          .readdatavalid
		.mm_clock_crossing_bridge_1_m0_write                             (mm_clock_crossing_bridge_1_m0_write),                 //                                                          .write
		.mm_clock_crossing_bridge_1_m0_writedata                         (mm_clock_crossing_bridge_1_m0_writedata),             //                                                          .writedata
		.mm_clock_crossing_bridge_1_m0_debugaccess                       (mm_clock_crossing_bridge_1_m0_debugaccess),           //                                                          .debugaccess
		.spi_0_spi_control_port_address                                  (mm_interconnect_3_spi_0_spi_control_port_address),    //                                    spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                                    (mm_interconnect_3_spi_0_spi_control_port_write),      //                                                          .write
		.spi_0_spi_control_port_read                                     (mm_interconnect_3_spi_0_spi_control_port_read),       //                                                          .read
		.spi_0_spi_control_port_readdata                                 (mm_interconnect_3_spi_0_spi_control_port_readdata),   //                                                          .readdata
		.spi_0_spi_control_port_writedata                                (mm_interconnect_3_spi_0_spi_control_port_writedata),  //                                                          .writedata
		.spi_0_spi_control_port_chipselect                               (mm_interconnect_3_spi_0_spi_control_port_chipselect)  //                                                          .chipselect
	);

	DE1_SoC_QSYS_mm_interconnect_4 mm_interconnect_4 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_4_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_4_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_4_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_4_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_4_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_4_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_4_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_4_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_4_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_4_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_4_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_4_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_4_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_4_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_4_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_4_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_50_clk_clk                                                   (clk_50),                                        //                                                 clk_50_clk.clk
		.pll_sys_outclk0_clk                                              (pll_sys_outclk0_clk),                           //                                            pll_sys_outclk0.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset     (rst_controller_002_reset_out_reset),            //     alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                              (alt_vip_vfr_0_avalon_master_address),           //                                alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                          (alt_vip_vfr_0_avalon_master_waitrequest),       //                                                           .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                           (alt_vip_vfr_0_avalon_master_burstcount),        //                                                           .burstcount
		.alt_vip_vfr_0_avalon_master_read                                 (alt_vip_vfr_0_avalon_master_read),              //                                                           .read
		.alt_vip_vfr_0_avalon_master_readdata                             (alt_vip_vfr_0_avalon_master_readdata),          //                                                           .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                        (alt_vip_vfr_0_avalon_master_readdatavalid)      //                                                           .readdatavalid
	);

	DE1_SoC_QSYS_irq_mapper irq_mapper (
		.clk           (pll_sys_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	DE1_SoC_QSYS_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	DE1_SoC_QSYS_irq_mapper_001 irq_mapper_002 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_sys_outclk2_clk),                //       receiver_clk.clk
		.sender_clk     (pll_sys_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_sys_outclk4_clk),                //       receiver_clk.clk
		.sender_clk     (pll_sys_outclk0_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_004_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                       // reset_in0.reset
		.clk            (pll_sys_outclk2_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (pll_sys_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.clk            (pll_sys_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (pll_sys_outclk4_clk),                //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (pll_audio_outclk0_clk),              //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_50),                             //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
