��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?[_�V�$�]ц�%��\S���f�[tֆ:[p�f���]p8	e�<_j� �|��GQ髞镵�vIl^l��Ք<�c��l2��)�U�����\�$�2�]���1s�VQ�!z�����J\۾��ǆ)��;�߾CH���a`'���2ށx����	���0�x�(���) �@e�z����J���J �=�^}f8����"
4�1{qYb|��K>ci�����_л���*��D̮��������Ic+�h�IS#!��]�m�4jYn���|o=�N+����D�:�n�[v�8@�������L�,nQͳig�2/�#��T�M��3�4J���oM�m�ѣ��ڱ�P����?�!N��l�N��Ak��4�X�Ǯ���c�4�9����SN��"�|M}�0ϓp0�[T��jP���H�S`|�o��4D����)vM��� ��;�+��n��I�֗��^�㷍����
����뙌�G_�iE���}�#y7o�q @��1
��c�k[�>8��D�'I��
|i<��Μx� ���;�8�r�����p!�Z�.������ X5^bP�o#;s�,�Pu:��װ��I���=��Vd}<���Ip�B��ޫ�p߯�j(��ǃ+nX���*�rx���7j�YI
�^*�#g3�o%�x����Kjk���͉s�\��c�5���ǟ;1`2�[[FY�ʓK�|�9�Y�[$0I�S(]@	֒�Ӗ��O����,�Y�ؐS0�򈕃 �&Bl7�Jѝ���rQ�<_K��0S�����~-'E?k�Z-�e�'�q'&��aNܝ]�,f�i�_Z���l�E��τ��xѨ�5����v��f~��B�i�1���9\��[w�(�b4|�r��j��� l�-��1ϕ�1�o��%p`�.mp�\�S2?[D[�L�;T�}�d�^Z�������1�F�R�D�}��>%�%!�2Yv������xA��]s�dQ���5�Q�I���r1x����-r�T�W|aZ�I0�G K^�U����~������Mѕ���!T�"���J�9�����'�Y�Re˺�iEpJ��s�J�4`O��Wr��z��ރ~Go�E�u�e=;":�(��S6�h�M�Ϯ��q�Y)x���m��N8�c��f�ֶ��.�֧��=E(t�S٧R���rr{��I�>�m}ͪk�M`"*g
�#�i�*no#L~��0E�w�_�p�@[Z�I��ˮ��|h %�AĢ������Ez��f-�+�mT1�(ճb<ťy0+@�E��)�	
t���f�4e��MlZ5�/L�Dpq�4j<��=��w��+��׾��$/Ӗ̒\A��>�j������Nc@���:�KљE��c���i����J��#&�+����s6iՌ:��0\^���=�6���A�I�V��S\���b��%�%ӊl��C�:F�E��G<��Aa|����_��p�Fi���K�v���3�ٜN�}��=���/�n�/��qO��9gK�sAk�g#�z92M���v��|���td�;����0�KQ�i>1K;%8�Ծ�Y .���Pz�d?�7D����t��/hC�����dW�d���5�-	*Hr�5/�6$ފJt���a5�d�>CfE�x���$Y4W{M�%�ʡ60���Q��-}l q��N�����uC�sp���:�g|lMgqr�J��\��ڙ����?b���
��+4퓖��i[��O�H-J&�x�����gf��X��̟W��$g����������|wvn��g���y���b_�[J��_I���VA����mW��IaE#�\�6�,��e�s���!�j�����o��]���n-�������!�-w<���Z�yP�qI�&'�9AA�V>��x�U�` 	'��+���Z�^ۥ^P�fd8��X��!�E3y��m�~�N�kM�H��f5wlq�Eq������W\ �c����Kq�I��с�OVmo?ݞ ��l���V�lB������1�)X�w+�������!�ʸ:�OX���'6�����5�w��W[d��p9�1�7p��M�a6��m�h�M�����}��� (De֧��EH&�켵F?�p�J�bt	w�jq�����o�]��O;�%0��'Ȯ��#��=RH[C���r�Nvo��y���I��d��,�,_<R�7�)��C��A),�%ػ��BM��4��q↹v�ʛ�;D� ��a�	7nGH�,��v{��n��cƚ�<=�$����m�A�{}c4��������pCż-�p#���N::����-��<^���,����ؠ��7�A�!�E'e�g�f�8�tU����������'Z���>D� {��`��`A*��wz��v�+��y�ω&x*Ґ�8�'n8�,���U�4H/�j�Y��ל����@��w�.yI3٠��Ka�?�Hg��9ތ�c��o�%_q��Đ1(	�����w�8fr��,g�'3���g�ك:���x�="j��8�BhO/�����hB����/��H�}�a�՟yp��0��Aǈ>z��?3��d����ߘ�,#6G�9�:��l8���ܕ)��4
��#����
?+}R��<�������H��*�t����|�:!)\��B��(�$,���4�p��@��Q���G���F�
�!>BHp�`�����϶ƎHU�⺰��� ��Ȼ�꿬{\�w�c{e���So��e���^�9\=�	���֖������@�G��&#���K��|Tf���k��`��a��׋C��<!�
��ʆ�nz��/< ��`�����os���ʾ,"v��'��%5��5h��Pͭ�9�W�"h�QlMMpY���p�������L<[�#kMɎ)�/@�̉(Y�Bs�(v�ō���i�<I}�m��c�#��c o��K��'7�Ё�(F(���E�w-�G�>F?���]!c�W����"ı��w�@�${�[%$�,��)&�a^h�8>��� �V�d���&�~/s��)\NY�v�d!ޥ߲��0�\�T��\�x-����}@���B�	'��舼['D!}َ�y��&��y:���'T����)�i�k� 苫8���a���|����\�f�'���G�u�������7�`EnW�rː:Yd�(���q@������L�?����U-���9�B� ����?��!%2l�^��R��$�ep�R���?d�a��;�6��3�/�њ҅��n�΄E�����oTDP��~=,X���8Q$������y���u����v��<�LT�Zf��Y� g#t&ð�_���X5^�gc�d��I0�?$�J�TOgw�H�h~�M��X��>�2�y�}�ASC+�B��/@�:ټ�%\"nfV�������!��A����ĥ�cЂ���Q9"�b���F뒝a[��NDX������+d��_�S�v(*�3�ó��#s� ��'��#�4]!�F����YlՉ��I �j�G�m>l�,�� �K�1ʘ�c��W��e.�%�%F����1�7�d�?^C�6�N���L�$1w�=1�Sj��b_V���	Ӭ I���15�a���/+7`b���^�1Y�Hʥ��G��$-����-���h���Z5�ʬw�z�t�쇶��e�����P�m�v?^��/����!�8�v��z���*�c�cD�P᜞��l���j��?;�X%��.Q3mth!�m�ښ��DA��ʖ�/��<��
2Q�fƤ�kc�@�²^���"�F��u��Cv��|��p��F;h�����Ǽ|���_s��ڼa��D�>yq��,���wP��`k�i�5B`aB�6��$OD�z��X�&��>�*�qoA���%���<�ʰVc��<����l`<��H����er�O�	䓄�{�ЬrpJp��gXVR����� P��*�E���&3M�G������~,��M�QX6����7�$[8�H��X��/B�� ���IE�ϛ౿iNϻ�O�P���	����^EVw�������H3
T�^��0]�,l�b�p �K�p���Fў��!���V�-h�p.x��~�&�g�Ǻ	�$π;+�|Q��n0P����d�u2	�٩��	�̀;&�X�{����)fc��3uȑ9�V���D��Κ"�<βDeq�f-�
Z�uj��h�/��Q�f�w��e�i�:�7J��h�Q04�������vw�]� >>B�z��@�u)��)��#U��N*~G�B����}F�U���O�^RA��&y��ݞ;�� Y���_
�4��ߑ��+���b��I�����2�]~�z����2i
\O��u4�>�3�W�3�	�Ӡ����]��
}a �*�Bx�aeп�2B�۲V`��L�	u+�7�7p���5�Hԓ o�d4!�fL��h�����i��5B�-z�U���%b;�VBj�D�F���>�N�3������P���H9��r�ƞW�I��F-�0�/�}AsSU��d�#�����T���[e�L���L�5�6�LFh���a��b� ��Ҧ�����,�[�G�/������k��o��Ũ�X�� �LW��F`Y�^�Ri�p�H)l��j�Cɡ17���<u.G=POtp�Q�Jn\�鲀Ǔ�Eo;I���1��e�$C�-�>����
�h; @=�.p��� �ėo'-��3=�/����CjT�qr�	h�]�|�J�1���B��
r'���Vd	Ƶa���ý�����Ѵ���n����\��Lk|VS�c�������y3�:�������m��e��Q���i�͸1�Ig�-g���0���wY������� ��<@�gb#���t����Ъ0��ktD�K������S}�pߔ<W'3©�跾�另�h�/�c|(28���g����`0��o��]&���ΉI_�}բ*�mF�[n��<W�-ᮉ@��GT$f;o��B&̇�OD��k%���;�.�]C�>���K![�7��O��>�'!x���P�a����?���l��y���զox�������(���H��+Ib���H9�����7�[�/��Se2��DW=c��~���Hƶh:P}������]�{��������Օ��v��&FﰚF������'4F<�6�;l�d]��g�t��n��`_8�����N�{�]F�7D$������hY
�<�?,��;y��d��wƥ��e���^�-S��QO��C>8N�G��E�}C?��t!~�t�L��@�������?-��Q�<]o۲ڂ�z'�3��t��?{G�����m�b�+i�;����]��K���bgu����x|U��!a���p��N(��&�]b��c��an��? ��r��ŉz�g-3����3�NQ�%�-~蠍ϗ�QK��Y�JE2��-�:\dR�3<ā�R`�Y�����i6wG`V�f{��Y�biX��_
���LP�H?�w6�|�n�ڞU�_w1��=͕�̂�����=�o��\>K[�֥���qd�Z����;;�EV2�t ��Y��TYs[�c�C{E`����t�˔D�?���`	T�33p�ͻF!�OL!��:=�́o=�H����(��7S�@��ͥ�:��C���S�? �}r�"�n��q�ZL���^�h�f�<6�V����"QA3��$s���5�adx)�Ҳ���>�$���]�'��*�s��B�����~Z�a����T���cFG���J	o!�b���K�)y��V��&]�=]�c���_�?��k�S[O� {A�����!*�"�R����.�%�͹Δ7�ŭl���bR�E�C|�L�����N�3.���caNW�/��'�?�tY�J�"=H�5��D��U��׫�&M�8C~b�<{c�;���ӕ<�s��O��-���-ƶ^�״�^;'^�;.L`��-�[sCnR��	Lw�zZ]�H��&㩧dɫt��}��x���C�Kut�Q��t��_F���U�G��&K+��8V=A�ћ��V[�!���!g� ^�ka��گ -\P�߃/��\�Fz󩢡�9��&|}��
�M&L�C0j��ͦ��WGhY�qjP�,6��
!	��n���2���&�i��#�ĩ~�Bؼg�>iT}-���4��F�oC�W.k��a���_���S{���4��k�>����>�ܨ�"m�S��Ϻ�\꨸���-����b3'�'H�ju�h�\$ ����e�o7��AI�思]�Ѹ�GR\��3�@d)Q|��N/��b Uԗ��	�͍߮��΄&�Xh[�?v�"�p��n��p��C3$��2��D�K<���N���1V�W��[�o�s�R���{�#�Yp�{e�b�n.�$w{���]
յ􈨁֞�P�?~��2q���u�~;S~���{~	6;)6];g:����D��6E��bSdi4�y0�������*������9�z�q�^u�e�t�� f�,�5����"����|��ݾkEB�Gn�����5�U���;�2��}�y���z�ωڿ��-=���~���PEѳ�F5��Ykx��爠��z��͝?U�Ic3���
�k%���������@����c�)B c��"!�H�І+�?wV��;o�G7[sq%�7C���a���-�ۺ������څ6䧥[jpi���#���u5�`C�Z��j��6���ڲ/��\puv��6�^��{�]W+��{�Q��6v�(Y�[]���r@qX�Jk�D��Ԗd �Q�
[x<I\wt`a��'L��b:=��(OA���&d�Dv�)�"�ּͧ���ZF7&�)"�C����������i����}j�W4��q�f�%:�
K���<;��z�6T^s/��,B#����̗�	���9��z���j^�VL��"ҽ�bJ���J����˽I.e����*�ᓓl�{xn��i����E��l��9 ������\/�;ׇ	�����[RaN���*�$G*�*o��9gA`ǂ!��p��l����\�zo2����٫#�+����׎zcG�+H�B�g�Y���Xnٰ���l�=��z�u��*6xՠǠ�
�!��"����0X� "�Mjp44�z�/��`'������2A֏ʄ.+y��X�{C��Չ����s���/G�<�^�;�!���Z{TC��v4�%��T���T��z�,�����n��j��.B8�{�!A]���5�!��>����<���l8�i:1�&���K���Y���C��l=�k����ԩ��ȓ�����d���ѱ�J�tA$�+Y�B�XMv��aF�Թ������],*v�s��v05󙌸_����ȊMC�܇N�A���b�F�(U���Hi��q9��A�(�}Z��e�3����0������7��2�r4J��ݛ��O��Ee��䊱�S7y}�Vf)�>ɘ�(�7�R��(;�	=m�����O��ȉ7y����\�K��u��Ǖ���P{�5�¤�Y+����G����\����������������[$�g�����[D��r���Х0P{���
��w���,�ʼmfmT�&΍'A�A�M�䗝V�O��3�� X�3	?R��C�����JE֗�g����H������z��=S?���uv�M��{�u׶CO��&|VL���/h�O�)zb#ogQuث��0���vF���o+ r�Y���]:��ub~),�{ey�w{�M@�:Cz��vZp�n��[4<���'�!@���8�1���D]�f��R����>�o�m&+Pd�K������řk��H~AVY����9K�N���G�$҅_u �B&$u��t����i�^����F �+DR�픈�J=|o�ۛ��c;*��I>U`�'����D>�l���7U*q�^?�M^h1�����_.���O���]0�g��[��KwW����=l!�xF%�/�`(sr?�`E."�%�\�ws&�{��o�������I\����V�"�6��jkh~�
~����rs��y�W�Ċ�v+��r���k'�rA"�}Z�I�,���T��FL�I��ok3X��V�ة3U�;����~춊��m4��o��S��$�5dD�`I�F~/�M��_�F����w>����E|D2qc3i�Ev��q�Z��r�%i�[�('����n��{+� ���*Ƙw����e���!.��o[.�Դ�D�炠\�ۨ��|���q��ƣ;�^TP_�͏Rֵ_�`���!����B�r�d,�n�%�
(d0�V�E�P5��] f,�9f/�o]n��ty�V~@
�c?�ѝ�K��g�g�Ҫߢ�C����G�{��G�1}W�(e| ��Y��mk��ͫ�\Ƚ��6$����q���y��e�O�Uz��4���h(���E�������XQ̈������ O���7�w��@�{�$D���&poē]���NW���ڡ�`~���=2G>�Nm�b�v��p`��*6
R�Y�a�$^rIXd
�Wab���?NM����v���ŊP�C ��v���� t��F�ƛޯ����Ϩ�f�\ l�C�.ӳ^��:�B����9�L��MRb6�0�7A��Q:��6]��=6�:��*l�zɿ��W������y$�g�����/�Q�i��t<��2�ӭ�	���\�'�;x����b�LpVG]����뮡��� #������4T��L�}�n������ګ�1f��ղ'����[r���UO�rh+�6qzM���,)yY\+΅�|"�0��a$)�}��$@������SY��n!�L��߹�ʙ���(����"�|_pc1ph�5,�.8:HIx]54	��k0X�矀{JC�]x�-��A֨�BK�~O�G�(��O�_�,��z���jh�s�4I������
 쥇yU=�q��ͳ�� �A�����d��(���f;e��VQy[����r�H1LQ���I����)�n��/�a���ʍ���,�9~���ᅃ�c��+��?A{������8�̤����1��&q���FR���l�������B��p���9PV�}ثT����U�����h��"������^h�I�L��K!π��J�^�H��h�
���Q���8����������<��	�2�2���@^���u�WZ�5f�*)�d�F[�d�-I��奴��D�M�E��^����T��F��U��*o�E�n�F������ly}^��\YS�����Iv�!�,�J���4��s�dּU�/�tm����_�]u���>��)�_%Df3<�9a8
��-�-�'����*u�U�5���h��h��Cű�9���.��#�H���F�;a��;;�D\6Vt�x:z·I_
�h)a^��=C\��ezYщ��C�v{��3�8٢��sݽ�'�B-���2�b�a�i���������7�D�	�4��B��E�k彯KBN��c���C�}��h����I����c#�Yzږ���,�RR��p)�Dۇz���/������(�$��em�� ř�6�J�ok���Ѝ4N�?1�mA�@hZ���L�"�4#H{j%���0.
D=�J��?	z�꿑�@�� �u��B�w���M���a�O�]ǠsCR,���~2�)��۟�֌!�{#,=���ex�6y�u����ϖ�-��{�=�O������s\NՆ������Qz"��7�����d�q�*&�<�;{Y-�Q�}�o/?���碕�@m��-��l�֝�w�y{Pt����i/��a-w���w�I&?&��o|,�bi�SG��\՘�}��˥�d�z�?�q�I�J<3�&�-���LD/o�BC{}��v�dQI	������ǒ��"�j�Oy�c��.�NL��gj�!��8���p��¶��7��<]��O���2Q95x{�M䇡��;j��.Q�C�ݢY�?��#��٥��х��Y/˄������V��O���Uk��L��y��%������[Sr ��C�M�V���/ӈ��-V���@u;�t���o7����t���34[��t�a�3`��~�*ٴ@���}Y���9�ٓ
b8�/D����[��	����q��t�#,8TP�ϻ�4Q.�5^��x��NM[s���N���Ed�^\�gp�*���BҿHO�;�i�؞8�v��=�AO��c)�Cp�y�Y��E
\~��慰�����������u(K��vT�a@ב�N�c�|���ĄU��Ɛ�0(b�w�v$ �fXi�	���t�bm��l�]���+O�� ��k��;2��U&�H��7�=���A'��Z�W�m���7~޺�	 B�T@���WÕ��St������>��*�X�>A_��u�yu4fw���AG����l��$�9�0�՟aj�O��`ZR�Cc9��P�Kπ��Hgܫ�Y&�����8��R��D4c���"����g#�-��:���iV$�!Ef*?-���QM2�Ql*0,0F�_��b�%�?˭�JU�����q[���\��c"0�U����[�kfݽ+m��$��da�n�������@ա�ؤ�^����!��{�T�������e���̼,3�綶Iix8\_��hN_O6~���+X���0��6�	Z*�?M��σ`~�n�:�!��S���	J�Z��#֮�J�lK�'��Ckf�q�Y�H�cB�I7��-Zk��ǘCP��Y< ���@��O'�>u2R܏)!w`:�<�+�z�U;���@��w�K�[BL�y��`�H�	�r�
���+�7�6E���:�O��������]�d���i�(8K*�b���O)���� b'� N���4�\�X�Q8�J��t���n�v�	qnk�>P�|Z�U)8��F/bW��/����?}�M�iK�I"􌳹n���Ģ��\Xh���/�*�CF���"]\b�"d9
ruKa�S@����E�O���4����I��T �`YB;Y6�����?���� ��<�b�tL���S�C��/ӭ>,@�fh$�����6�����և�@?�)`����l�!7$
3-��0����x�_{�(d������HN>�Y��>����R%#��R��Eo�z�A�'dXD��	��Z2��"��S,���f�'���?%i���v}���ÒL�)��X=�W~�C1��������| ���ʣz�;��Xɭ�����9]l�Se��'��r�5a�'#P�mа-@1}kH���)�:4�Zřf�L�h��N�nGzM?$f`�������r��EB���Ȣ�}	��P�r�"p+]4��'o |1�H�ސI�)�{u۟D��c��<��<$��#���N���t�;���la1dS�7��1E��`Ɛ,f���7�!`�4`�TJ��M�vG��X� ��a�$�i�x�Y|m�.�&�<�3��L��-6���Vvd�5�2�d#uC刿���R!�mn���r,��D��Ci�\�G"��)A��KMK6N��Yq�A5e���U-Wk��f��ҵR���w�U�oA/3�2�O���	Й�D�Z��n!��pA犽�G`�$�o�3F��F~݂;��w�1\��ל��A?���epۢT�3/{��H�~_��w�]gQo����~���V��,�98l~�uJ(�,b�-)��_LK�)�,M�:D����C����"������9�>��#bL,�dA�zhF]�Uu������Ѱ�>�/���y'jj�f;0^{J�ɩQ����a�V��ui�N�z��ħ\:}Z�[�[��Z�	J�`�i�V;A��H�5@�&����w��~���Wq�0�jEp>fVG�f��o#x�ž{bl)kb�WB~�P=Z�gz�!��	�Yf`��Q]����)V�}�k����gNվ��aT�]�<Kv�%�R"%�`��=j�	��Q�@�5�WT���Z�2�,����ϧ�%�i�
�i�Mh��F*�R�w=�Gkn�/Z[��{lk(�Y�,KI�[ՑW���"��p7N!V`�ڴ�WN)+�(q,��s��,�Z��cۡ	��<��L����o}K~�^�����Nǭ�������@�W�f��/�um��������V
�)��.&^+x�)V"
y ��ɧ��7�nhz_^m3Ld����_;�a@��㴡��&�^���Z�a��9��n��*�X��(<B\�z�
�7��w�
A���pBo�6�O�R�.�L�ޢ
4��3�6
vM��Q?
��#�>�>�t-5z$���vnG9�E�+Izr�')as$v�;� ًF3��5]T�����*��ikb-��n�Q��M���gX4VN�B�L��^�N�\�;���Ԗ��Q]�77N���mm<��՗�3�ո���K���B�jrҧ���"�R�" �U�0n1����-.S�g��ʒkO���-	�%ײ^7R�l��J����*P0�v�l�5!�����*���W �����X�MƬ;�&�{���u�7�:�7�����ع��oA'�%��-1��k_�2�TٔWw6��.x3�O`�D�#{��=F��q1�x^3W�&��aD�@27�f����+���|D�Ynz{H��n_q��P�׬7Z�H�XA�{���C�"��e��)��X���-���wu��p�,u�7��#��+�s�A��a��>�N%<$���<���,n9��W(�+��A�R`S
'<�ma��p�)�.V�"��PK02�(�3�y���6c��<�:g�@"�-�͎�*���`���)'���}+��Dۺ��|����+�2���K�{�hY�nc���7�BB���A�KV��F����"K�&�a�#�EKP������(�XZ�+����N;I6X>5���Yߨ�#��T��9��*!�H[�'�|R�]Y;9i)=��o��Ig=����NҴ�D��+1J?� �z{�ul���ա�����Tn����iկ|�:�,A�Q�x��2	'N�_�֎�k�|���G<��� ���3BR)b\�0��q��]�Ա}d������d��{Ո���� ��"���G�ϋ�����!����m�dp%UC�� ��π��5��ܗ9�I�7���=i;�=P8��Y�U^�\T�`|�	�3#k�()f�W9#��%o�L��w���x	b�����H��$�-f���W����>6e/jH ��l.t�pK��f����\��o�3�Ln����?��m��mn8�@Dg(�8�
\k���F_l=��a?�C�������}Q��>/PC6��&çM|�?��cWJRZj��*_��O�1����#`<��/a�~��9�a
؎}�_�$g]�qm���ږl1��^Y�Uƭ�
|oJpm�:o�{ߘu�. �H��� �/�4��όkr�\9�N~����Iى׬�y�a};�YY�`Lg/dǠb�Z	6[?g��ә�����x�D0F�h�G�5����˵}a��kF3�-�����3sOw��} ѭjD���D0;oNUlP��Q�v���ټ�d;�<�l���""?]���[����xV�՘d�~��Ay�y�@R4Z�hu�����k���)X��!�pxI�e��.����Թ�KE-�)k��N���u�[n]X��x.~�{ۮaˬ�4o�{�x\�קGP$0��:�z��B�^CrGp,|q4� O#ؼW	nӳ"� -ݔ�tZ�]G�2Wa���^�K5
����$Z����øNr(���=�f5`$}-�l~~4��Bg?����i'fT��������0�+��f������Y,X��rϲ�aeXxG4�@C3=A��n�������S+�N�;�ۉ���O���*���T�����&�H^�<lN����lW�ʇ�`.a�~�wc/�2����+OŁB��9����i�}Ϫ�@��}t�ܔ���wL|0��b/޷�HP�+ӱ�l��b�TE�����s���
�<*.������r`�b�ZEVV]���E��\��
O.�
Ej�8��^`�Y�2l���G��b� \[1�74�+`m�񙥴TL�׏�&Lz���$|�F�4��hhB�� ,b5�n�ݓǃ���;Jj�p�K�C�&���HYbx:%����E4~4`�'���k]�$�3r�J5��ݴ�CDt�N��Gɸ���3��t5��[���N>�>PQ�y�Q˴�����<i����{��a��I��Z���{�΄ԧ^$ RڥO�ɨ6:�O���g_V�(TBa+=Z�CI�q�����Z�Saǵ'�U?÷�M_m(w���o�T�(|y\��&þ��u����i������{�{���|hA����Hk�hE����(�B�4�Q:���4r���J|�G�)�mgb�<,���A%�H�<߽yf
5�yD��h��Q�o�t���DwtpN�I�C=J��K�:D&����|LO�e7iY:�l9a"I����l�'�G��>_A'/����8�5[ߞ؟�d������%H� �w�=�@0��xb�&�%���G� ��L�����"���%�A��0�oP���Y_����9�U�<@��9ugG_d=.(@��p����f�����r���7/���;^5��=3k������+e�\�g5��,���ڂn��o�f�����|sv�-��VwN`�6�UW��@�D��o$�7 8B	�-��/A�̛$��s��v�dR$Go��+����h�\��/$�Z���΃4����X��r@/��a�f�}-���kڗn�$o���	�2Շ�.;�9�S#@�\-i�v(��rp�����KaǢ�4D~wM���n�	�Q�V(�-�d(����䛯$[��+�ڟ$�^��'�yy@�Ӌܫ�<�O�J�§��O��pB|^��}�xu�E#3�U<�Eom��y'a�
�vW��IEg8-�kT}�'p��`��)!v����lf֭G�����{���(Z�#?�6ij�aglpR7�lDJ��xs}N��'�׭��9��IWYD�GH��°jкL��)��H6��������$C����%^|������B=mUV�g{�1��pv�)?rq�?���-�&Ӭ�϶7��S������ۧ2�YQ�L��<����7>�b���7�d��,������x���R��*
chx��pXgS)^v��?��*F\dUV�-����m�pQF�����Z��ocSK�>X7�͠7F���'y8��*P��H�L��D�T�6cv:?_�ُU�U�� ���R�"g{U��B�}��Ӹ���b��t/����焭����`C���BhB�DB�@�H|�ϖn�F=�"܆�z0������l|�O�*+���c���N�e��rM�w�<Ҫ�Sի��8Ɏ�/TC�.?�7��}X�?S>s��
�����3�Jg���r���ʋ'<y���9oG�Sι�����iy�����˨៎��g�1 ��"gM�LA<� c
o�.�\<�{|��n�Y�;���J��G@M� s��`g>F���ڱC�l�l�Z��͈�:��I0��W;\4��h���V��P�i ��D"�� �w�CC����wA[,����L�хYd�a�ג2E���%
�r�$q��<N����'�ťx>m�!��>	w����B)̙�rؼ�B4tB =����o6	�@iC'��D-���IsT�
O��\s8FC�'>E�Y����(�f�/,���;[G46闭RB��6r�]�!�5 ګ���LqzDO�8M%w\^���aI�����u�r�W�������<����̴����#��4d�Г]Y�I��x,����1�z��3�A�R�ߢPz�<ί�udS�4�V��b`�N�󮟡2	��qVB��o�#�^����ۙ�j��dL���Fg~�����F��I�YU5��2�n�ne�p��EЎ4}0cK�ʂ���|bw��H�͡��Hg�o,J�ֹ�XE��'��E:�n�h��7��3��g�~����BP?����~��},&�#�����c��o���*A
Ա6\ө6��.��=�0��]���w���K���.M�F�#t��$4]�@��r�2��/�r|QU	H��U�$�����4f�9fZ�V �PR��$*��Z��u��#ـg��%�Y�ӊ2��o�6��E�y�3�y�!-�9�l�WvOINW���$���bh����Gl�2�韠+�|$��6�H̓�\���&-i��1j��݄�a�}/<�' X�}_y��?���fB�w?3�]U���K73u���K���Va�p�F�Oh^UzI�	Tә�Y.�}Z�܉t������:�x���=J�%ﺟczj�xJ5������46s��lT�LV B �E&�t<�}�O�1�^!�YfZ"�����w�Cd˞bD'eN�hV��`D3�XnB,��*��ek���E��*M�?{ZhwS����G1dk�,�q@�o\og5����c�4j�_�l�'n�G¡���Zi�m�L^KeoR|'��AajX���4�3���v��z���7sT��N�ˉ3z�)���L��n2T�/�$��R`�IN��w?�T�����@���X��"o�R��Lu	B�j))f��B�<��Tn�t����_׌���j)���(��N1�g1ȇ���*�2�mv�Au�i��lv��A\�#aSزP�H�Q͌��(�����µ2�yH3O݂˛�?��'�]2;0R��-
�k����?�ƕKCzLNF�������V[�bm�d�>�I<��x2�>&����d�1Vܕ5�qh
�_�~��m�����׶XK3�o�=�a�1�К
d@�;��:��Ȗ2b-�Vװ���WdR�����8���mX��	cy�]Utܧ�긻��؜�'�R�;�_~5=�M1��M���I�Yj�c��4g=���G�A�Tm"V8��O��y3��E#��U�E
o�+��To_�V���d����y�Nb��|<#q;���0��~:�s��U7x���e=m�$v$� �j�jC�e�B#3l�9�(xc�w�T
�|�-c�~6Ӫ|�6<��Q᫟P:{g\¤�û��P����Cd�l֯J �������q��k�Er/�bh��d�e�Ʀl�X�~���o��L�b�����?�-�k� ?��3m����a5 �q�"2�!�p�F�J�e?�q���
�[q_���+"�`·�^gqs��ɨ>�NMě�q��n:�.Z��-�V��L0���D�?����4���N7tJ<<�?e�*���7W��W��o��pB��*��� ㊥Ro;?1p���!Y�"mOǙ�{���� ��;�Ӥ��m�u*l�v�{%g�U{��esE��a����6:���n?���I�4{��Ƌ榠��cv >*X^@EZB:�Ӏ�*�J��,o�g|1L��Mv��|J�1�C�ϔ��t2�$dN���@dy	����%������X�@�IO�K��;�@nk�C^���.�n�No�o��@|+����M)ʃ�n�4$���D�U��d2 "|�)�m}5�r����ʻ�c��� �*�L���W���_7.�k��Iҽ��	sa�WN�tIIY�q�����}m(Fk6���8CM�2L�E�]6����1F/�y�S:'�� �ͪr�����a�Ƒ�o����8�Ѩ��WĈ(�U�B)�������f��S�>�牕=azne0�X9��#��og�q`ݾ~���+�İ(�6k��_�Ԥ��d4*.�I��H�.�Xj�W��
���|�NP#L�� 7�v���H����ZU<��2=j�ޙ)�dl V^�J'�b���u��u�ڲ�Q4�J�҇���c�Aؑp-Ė�n0�ȿ�=����L�"R���ᔠ�p"�i2��'�%�"@q0c�s2������v���8�d��0��u�9�����m���KY�j���	<OҠ�`5�YY���[umt�ӇD���,~�;��Ǚ2b�PzJ��3��B	;�,iOļc�Zo%�h��{��7x�C\N�$��,����$����K�Fe%v+ﷶ(�A�j�!F|����I�0�?v��.��$9<1vo����KK�L#���b,k����/����AmV�Q�|��i7j{r9��� �O�N�����.l�H �v6k31O�S�8�+��vܣ>;�y�"Nق7?�� ��T����C�zu&��U�^
@�s+�/6k����z5,�v�IeI�]R��V�Y���1�keݒi�t�����ϐ������O��z?|<n��22�ɠ8��^MK0;�so݇�x!�7��s���K�c�D%k6�����uE^:�T�韑Uwgp��J�즑b �Z 7�

�Q�p����MY�s�U��:��}Q�d���+wF���ˌ>G����Ez�W��죠����9S�ڰ�6���a fRI؀�j�r	W��(�m?�~7#��	1�[v�<��
����Y�=L&�����&�2)�Q��/�������OP=� tb��A�h�Vw����s�y>�{^�0b�( 0�i��n�k�f<��Z�;�@»�7'"\UZ��'	�D���T9��ܺɂ	�/n�n��<w?q�r��o����@�O��T�vb	^/�CV�4Uгϣ��d�8�y���[�U��~4��*VJ�z����Lփ83�=ߣM�`b&)lt/Wp�$�݆�dމ��ۢ�bf��J�D����np-
*���Pt;r����5�X��$� ��&(���8@��o�@�oO��k�K�0��h0��9aB�5�)�����4�1.2T�du�},%�.�ZT$�$U#w(����D,m~�y�`6���[�6���a��$����@�{��,OM8R=��['����(�]�Wut�oj��wK*|GVwB@�F''
�։��ϫm�v~]�0@���K,&�z^cy�HN_�8�c�s?��ښzJ;�8�*�����"�-]aј����G�w��&3�a��1jS�u�w	�M��,P/�m��f4dr"ҿ�Q�&�����7�&*�$Hv�Y�Ը���[<-�5y�\��ӯy��A:݊��������8yVI-y��|����S��� ��t�~%K��,<d���uc8#����V�`t��tU÷��[+Җ�Tz��X�����Z⶘�j����)������t����#�6�����s���S���K��p�T�?�վ�I1�/�7!��Eѧ�f'8���S[K�h	��c�J��nO_��
�BaW��U�) J �̤D���C?�a}"��Dۣ:EE<3�Qc��E�z�^�i�K�ּ��1�דm�d�m���ᔠ� $a�&�I��K��|Du�������i�G4^�	�B&�#�GB.|WE����7T[�[^�w�Y�/S	���+#���{�k� ���-�J�z#�����mG$����(�y��`i��8�!R�'�.e�+i8�E�	�'ǲ#ι����_�u��o&C�3u���I��t=�.W����g:+�FGIi���!��6g�x��<�5�gZ>huN�d^�%H���h^4w�M���K@�޾���>����C؜
uu��̨(�3X�^���ú��0 �m��̼8�Wm��Χ(��%<�>�2Q��!���uK����e����`�H]R W��z]�1=֘�:�׻.�-�2r|���%B��?>։O��znD�TJ�Z�N'�G�W
ZU�c7��o�����y�E�B5\�|�˘A<�6Q4��"u� ?�!W�*��"l�$�������@Ȟ�����0�˩���,��)�r��,'���wk�����i#G
�H<�s>Jʖ��.qv��\`�>8?Yk��"�[ST�!��ژ<Avi��4d���z@W�z>߲"��BnN���������贊�ݢw��B�g�˙�tq��œ�.��1Z��gێ�+c_��� x\���A?�Y�3	vu�f�&�"h�K�PҡMQ{&�{�̹A[��U*}��	k
�{)�	"���}���"��+�1�*�P����:��sx�%�S�Db}}e̾O��739=��BL�4R�R����T�@b�`��g�{�֜:P3�%�?z�Wt��*~��=��.�Oe Z[�b�t�SE���5.,�ڗ�b����߭й�\5�&�\{�sv/��oZ��`A��pMbL*�4Cٛ�k�S4�d{IcB'�(�Z��fS̃i��Y����S�f�n[��Jgפ�c#UUϊ��F7�gu��W*�/'�5�c5,G�x�q-�ՎB���x�M�=Е�[��4�=꧈�`���&�Y���MLU�n�D�	̑8Nn�:�Ն޿73�&G�!�#k�_f]*�Q����z��0{��ץp kcY.+�l�K
�����c���<8�/I�:�E־~m}(�`�;S�q&���5	$K�r�*JDޮry6j�[t-`�_�M�/�u�JL��y��4��z������@�ko���`�^�_W�-���n��"�K�1��t&³\H?�1��K��ƣ܀��a0I�����(������uJq<��wKd.��q�#���ɇ2E���TB4��3fU1�ߌ6�/�AT[�d<�>D1b,;������}Y��/1�s���E>���8�';؜���4�Yц�ƶĭRFzDma	ۼ��W-�_n�xB���{��U�y:�x��>�;0 ��}��၅�1,1�T޽�)�x2hl�Ѿ=Yν�L��,u���U/���1+Ѻ�`㗍	h�i�,B�}�p4x��7���5m;D��qbޕ�^�V�.Q�#7b��ܴ��H�(���ǖ%��4LI��� ����@�r`[o�����z3�Zܦ��t@A���޴�/;+C<N��Q� ��u�k��q���nbY#}���������cG�OU�6	�@��  K�Z�6.�ͽx)a\��J!�z���M��k��e��E�hu���d��b_�N�Eᅮf�tᆮhnMh���s'H����/��'jߙw��X�z8W %������?�<�Q =�{��;{O���j���k,z�-�f�Y���H
Q�,k�"�"D0ǹ!�X!�%[�ֆB�N2��^DAG^�oQ�:U�h���Ў�J9��*�x��a��W̤���d���=�϶���)��Tu����rL��@jl..L�ygm�2�I�������ah!��V51˻T���J�#\�RwN!m�T�>��z��b+�R0���S����;���1	���^!U�2��Е�Ĭ����{U��Ľ�(DB{^�<80�]ix=�����9��P�������h'�o�[��%�n�w@�pu�o�[i7�rp�E�Q0{!�A�q Њp��Y8�����8H�x!�����6{�|��qoD��?�lWuԝo4�G�p��Ø,a����0Ht9���o�IU��V�����!f����'���e��z��/��?۞Z�%����Y�E�����߁$>�m�N��T��ʯ��P�{8d������J�}z[�Ǭ�@>w��;(�<x���q���m$�&�?�"�9?{ϳ6sﮆ� �6xN��� ��@"��\�2���o#��C�7߷ŷ���8�J���֪}ߝ���cSƓ8n&hK�%"���l��'�����-�~�+�穣�qk�+d_K<�\����q�RD�A_��P%�!2��^b�(�j[S�a�g�����5��X�$�~��:ng�+n<�ٜ	pd�e�]ZR]ɞ~֏`F/�n���al��ܧJ+鐀�i��E*����"cE�'0gLD-1�(~V>�+ ���2�D�゛ґ{k(���+3ͫ���%�-�f�k�쵑�M!'���a0����ɨb������q�N������>����Q�'�	���3)GYWe2R+�pq1�[Ah(Qj'�|xP�;��F5ʙ��T�*8�/,���6�%�r(qZLuG��)��8E����\���*r+y����>h#Cq�U��a:��y���,i.n���[�	���2J��!i|��%_���)h�����K��$/C_A^��+L�����E�9!1R��!;�O�I�e�J"Ώ��J5����&��K�Z8��8h����Z4ulо@�N��E�+�Χ�=հ�Υ$�N=�pw�E%��Va �P�hL$�4g�=�X���v7A�M{aO��f�}r�!�R�r�p�Gn�Y���S�*Z�$I[q���f7���J���>��,��93-bǯ$Kc�Ǔ#{�N|�d��s0�Mm3 ��x��Uj�����5vB��+�L�Cf�n8�b� �N�4��|!�t ��w���u�<���	w2ɭflp0�CU�T|��M �c���$B��e3���V�����i��;D����Bޝm�|��xM#���u�#�K-7��X梡�[�\���1m,�)�F�LR��P\6k�V�_����,"��%�i�GD����/��I�մ��y}�����(+"$��3����a�KS�y�����\Ҟ�)������լ���VيfQɼ~��������h7��`��B��b�	�1Z���#͕�V�[t�j�lDqn��y��� '����'#t��:����:��΂�3��qg���	.��Q4Z?'�.�0O��s@j�%3�=�0=���n���v��)8�{��MȀ�!�� �G��n�b�$����8�����������	��󍛉3�������<��q����߉�g����9V@�f圃�����`"���z���
݋ì2�ٕ���o��*���gd��@�\u�#͇���G5�c���j\�+��5b��.�s�j!PQ�Pm����2�"+��n�(�;x���c���F����-fٝ<�x-w�1� i�2XC��g1����	�(�G�{E+ܝ���7��o߇9C�C�w�n��R��$ߑ�7�%�H��uῊ�V�ͪլ����qb���#F�Mt��Am˨"����\�w�[�[MU��n�E��dyi�U5��9\夥� zaՀ$�O�X/��+�k�um
+Q���\���ԮY��'���W�3P ��f^����m1G*�1����	����>~6³K0��4#c�ǟ�.賆5�uZr�� �C^�lԇ�IV�����k'�&$�0�g:IC�y�I6l}��8����D��/g��˽�"i�@k�T�}��"����b�EH�<q�q�) zs[��H�:�Ѹϫ?Bp���d��[qzV�(*ީlp��C����g���0��M�'�&���s�&�t�PCa,@���w�]�S���s}��r,F`ܯ�f�Y�������gi��i
�)�u3X��i-��_����٪3.ˌ1��^Y�θ!Fvu?�qm�Gé!����{O�i�iߟk6�x�.�ؙ����N(�S32����bIG�YB��.�fT��*�}lׂ�OH�0K������^�{��ﰭ}uznKXa��\3Q�¬�`Z�צ�A�1�eR�Z�U�������~'?	c����X��ց�?lG��;��/*�D���r��)��*�zJ[������9�����nY��۔j��	��xz^[��-�����;�@�0-��z�=@���{kP�Կ����_��ip��Dy��؊
/B"����{u�Ļ��@��1�KI�����R�C֪������ K�c�R����?�:��윣Y�[�����C���p�����x�NL��xz���O�i~"@h5Vi{�@�򅇼��s�T���F�����W��߲ӴD7���EG��XM����6��;�E�CM_#����v�f�������9���l�EQ{w��ƕ ��&m, �?�t��E������C��%�w\҅�#�_[�7����l�c�"�|h��(>�o�u�H�i���Yt��@�Z�~L�sf0��pߨ��X��~����K|�ڡ��	$�~�b����7�G���V��܊�y�'B��䗦L���(}�A�Y@+7.w�7��+�~M(����}��W`�ȎiV.�.�Y�ߏÃ��2͆� ��AA�>B��}���/$Q�Ԅ�t�����k�dʅ�Z�1L�X��K���PѤ4ĸy�8;d�݆�{�mk{!������@*lQ>�FM�
v��v�k��ܵA���f\��P:����h�-�����Y�h���~oh+2���$j5��`�c�����
�*�\��%Kh[Z+�❝j��K�hը;�� �!~I�+��1H��E����#o����Aw�,%f�1�������,�|�I9���ƂWXv�^pqe����9ɾ�Q)�م�w<�7�l#7K�,���݋��a�� 2fRD�D��d��3'�t�#��Szf�Ә�f��2Vh_{��8����5%"
�E�pJ��β�1�
cw �9��e��F�Ŕc����?�!���cٯ�b��Ux��h`�*GLn�I^�ݏ�������/ƩjE�9=vb\�@;�o������rC"H e�c^��|�I������E�QJ�c;a�m,�#�ou�:�9D����ﮂ���K`GU�
Bb�	��{4F�	����m+T`�u���������u,g��9Oz���!���&z̜�)��-@��̩t�[m�q�t���`��d+��hx����Y�C���O����PI��.y�IA�F��61��8���D�D��IQ
��?�)�|8��p;`-7r���ϗ�Tɛ���e�����~�sJ��M�{����io���3�M�Zrz
؏��	,-��97<Z��6T�O�x��Ej�ݥ��8�D8����e�8~�9���D�}���I~�Ю� ����y?���byfH΁f��0c��w�/9S�w�ʅ=]����]jV5��i}���' ���q2�%;;2m�Q������)�Bܭ�ec���ԧ��i��j7c����0��LUU���9��G����U���z��z��ѝ7���I�@��͐*�,9ք���Bt�I�`k��TX9�t���/��t9a��H����-C\h���旚�g*u	�#^�����ID��U�����a�@	O�2�m},WÀ4<ǲ��s�[!4K\z'�[R�:s�Za;�B]y�9C[�0!�����g d�V���]z��\�ص�7�?��۞���Qu��Aw�Y!����b����1pE�c8RMԘ��&�7�(���������[����D�܋����n5b�^��H�B���NÔ�/�
�e�U��E����N;�˱��73DԣNo�NB�щ�~�̉j��t�'��=T)�J}�5;���{���ݬ�)��_Ү�ܟͭ�V�0�.���{;�l
��J�G\)�5�.ԫ��]գ�)��6X�f~�$���c}��z�mX���;�5���WZH=6c\ѯ1��ZB�9���_Rj�]�e+k���z�������}00��LO�*ɹT>˃�[��w���SrN$:� m��@��P�=zJ�ajU �@96}�*�("��L�B�e�oO�M�5�ܛ��L`�%_ą�&�j+�
Z!h��`R��5ٸT/���H���2�$m�fM֝��+�W�{Çh"-�V���200s,��U�-:q�_ ���5@�Ȯ�3WW��kMF�^˟�Yz���;��&�j�uh+k��DYF+|[nh����.�rP������] ���7
]B@
G0�@�����,����P�im�7�� Xd�7]�jk�|t,�ui���C�y|"t�n��^T�#l�6yc�{R���*?l ��H`jī�A�<s3���*J�ДM,�B����_'��w���9�����g�|XB(Ҟ}�fqW�����-m؁e퇦>_�ކX|a5v��c8�J����z�P�N��M�>��}��I�I����7����jL|�{4��G��-��A�ŗ�_�M�(�����	*�!�d���J6ۡ�kSc����д�K�j��f�Yu�|�8��@��K<y��V���Ҕ���.�Rx�!sSnE_����ُPܣǉ1��@U��fG��P*B��i}U�����%��u�����k����5@O�t��#�aȺX���C
`Eٳp�$EI�ggO���i<SD���=��d�3���k��cQNU�F�����O"l�Z��#��Ǜv��M�~6F�s�gLU֎�s�q�;���\�2z��%�KJߐ>��*�>ubC?�p���е�Է�m�;��
%��J�k���@w��\}(Dv�k�t)��x�^{Uł����Һ��]剰��D)pR�OfbS!�|�A]Bΐ��{��7�X����%Y��4I"`D���Ɗռ�� BL��H����	a=�m�G����:�.�w50I���֧lva�;\����k[�P�h1���B����i;�}������[D���p��!���G�q��ά�:iUiHE�|`��%S�4#J�~W�l�I�Xs��Ĭ�	ިi~��oS��f�^`�6	����k��6�%?�>+���V���W�ɟ�z|�1GM:�)�
�@]I&8���wH�$���F�Pq�VP���s�!�QD���?����2��y;p��>{7k���X&5� ���YL!5r߈��.�â�!��Rb�|
��E�?8�^	�!ȧ�_5�h���8��8K�iQ���@��H�MV�6�͟����\�}�����,�CȠX��G&;u�-2 �ͬ��o��Xw�@�Cө7~��%��7Y�g���{�����s�tp�s
'�����ď�M"*��S�H,�XRQ��k=�0��\<�����׀�d-<�7ѳ��%�.������cˣ�Z?����Pp�C�'0$��}LM��Msæ!H0�?s�[�欫�P��
xy���Y�c��f����0��-Z#�$_��l�8V�� -p? ����)�h��˱ݺn��J�^��#��:��L�ğ%\�B%��گ�=>�� �����4��A��G�z��?`ȼ�5����ߵ�z��a���K�Ȯ��jul�74C̼��O�L�٤��@��|Q��U�����h�l�&F\��*���MR���B�����'nr9�h�T�$U����^[��55��]�s^�N��䃧���J<AH芝z�(�*>��g\޾����'��Y))�3*T{i����_�]��Y�*(��[#�B�i��AO4�����n�8)X����߹p���/�(r]��%�O�r�ʰd|�w���!�c#�g�$=o�}���~�� ,Y��O��0�Vwϻ�P�����m�BZ��p0�LF�M)4JB�^M�T�X���#�=��^�P�����n�V9��̔��{쬫�w? 6~>���	-���cީO	�-��	�7�=g%��fsQ���X2�QC��k�DS���؋k����m���~u�h������4�#����Ƿ�Qvւ���/@��>������J�	�ߗ*�D
�x�|`|Sbi��%���U� !��顉M���pX���g�iR�,r������r�ip�k��9ȸ���M���5#b��3���0��Y7�GSKk���]�ك�w�B�|�yBH�Q�EԶ��O~����,�'�R�u�k�̤%hs���Sf��D����x�%(��d+9zV!!��J����Hj(����Ӛ�(5��)�(4�e"��;׭�Wb%z���.�Ӿ'3:g/��BA���b*�D�+$�d�R��\ccq8���-���&5L4�}�E��Ƌ�S��Q�E��Fv#!��;@����E���C�c�Ⴚ�hGh>js�����fԓ~`��uJD���yN3b�y�+��Él≜�G$'PΚ������Y��MOd�*6f�;�Q����虉.W���� !���
����1c����a��D���c�`xc�nv�q�ϩ�Tv�.4*�c���m�Ru���'�~w��N}�!��O�U�ZU
R�/0������U$0�A�iR�G�SH&��a.9$Vs:_sg6��3�7O����o:��ӄ[���*���ng:"�����y$?،�����/$5���ap�q�4�BnLk��FgX�����le��E}^�A����eM��S5�X�֢# ��n���O�0�N�����|�5�vP�j��SN��`���O|���Q�Ħc$��q�������^2��6�[��#��dH��aR�;'���PV�	4[z��dEJ���~r+�s+Xlj�m�x䑅���&Do��/"�^��ɐ���p��aLO�3���~9�?����Zst'� z�Y=�yޣ����*���r�nv�BB���/��ݵ���[��lq���ct)ȋL���B��](��0�+�k�#���J��V����c���`4��;7��[���xf�-`B���5��׷A�s���hx���!)�g�/��3��T���]?w���%�c�[�>��Yz؍�՘�⾔{�����(1�(��Y=\�µ�^��4�}ki��[6��R1A��]8���)���o*[/՝�����n~�R �'[�_ 눲��{d�Q�zi'Zʝ�k��zjk(�ԥ�e+���A:;�B,U����'}[�m+�v�23S��/߯7�kA_h��O��w�P�t����WHy�G�L9;�D�i�i%��R`o��j`V셮�A�{ɉ�_BeCϳ�6g�[0�e�N�	h �*j����Ɯ$F�g��넷����3Ě��NI��l���J-<S~���l�K�{�%�"xdo����<�PC(�K���N>�Z��dq~*�{	֔l����/sg\����E�/d@	��+�^��^Pj[-�8�$s�Z]L�XEC��r��_��6�>��(߇�÷$>�fǝ$��E��xF!CMz3��ڃ�I�AMV�a�O��"U��u0X��/�$�|�Z��㲓��|_�)w.����KC�{�;T�*O�A��gP�u\�0��ѧ$BR���P�2*����c��o��v�����dn.)�$��$��[k���+
�Ml�H��,��.�T�z���r�ԛ��[9!�˩����S����:�(�=���CD]`>x���4vf�C�mK�3Kv�J=>�n�z�9�LI��29�F��V(:)E������m�\^���0gr��k.Tb�������yS�<�*cO�9s�������n���F}�>������yˮ��C�N�mU�DYz�0�R��D�]h~[���[F�2�p��̼�fw���R�|Q��+�E����:��#V�[!	T�7F5g�*5q*�Ɩ%{}o�ˏ�b��yw�$T�1�^\�9�(v�]h��*�vkN�v:g��;�K:\�-j��FP;�Q��ܹ�v�%�)2W���
�9�o�_i�>���='�ꗽ�����ԐZ�7���
��D��M�pۤs�#���"E �ޅw�U�L�$����ro� �����oh��rxE�m'���&� ��7��;��0w���y  �P�5J�s��J�P}�ޢ�]��<Э%ʘ�	C�[�`�;r�^��Y�T
��#""��8����W
O�֞\�*bѤ�?��{�|@E�?c(�~��L��rC���U��&��6:t��f��#"�h�3��4j+3�Ú~a?��UT�|<�<��@�r�n|!�z]#d0�~��n���g�}�T#q�|����\YjR�A�n����
�Db��z�g˩�=4ɭۅ�1���v��W[�H�w.�S%����Sy-aQ�j�ubⰜ	�^�[����%��/H��8��?�x!̉�-l���+���]2Zp1Q����?��Ǖ��l0h��Cϟ5 ���	�Ż	��M]�/�PC+�K:�ޛQ[X�N�L����n��k���? 7���5�o{�)�5I�����M�!���iO��a�7{�9p��LU=� Y�?9�]�Ǜ��{\e�dʋ&#?ڱr�����rx�F�R-���{�4�t0�^:�Ts���B������1j��|R�0(��H!J�PYh�¡#`���WnĲ��3�‑�'.he�c5�kg��f�C`k|0��A�ۄ��.��>$.�۳���l����$���.�s�o����<�����|�?Ġ뚏c]�OΉSW�(L�I�d�P��9�h���2��^�V�Lx�`7�c�����6�&Ҏ\�윾�v���V>'yduu��#,�|�NI���I>�UcZ+�C��Rt�J���&�[G��ґs���mɁ�$��<RWv�Sf!j,�B7���m��0)�7��&�J�ƫ�2]����Y։2���y燺�;&�߿�%t�I��\��S8���t.VY,pم���;��Ą7�O<��4-lY�:UHB/Ϣ�#Ґr ��Z�+`aX��|�����U�A��-�4�f��KY��N�?H��_!#$�YE�R����;r��Vi򘖥|>nJ@��I�'����s`N�f�È�;#���=��>Ե�E�;�a;�޺���'���������Ri��m2�4�P��}<�{�g8�_Al�����Bvx(��YHB}C�$�d�����#���g�/m�.5{�u�'�GW�����6�va��C�r vF��Wv-RL�����E�T%����\
�Ю�jUYz��3�C��W� �s>������=�����mA�e(�`��p�.
���^�uȋr��Q�p�[�[N�e�L7q=�D����(�#����dI���ô��h�.}�q=��K�uݔ����fP�g�2��\_Փ�13@$���SaM����J�Ya�d��А�Q��M�oC�x_����o�I���s�/ۮ�ο���[m�����J+���~-]��W�{�n�4K��^����&��~�29��؎na�KF�hX~�ד_���w���"�)H�����Ɖ^���Oz�b�H���k���co���e��I�13�L��xH�٠�o������w���;"UB���d�;[��5�~ٱ���b Pe�<�
����1��e�U��L7mG�OТ��O�j�~ )��1����f�$"7�vT��}A�=�R��|��@ook˟Eg���wn΀�����JG� ��H�집�~ܩ<��Bq%�ߜ5"�l���]��-O+�Ԟ�ԭKOVQ�(���a�vٞ��j��	���r�k~]�{��O=�z�.���y���,����l)�*`[(��E��n�F�w_5���0�J�� s�d����N>�����ƣ?Ub���>�İ��-��|*i'4��A4��2V�t{Z��C�2�	�y�.M9�	�@�D�a��'��9�^X.�MI�=�������є��>$�ɟ���9*w�o��!׀�j��r���]�i���f�0�>KO��=o��D��	�ς ?5&���.��9#}�e���2�5�0*�%,a����?T0[�Jt�{��}��.(���[�k+��`S����x��zE=zSwB���[(Tq�<4|���ഓ:���$�	�ߑ
��j���܍N�]�5�xC���b;k�q�4ص�Q��;��_(c H��|q��H^�֘�0P���r�&���º��5���g��s��0I�P�2��~Ī���5"����c�(I;LJ���������2�M|z��2��W��]�G�W�;B����jXE��c����d��❅U��D�_��&߄�gr��;�hD.��'�Қ��9��ɡ
��M�b��ĺ�|�l8rv���9��{�zg�9ۖ�_+,X<��,�v����d&�Pzh������ FG��S�H
���V���ֳ�$�����BP�&]�+;�;����*��KDze(^�鱿uL�Ho�
ψ8*ٯ�mPcs�Hͭq�Ch���Xa#�!9&�=Ε��G��̢�8]�¡�2"|�_z�Ș���K���\i%i��j.��dݷV���"n��f�󟒟.�W�+���?PT_���	�Ig[��[�A^c0qX�k�{;��7������9f�_ط�n���9J���9��$g��'�N��_�{�c�4yܔ���k���ͼǄ�)
�b.9rHiF���q���z�<��߀�U���7�~f�M�x^��a1�[��nr߀gt]<c�`u�hċ6.��"�=kn
�����`��&���tR��<�j��O��M��L��;�\���Ӏb�)Ch�n&"��G��'�!El���8�������A�"֞��2ΟBa�`�4�\~�nw�����<tQ
~� ���C�q��N9��2�Q���h$%Z�v��..*���E�&�p����_=_�&�!c�F�ڏrS��B%�<Iz�M��Q><X��{h���G��UB�l����ܞƀ�{T�v�S͍���ۼV�;����"^P)�����@�JZ�H�US�����`�Xě|<��y�+���������D��&�('����25-ۮ��:z�Q�2~�|����$�L�%
��0-;tH�9.�O��g��v;�fC�Z����x�>�pa�f"-�@�5��~�ff�|����f�;s":�9v�wBǢ�	%,�*x$8>��i;Zx9���C�s�Ԅv��մ�qN���\��7��qF
	
]ء�ӆ��{C����`m�v�\+�΢Ж�}�\>y>�#�u�5yq���o��v^���p�*�0Dt����X{���Q��{n�|�ԹW5�C,4��E1a��=��;�4B�auc��� ��kh[�8a0�b���(���	����jB��	X=}٭��:���}��S�(���o�>�n���l��I�l��W�&&��!�^�9�
�,e�å���:�u�-\J�n�w���82���h�:��:���\b��h�'#����U����gȪP+���n߆�,��ün�Ffܖ��	ؘ�4s�\��s$����CC�k{����YsۘXY�4;��5��fدeB�ș.3a��|���3�w��;m�N�� W<�?-n�g#���

�^c"<�b�۝*�
DԷ�t^ ��<�ت��a��b��lp3q��f
!�����ů�t��r����m���!��^ms��f]3:`tO�}G"C�er]S� ���4��(�\�bo��Q��B{����xn2��ΛO*v��"澶��� ����i��4�AX�"��L�@��l&�&9����5��O�xH�'.l���p|K'�Շ�x�c	��0u���Y4l���6"����։�i�;=��QYD��r
�V��`K�����e�&����( �Z���<�bVAfc�Jl!%�5h����A�P"��C���,ʉ�Ί� -�04u3��D�T��7�&8(������h�8�@����SW��1��o�R�XH�q������w�7M,#��&��ǂݿ����P?|b�k��^f��K�{���|T�i��+�����cM38��O�;�`F��
�5�_� �`�#>��n�G.��\�+���ǆm�L�>u4&�7 ��F|ʟZ����&P��hi�`�f�R �
A���0�;�6�論�o��P�wW�E��\?Z�W<#�L����;�|a����ºVKN��ڞ�W�Gr<ZĚ[U����=4%𽌅w�(Cl
����;�����٥�$�R��A�2)i��ǲ�Im*0V1�	�ОF{П�h�g7�p���W�@*y,��ޗ?~��=������)���)�˲����F���`�AQ]� ��m�2�n�P�$?�\�&�����8�H�z�ͬ}Lb�w�&&�����Tf�#�6�034���1��I�*�>�*ݶ�A��4+n	iN��S�j�� �s�������9]0�\&񬜁U��|��ʹ���[y�ڻ�9��D��r ,�W��x���&���1��٪2� �N$�vL0�D��Ǜ��M�nс�#�d~�Uk��
��P������8���z���P쥯��u�<1$����nE�	�V���CY϶p}��l��h~ ���4���_5�6�X��y�7۾��O��J8/�>��d��������2b��ÚxsM���!�~����ӌ�<G�E� S�<�Ԅyd^�G_
Bl0]0�m�g�^�{鋏��8�'��$�'�`������H�%�^oP�λ�v��}�H�C�J$ C����H�2f:ϲρ�J����L�;S���nM�]Ś�p�:����N�|����m�d����D�mʭ�}��V�\����;�P���1��L97�?�����O�a�,el��	�}�ݭ�C�j�^E�]�r66�{�5����'d�2�m���Ên�؍��-l�o+��U7\�PQw�J������3M��]ջP�cN��$�)��+ �3PM�eB�Y�F�hT"�$�4�~v9{�#\R�u/�Tw����Pu���z��둉{3d �Il_�w�B]m��(��|�@v�b�z� �#a�&�8��1�$s:\���� �9��g���d;�A��YЛ�s��T�����&�Y����=�E%�Sn56د� ;=*�Y�<��F��v.1i�i�Va��v������ȂJ����9�ϰL
!�gE��ް)}ipС�S�_���!���݀'�����j�jա��-�mH�H5`}w'�-�~V�j�����@i��(����ɪ��`���m�������؟��(*~�3�}5�(����j+�KO�^IE๯b��w�{EvW�j
��FLO��q��o����e�e�1L֍={��d�0��Vfo����?�via�Ū��̿��}�}�� �t��zx�1�t��݋����T��!�������$4��km�:zq�z��k�_����D��������V��QK|MJ�jo���\��5;2�N��U*v�X��W�OUll
��,S�:���Ǫ� �ŚN�'��j��N�E30�@���`�Ur6�G(�Kur��~��<2�$�Jn�1�5�)�D^o���m�s��䅍Ub��l���e���P'{!Ez�b��%�>���(q�x�s���w2��<K^���� V2�W�����7�����e��j�Z�&��yQqꐍ^���Y�Ƴ͜k�^��ɛ��dzɔ��\��G �:[4`�p�R1oD��=�f�:K���=�|Yt�D�p(���|��_�Ktca�m��PS�iq~#�խ��L<���qԡ;L��d�'T�}8X����M���y�E�`)%S �R��`�3.�3#���V6A>ũM}��}��ޙ. -ϼQ]��ѹ,g}�@[Z�ٞ���5 ���j4+uL��2�w�$�s�n8�GW@$;���.�i��.	 �=��0��hJ�'-���՛0�cY�]ܨ+z��O�!P˱허�0{%�m����,K۱�[N��3U����\ˠ�#u�S��붖��G4��&�SZn�s}�U�HH���JX����"����Bx�(�/Gh��&�j]`���]"dJ�8�T��R���ci +�0yV������A������T ���a��&^(F��"�?��B��2�
�E~_���,��uu(�D�┻��a�S��7$����4�5Gx"o� �KB�k�N�&s�z/p:���&!c���v����'�,��3��k;�3�w�U_.��h?=���G�{��&�a��AtL+�;�^	Պǭn�e���yŢ�CS��K��H�ⅈF�W\�V��O�1c�N��}�������^�E=
���ޤ8&��UgO���	�1����s�h�Ý)��H���MA6��f���K���bM���@���Z�--G/iI�%R�h��~�6�q��ۇ�]xC�� <�S����<Gtm�ǰn�V*'��J�F�f^v)_��v�i�
 �!��*�x�r)��p���?���[}��j�X��Y���{�s�K�	n0�s����p�a� #�j���-�	���͉׺$M�LR�3>~l�5I��n�<���k�܈���לЧ]jP����(X9a�[����#"Q8��A0�Q?�l�� XԢ�1n��&iJ;a ��єC�!P-A��lI���Ú����&�m�`*_��?Li�$J$FhC�>s���ϰ�����>RWў�a<MK�J��Twz'6~
N+"nӔ�n��ex�����p!��di�Hj���o�Hy;�\�9�Τ81"�1��w��̱��l�c������SKtO��!��h���,\���Ys�O}6�˼�T��5뱩���F@^7`��ޡq�*�lŤ��TVs�s>��0�W�!z�P���G��7X��rz5ߊ�����f�� ^K^Iiq���he{��k��] F�Q	�TV�Q 7'�����aY�����7'b<�Z��~!�>G�'%�t�k���S���,�����UJR!�t8��Kx'��<|$P ������X�2���>���__4�b��B����ٳ�t
�V�~+y��*�����Q#�#/���#A��l̇\�s9|����Z�⊂72ĴF�ɽŁL�����|�s|8r, �t��u	eR����=���{�n���
��'%H� /����2t~DA�|Da\zd�%]��Y�!�S� 0���F�`�߂H���{��3�\�%L=�#�}�;0a�g�x��ֵt�> � 1����]��C.����:�	l�O��u2S���>E%Ạ͕��W��BiNK�
CI�a^�6��V]�b\ݞf��G�V���0*w�����w�T�4���C����e��d�F�u���)NC���.�9	U�,�ڍ���s[D��3���(�^/9@�L#=���#֢��?�n*(�1&�֪��3�j�+fbj��!������σQ<�/o��$D	���
�������LA�p9��M>AV�n���,�6.,;��ٞ��1�!����죨�R���{���綣tz�Eh&1��rB!�3��C�b,�*�c�Bb��(r����r���Ո�g�`��8Ϥ��	Ж:�)G���������A�w�bqDങ��jȧ�z��=��c.��n2��Dk!v?����NNQN��������ԣo���,0?�=�Y� nQ�f����˛���H,c�uo��)
Y��
[0mTt��ru��9��5������Ѐ�壩5 �OK/�[tl��>��ٶ�)�b��*���ȁ��*yo]r�ls)���;�{L\�+�<D3���'�d1���D_�f�q��N���"�|�99��|k��M�GXpF����	�]���	��V�F �O˙����ݪܷ���uc�4��9�B���9_jL���Wd��1���A��58dN'�^|.P�0��O�Bك��Ю�#.B�\��o`�T,�d���C��Tg��>����e����CaT��R�ٍ�q|�ִ%�ۅ�����G�6w��D���O�a@���u0ڤ�]�c+���8�qQ�z�C��r�82ϰ�"��	u8j�5�n�����*&9S"8ʓ9��������4��^�9��zv+� �,��H����h
y�4�K�c��Z�3x�A���2B��&�^z�"�^`tY�t$l�LTi`���xY�|jo�xXZ��V�}9_��
,mG�ˋ�����|�;2�E����pS����Y����ߜ|z�6���͂(�����g�,J����r4хS¼�3�r~���$�*�B&�����8��\JroR�:�") ܬVx���+Nc���Z��>��>Zˬ��� ����
;�2h3"�ߴ����p��8�Y�-�Z-�(e.:�X�!�'�����k?G��V2�o,pu#��(4)��O��1Z�o4/.�$��)��"��B��!	�Y
�C�
o�-L�.0f�,Xi#�˰h۷�B0݅RŔq�;�زf�Bo&�(z�l��ŋ[OX�}a�2�a��6`��W��P^'5���P�L:��"3�ӓ3�rr�/Zl�/Q��K�xC�)0��8z �����>�e��p�Q�sL���Z�Rcx���^�C�����{ҵ�&�7w��:��+Y���@����>O�|��X�}q%)�?��mN61�,:�Ս&�V���2":[�?G�T�[�~��5����Z�2��E���l��I��u�ՔłL�Q7�4��������V�	�����%�~S��;��+.��a�-�;��/��&�J�,9����n����`y�k6�w�ٌ����Z��~��� ,��O
i��������8G�������|k�s�Ա���!cN,ۑJ��khp��=f����OM�}8�]v�W�ɨa6D�g��� nD:?��_6�Dv#W�|�'�>RH�,��g�J�YZ�$7�^�g��1�Y]\�fg�%j����^9|�VD��{�$)�#r�@m�Ԟ/ۤv��1	<�/�1�mi*�K���&�ĕtA���o��^�>��
�-
�4��!Z��<�[$9Ԗ��0�D�_��)sR�U�ת�̆�����#�с��Xqj��/�a5*1�%楥ؗ�W[�J�Q:����[��"@7��ƗD���t�%�R�}wv���6�@_��f��Nn�i�`԰yѬp�����*nno�FG�BF��qp}�������N��[�"�A��!T䍥�Q����^My�(N�ө���IZ9U3�|4n^E8*�g�Gp}�3t�[�j�A28�XT�~cw9 �$�Y�*Ej��Lvm)ZZom��U�A�=���JXW��: R�䰑�-��" �֬fZ:5@zXC�r��O�nC��0���>Y�.�������cS#�^R� H�;���ۓN����g�g�C��"[�4~5Jd$)�A�\%n/�^�ڡ��rw�d7
C?�[� ?͠�+��� �]c�j��P�,�_�i�;&��@Anٳp��JJov��p��oE��{��>�9�X�<��+��z�j)kS[uk+�qvi��<�\k�A;\~��1r��12�b��N
��Y�b��7�+.�ǋ>H=����kSk����su��L'D��� iЗ��Ĭ/��s~�co��gx���x��^�w�=XZ����Y5$>��_v�j�=�YMtx�Ӯ�,����a��^���4H�u��O<���&N��*�)b@z�o�/��d�t�'�y�����}��y0�Y���,�����l(�Ŭ)E�5��Uo?���`�Oa���e*�ϡ�w��q
����C4��a�3��Ikn�v�*y���S��{�6jiY��,�����Xt���O��\l��
�v�l磢��>4kw�����1�ge��8�1/��s�2Ò	�~�@[�'��f*磺�Y�>$O۝�����T$(���_��^y�&I���kt��$�%eK)L�^�[��)���r���sˡz-8�~ �Es� �! C~c��r_�_���v������P�ncTƟV�(���d-̎�bS�	F��&��T	z�aGr�(����@����D�F]�Ѵ�n^��q�MN��=����H���Ei1vB.�N1a�O���UF�٢} o��!A�P.e�5d� �Q��BI=���O��Ǧ��R;j��@����B�l��8ȁ3����>Ď|�*$�����ή�]�P�HD���)��5�J��5Ȉ��M%⢇s����@rs��6���^LT�[�@a�7�'�R'2�{�a���6H:�a.�@Ȧ�&��z���I��c1�:��1n���ø�LC�l�b��`���b��q�H�G����3A�>�Ɗ�Ý/�y���S�XS�|���ϵ7z��������/1���3��ـ�����A'���ƭ��_�
�h��]�΄��c��c���`��ʃ��D�K qwV�FW�e^P`�h�{R�X�hOÃ`���t���$ j��3�1�z		��]��GɝJ�U_�ۡ����q��*���Ya�JM)�@��=�/���"���'�"�4�����~G�`�|�a�j��閯4�	��H�o�T���Z|Q������������:V�X��[!)��{ ���k	z��{�V<��@������}.Sg���R�&/����r�ҿ4�{�@{F��w�!E�0��������ʟM�R)D�я	���[��v"G~�M�_N��мn{4F�x��G�iD����?_��t�g�<��N�&)�·�'��aS�4Hr�H�
�過|���)�#y�A8�<jJan�����8� H���!�VG:��(9ǳ������lU��o>>Nh|5��Fok�N�s?*��>�X�"H�y �ӢV��X�<�ъov���Dm�p�]í��KՃh��ј���v���!V{�/�yI,5h��X�NY�t-�`d�W����D��0|�U"�/�r���F1h��$�_臲���_!`.غF0����@y��X{f��wh>c^�OK���ux�Z��x�Ч�_\�f"�l���ཏ{�Wq8�ڴ�xswJ��a3Vt #��lG�yV�:_����H���"X.g�4�hڲ��!��,�$���.a&?���Hv���%��q��Z�I$!��ǔ��{-��*_�О@d�"��������S��\�^�P�2]0�?����ӄ%�v�]�H�o���<78$��YK�֑�jzr��"��6WHM:�ɫ�}�&���D�_���D��h`�� ��bv�����X1=�!yz�t��3[{x�K�<����}^�ޏ=�=�����H�ʍ��4P�rnҸw&`l�T�O:�J3X�@@�e��u���\0��n*:�懰?8>(�9u�
��ᨏ��������՚3p��=�ի0��� �f�e|U9�ړmP7�q�վgl�� tm\�֍�ϛ�8qq|���8G`ŇN^�*uP� �ا�d�NN�0{��|u���ՐIrS��:>Ug@�?3��|&>;ڠ�d��u�9�<�
$Ѹ�B�(5᠁�|e҈���sB�$8M�'�!ii��	�5�ڕ�x����Bl ��s�X�=���9���9<�3A��k���]��-�\�kO�5$���A���«xCb_����$GZx�#�s��B���>�пϖ�4��'_Z��/����S2�SG��,;�S��C���4(���ޛ�]�oN0�mҀe�)#�U�U�g���Ar>�FA�?���P�����+�R#��[��hnyf�o��XceJ65fi,`w�lc�-}oŭ�蓽 ��<���1!�{ ��S�����}�Fl�
|��Um��9����3v�^)���#��y4���6�
Q7��sk�X��>���=aʙ�P7�{)|~8� ��c3v�)��A*� �T��l^O�1$Z�ὺ��O��rG�
��	;���v�+1�౬LrǑ�h���)��5"����˝�W���t�Y�4Bx�)c����P6u�R~cV��W�?��!���c%H�Mz��i|)z_{�KV��R �P��cH�L,�Ztn�d
�JG��!?/�J���ư2g�=�)��45W9�,��UW�c[
,R�0-dLj�`-Fx!G�lUP��CS�v�-����u�8�n����!o��s9�]�n�.6
A���:\<��Ԕyrr������q�� ��PeqY{o+U`~�bG4�c�����1c��m�S���Vg���׏��ذ)�k�kK��%ǃ�����I�M����4����樔q0�h^�Ny�#��?0�3Q�0��
�O8�%�-�QuA	,���@��	f���}2\�U��(Uz�Z3�5
�0yY���TByL�w��&�-��%oF��U	��z��~9<���?�Rv[u����4N}�hG�[fyTl���h�KF�����8���,�Nb!��j|p.I¥V�ս����
���ȥ��5�dm��p��V���"p}�D=G��|j��7̝���A11�gu��fB��
��4���jh�(Xtd,�#N�C�y��*��V^P_uo6]^]�
�I�����0�֎YuDlPu\�$CUm�����,��B�]iy
����w�?B���BA��R&(�O�I���j`~ML�H���gچ������D��#fnD	4>�d��M�c�Ѣ��#�E/\�J�X�R5����sl��,r�� =����'k�Z#��zO�GP�C:PS�.���?�t�Д�a��Ҭ���' �.�x��>W@�D��a��wp����j�����Y�;w�����8jʬ�T�I��#�x�g%�b�z����0bsQh��� `����U����$_�ఽ��~9�)�%GC��}� 
��u���*�84T�z'�xf��ֻ�PP���e)��5���9O��'�(QR��Z-���B#Y�*~�ļ�Xn949�qv���g��[����F�r�[�ղ;��hp�	!A���~�Dc�mv�<C���A�ͯ�����o��Q#�<����� �.�K�'OxOq��{����<\���2����6�B����;|B������F�J1�T����-��>~�S�#��b�&�V0�����q��Qjn�D����`G$��Qu����+�HK���_|z��x��!��K;FH|qL�m27�^���Ib�kNq��G֥@V��l��t��'}�i�|]��l�,��yx2^�v7��	�I�?bq�xH���m��3�(����4�zS�4��S�]��F���T����`��Hj�������`'xd!S�ݹ�=����R���ڛRM��i %�:&TeT�u� ��Ou��M���D�s}���t���цUk�d�˺�|9�)u�0�[q*��T�C&/�����	N>("���!����W5s�p��"���Y�[oB&�Zb�k#�tn�N Ye�@�v��Fj)���B�E���֕a�:��(�в9X�ȐE	y���o��J �K�s�(��Uh� �ܛ޾.�8�,L�!���bsӗ@ܜ����*���(��8�����	��}�S��<�ö.~o��Z:3��c#;�*��lcWɥf�"'��>����Ci#�j{�CT
8�`c�j���)�lB�#�4��G곎�hfL����U�d�u�'�͈�@A=OY-��o�2�W�$D7-~cUB�	���V���Yn��1�jr-�8K������Nj��9��Q�����B޿�_�;��?���D�F5�� �ŋ��i��xgZ����)�j�'p�
`o �5�ͧ��e�O��?uu��ao|����-^r�ʽ&N�ȗ�Y&i_3F���.��͸��>�Y X?>���o2o%����K�����,{wF���Sj5����4�q����������P��P�՟��w�ЄN
��5:V��5:w���wG�>�Qג � �!�Z�t�?�"B�hWMDA�oF���T�
�9��C���\1��$���`p�՟&z���v-
��� �&t�n�P/��]�t�d{4uѐF��=[<wUə.L��<mo�f��[���B\��O���Jw��|��Z	�b�.x*_�g�\���ZE%Czꧤ�q|�������\O�V)v���I�dX.nc��ZؾJ�އ�!����4��2Gp�N	ȥ�?��eq�-����y8�W�E�x,�-3 �j�T��K��F�������*��jW����ē0�����?�!��U��J�� j�s�!�av9O�f���7�1	٤�3oWg/��!TU�z���]��@N��AN��T��ڱ����Z͌mv�^>*\��=��b��g3O�F�>@aS�@���9΋p�H�X ���Kַ>�n�D?��4�W���t`n��$�P3�Vua�P����L���ኬ0��D\8�H�~C��fI�����z�A�찤�4��@C���NGK�q����-z*�83(��0D���O�r�)�5�Ȯ��+�$=�r��0d*��q��ma��nE+�G��j�1oB����(?�� %dF
�[6�+�P����S|��6����r������g�|�//��~�� �#�� ��L�����K��8F�?�_�u�Ir*�B�#���C�l��>�@"#�d�r�"��VK`xÅr�ڬ�qA�硺���*9�>�MkQ�x��1�sk���e�t�6�Y��*����w]����t���遱_���F�(ӳ=�~6W��Y�F�"]����������*�yR��6)�)^#3�V��0x��)���$�juk�΅�I�E3���>�K�tw}��~	�8��J/���$�ɡW"���x;��I�xn(��cm/v��9h�C%8�w���j\�s��.��X�S�]`���M�9w����#�1��)�HZ�+q��"��j�����!��m��\J?`2z=8^����ʴV=�m�Ⱦ<�z�_���(��p>��LSbt�����`��I����g�Fc�k�G�h�ja�OPs��Qz�$���Z}��xd\�%����r�=1�as���ӈ=�� B���Zo���.���^%kّ[KW��@W*�������T��X�o��"��TV���l��~����b��u�6�*�]�2��ZZpegp��]��"+O�0��<�\��+q�ߥ����rn��ɒ����L�ʮ��?ޭ=W��Q*/%z@���n%��A��6�W����b�De.��!�����/��u^�e�+;r��Y��>�� �*��X��/�S F~��_��|��Z-"Ar���Ur�LJ���y���/{�
��X+�R|S4����u�|�'�C����l�~��2څĨ��Ӟ(WOj?S'�򾂼���Ѫo+�6�����ۺ���H<?�����h��'�`��i��K�2#h?M�d��Q2�t�o��T����$�j�[!/��p���#j�pv���ThoC\k'&?��8Q����1A+&�4�V����,��~���0A������J�S�;?C�/m�
5j����2GM�#�@�o��Ye[#��������/�i����dZpΉ��ʒm)4D��������6�lL��
M�H/]H�~(�n.5ˣ�r����~̓�
��y�Db��Yf�����'��*�c(I<:�U����)��,{�[�W�XH-ؙʻ��fȳ���J�V�'���	����f����l%S��v�*L�H��§ ��j���T!���(�����I/�_JY��dAQLV(�qK�E���LO��q�w��v�H_�;�b�G�=x�9�؛�WaIX#V��� _s�|0��]��OX��ut�"˂3�k��F(��1�6%i_���wpxF�1�}IɼZ���]��
������Ҫ9���EJO�{FH��|����	+�-����d8�U����p5ۅ��9���Sq�� ��M=�k���{�\� �y��r��,�3Ue�y�-n�B.���]t��n�F�Gj�~��|�&4�6U羨4�e�pٍ��R���q,�>R?n�?�/��pN�r,;$�L�ت�N>ebZ=n�'E����uz��_WB��#��:����Į��/ +:�x:����d���P�,� ������a؁Û��h��e���:�������q����l��U���2���J�%�!ND�ι'B����T��}�}_�wJ��v����1M����y��cq�}>1�T���$�=o�N��/���ʳ��@��Az%p¤��KZ����r��H����;�\��ӱ��T�Ckj�t��зD� �[qTTH�bTЎ�O��^>_�f���^�}ٹw�j<7J�BH3l��ͧMoH��������+�"����_�-��2���V���P���Ps�ED�Fz�8 ��o��W�7��!Z͋�� "R@�5,(f3m�X Y���	����	�$�H&�O��Bl��â&����f	b䭇�$�`�Ɗ$�`��b֘��������/b(����`3jn�
�I���,Z1���69�S`v��N5��u��m�|��s���X�Nf��X�W�`���
ס����ib�sZ ��V��P�!�DU`j3�b�U��ߵ]�b�����*���`4|hI/w1�=��D<E���h���}�;O�G����ϴ��&!�rؾM�q}φ��(ċ�M3b���h�Dq_�[�"��앢��y���"VWk]��T7���E6QЁJj&���U��u,fdK�&�-ݢ����>�	�o��w���qr΀��~'��-AHG,��k�yQ�JT�NE�(#��~w�s�)S������v�M�XZTrX�J�-�d͐j-Yv���G�'�{1������Mu�O#�i����{�Y�5�%�ѷ=�V��7uXH�$�Tb��ղ��]xx����p%+e~��rI�SF���G)��*\�9KĤ�6��e�AL������T_���S�'u���g
�E�V�ԆV���B����ν�@\�rrN�h\m��,=�4�q_��s�0/>P�C�Pp⨗w �!QU�������2YB˲G<Zm�7"?���N���_н����,!�}��t�����Q��༹��k�i8���q�?w�^�ˤ���5c ���e��t �0�v�;E%��Q�ǣ}]4������!�E���fڰ�����ry��pm6��H
��q�ZD�^�4_����K�o ��Ѹ:��:5��~�]�H��&/�\
;���Ų
,���o��{�M]��,�۠|�َ�!/d��Z-�!uC�z�<9��|[!X������d%�a����\L:j�N�k�ށt9Qa��[y:m^;���k4�6-3���0J�,�ڄ�9����f���0F����ً��c�9����ж����4N��,����;�t�8��&�.�nZULs�T@9*����H���r-2����q�s��7�[��[�b�f���,͇<�w��8/�c*M��P3[�hXܨ����*���K�q���s�LW� ��K��alډ�gU;rӟ
8�3��d7�
TT�&;`%ք^��X�Th 60]�Vm��|�u��ͰR<=�N17쎭���M�ѹAᰀ�_��,����!�ok������ن��b/0�WN�Ng���=Q0�X���6�|	��!�):m=O3x�<�F]@�ci���iU|�)F�d�<���@�y��-]tja�����!�h�> ���A�A_��H@�?P�ͳ�-R�@��}��8A��ܨ�erWF�=�ֽ����̐b�u�ޮ&Sa�'���HeO��D��z�ށ�F#��1p���C�Ϋ8K?�����N���\,8�MQP/i�-��O�A�6?g�mZ���O��'*�u�#קGe�ͼ�R�MO Չ�*�5ha�u�'���;�:)���M-7��V�4p���l����9�/#ЀZ߿$�CP�t'p�$�1ɣO0%�E�xs�KUP��_��ِ1-GB���1��b��E�p1��n�c�<�Y�:��/ªM�)�@�b�g�{��������LE}x�3��=[��ۮ<�&�7�՛h�^�/�i��lG',���2ʂǻ��z+�{��������lJ��$X�&ݨ�
�yC�\&�����3�^�&w{þ�>Z�m�(ay����,~�-aH�(Т9Q����X�ơ�^yl�5�()gR.�\�v˄��!F*벽(��Q��{a�х�=}{>��6.��P�~0��Ēi����S��c�w�6���>z�AYk���J?�U�6Fؘ�
�T����3��ࣵ��Y�E8!p�g��p�-�G�p$VT�f�]�>�>��+�t�˝�@�.�®��?����9M������eb�J-.x��F��F���UHv�zH���KaiaXU�eo}a3��{����q���7t�S�U��M�݌��Е��0[!j;�<-��.�_P�K��MǏ�|G8��L�㣈'X�������N��>�%�E���Q��J�t$�xN���vĢ�T> ;l�x�7�8pn�|�����K$RQ�@�d<%|c�}L���bUp$u��ɥ�0ʭ��Y�y��G��n��A]&Y���|S�E��@A$�)���tM�9��jg��!2y�����l]7�A`
v_ysQ�/ ��iz>� e�N78�oTkffC�!�3�ڸ�0˪tNhV�м�&64j�p�6\/�m�vx���{eR�T�ζ�������]ɉ���b�{c5�O�i��sV ��C�ʇJ���-�_-/7�U��	[����4:6~J�4X]��i�L7z!n�����Q�x�u�Q����z��Aʴb�C���gi8䟯b#�^�H�1�R֣��D��� (����Y8��F<Km�}���=X��cp��IoV�{ȣq^�z����7�i[����/uP��&E��f�#ڳ���H}�ͦ��������`�RPfXb2G޸ ]TKl��d�Q�O�@�v��ۮ�$sf�a��v��T��XZ�]�#�X�?r�e*�X@\�����Yx$|��Ch�U)�<��ޘ�l�e����֯uCbc܀g��c���*:��t��Z�{C�D����]��=E{>�N��-�Ej)FՐ!W.�g��.]��x�����B�J���ӹ�������� �Y���G�����ũ��<�rT��k�=���l��]�.%�-���;�s�3Kp*Ppl��J�U�Tyǯ�� �󰪼��e�#�'|4��[l��c�bjI��*!R}�gc��x�q�b��1̢"�UҮw�2,�s/����L��u�Yw!��S��
:�[�f0��+�4:���rv��%!둟�7�Ha�p��`��1�~ї^��#�����m�!bF���G��pv'�1�Մ�FS����@���"��k����r��N�#%셇�B<*.�:V��¾�"e1+��zq��Q�ү��k�~��[�6+}�6��e/�����[!���L]-�%��41Vs�����;�l�A<fiCVG�7���&m�Zw�z�l�PQ�#���"/iڍ���*K~(�{�B	/Q���Pi�qZL^X���U��C�~���F���n�B���-�;�#>!����Pk� ���X�S�X�`R7�D�ВMO�ΝtV��AN�32yQB�2ƾ!`ʅBR)�r2k>�t�q$/{JT�/wk�ɬT��z�en�ƲRC�E�[V���nh�i�˅y�U&��2k!���F8�Dk�跙�dx�C�(���qZ�������w�o��0q��i׃BPz��Z0B��,4���W�g{� ����Z���~�k!g���_��K���0 �d*��/�bο	n_��K�W}���b���1} � ���|�bH<[g&����L9���hB��NXނ#�/̼�'`�Ԑ�x5-���5~����i�E߱�"8j��������+�I����G�N4&�@�}@*ܚ\�[���2�fHO^_�e"�H��C��Pn�q�Ʊ��]�aL��	���[`�K��t�ZV�H�q��jȠ*1�DO�ɧ��%���y嚥�Yߍ�+h���[�&��բ��Xu��N5!I=j���d{���٥�P;���$���|��C�feJ��Xo�bv0���4*�1�~Ì"������$6G�n�U� v�1��`0.�������(lf\Kn�V��G��]��/($��w�4�]�ҁG�FV/"�"�?*������ӑ[�K�d�S�{��$!�����B��}�	��%W��w�[�h�ݵ��t�_x���q7BC-�T֠���a��)GVk�ڋ��������ȷ�Üܲ�3��T���mؓ�Y1\Y\�P�;o��	��,-�.ŀ����u��X�hv ��#]<bi�hZ�G���[b���03�ج�������GhB-ՔE���u���R���_O���,;�H�d���D���p0�uo�q��Z^d�;�� �<�c4 �ЬM�v4�y�>%�c�Z��F�VA�'�I�E2�WRpVdI��ꕡ+ f�Ov2|�}�����L賄�||M�
�̀l��~�6�5��~�mC����le��^�T�x
	����mlp��.*�8Ɨ-��hz�-=�֌��ǭ��c�z���*qk��o��]��׉�nݟ��b���,�h_?YNV�X�1�Ԣ�]��El��,�<ַz���Fv�q�����c��0�G����ֺ���@��ab4d5�>�ڝ:W�`ko
(�>Y���:c����.�͟��p f��:=�n��w�H3�����s��7#><�	�\q�#����%�u�D����u��P9��l���}*��y��<>���:}m��#���v�+���mg�X U��K/�_4�$ kʱx�9gdHh��NvgSÿ��ği�l0S&�8g�cT5� �k�ݯ~���]�D�Kd&����r����$����䴖�D$�R�x��'H`F-��������G��%�Ҹ�<AP�3%.=�d4����K���I:!j\{���V�M�#t/O���mhH��q1.�߸�D=�]��7�P�=�����%��y�F(`${)t1'�W_��͊�H�m����7Xq���a�>��VōZ���,��Ĉr�f�B�Փ7.���Dz#,H��Gvvv52Ȭ�f����}6e_�<ps�H�*%�����mQ����̓&D��z���s=�}�pZ�} �{��Y�F1�[�>�Vx���v3�6��J��o�����::��	O�u�����:�D>K -�o1�j[��b!Hv���8��sG##��S=�/���E'#��:Ū�\7B��$���萶��e��ԲZ���8�٩XTj�͐���	�k` ǉР�bF M>�T�rG�8$`�(�`����V,������Q���
�>_�v}���԰Azw�hl𨭔ȍ�i,y<D�m��>��Dx�Ǣ^��������t�*������.-L�Z�T���lW󔨗���y��k�H,T�F���%�4�d��3G�����#����0��k5�9�k�����`c<���3��CVăE u��v{1�X��m_1�i(R�Pui�d8�MKkv�I��Q������C��5�9�X�*w(`B��C�g�v�|x4nk��7|��#u���e]s��ĸ"#WR�,YG��N_(��1r#x#uޅPy}˥�+�4 +>EU_WUw&�Yv�w�X��FRk��8�j�?ϐ���%�k��|���@�|�.�;ţ��b>q���ZӮ[ʜ�e�䮍(0be��ꪴ*�qE�g�I7�?Y���A��
j���
E��nQO^��v%\j��j�C7H�H������A���s<����KN��^�;+���X[��ef!�VvmS@��$�á�7�~����(��N� �Ҿ3~�lY��n�w~���P��L���* ^
����c]b~��x�Б
���p)ԏW�%
G�k�8��$��P?^�]�s�e|sOE���i�W.A4Յ�	��P,�^:��F����%�ml�	���|]��8 M^��E�\����	I�7�����TG���u�̼��-2�
	��6^��	\c\��	���䅑"��V�M��)ZYIO��max4�S��L[%Hе���݈T�����|�K���$���ibv�����it��Ap�`ްa_Z�'�Kg}���R]FCFp~^}��r����77 �g��m{2I^�4r(���Iǧ���Dj�`��`�%�Y��'�-h��;��P]�ixӝ�,q���;)��$c���7%²f�EM��:	#)���)�K��;��iSv��b�X66-�=�v�Z�}A�K���������|R��D�()����v_ծ u�`G��D��?�bTܻ� J�I1�p����`���5���V�)��x�F�3e��@?�3��J[�1D��G�&`���.�	���
���y���`�9뷌��:ßW�́^-�.~�#�����4�"��%�����Y��
>����� \t�S"h�-5���n9�/�~�F����R�}{��aj���O��$�4V��9�����7�E�en���rL{^������p���������@�U��gBȟ':��Nd�?�A��oT���{��<&�ė�ݱ^���{ܧ0�9�M;=Q�C�e`(���M��/� �������*��W?�/Q�
���eT{�A��*B�������QU�eS#c��x�8{��;&��H}���}��e� �[�?t��Ӭ�����/}�+�����9APDHs�؞�|���/l3��[���K2��3V���Z��Δ���v���3~Kp7ʢ���sA�F~I�#��a�Ό�d�Rٻњ3�j$�An�N����G�s@R�ؗ^5���ɯ\	�&����og�н�0�9oz�ɏ��fڳ@��������Xx��.�+���JǐBރ�@��6A��1��i7j�.	D�a56�,�dV����0&%�{M�F�j��_��F�����X�n��2>�GqU���̫���G0���@Ѥ��Te�Î���O����Kp
���(h�W�3���ܰ4
lj����"���'���f�t��t��h��ԑ(yF��Wztzũ]6s#b�ɧ�{�W[HwF�'{��K���f�XΈ�d��-�ۺ��ڴ�����Im�Q�	*���^�l��r���\ �c��|��$�Bi˲��iY�����a�+VR�m>��p\��`������rSu5ņ�`��2�ɳ�Y����P�ʃi�hm�7��R�o���S���ِQ�>\>x�{�*w���������u Ӏ(j����߮0��(�s�P���<�ǀ������s�l�z/;9�4��-8)�S
r������jٳ=�+�ȒՕ������.�wǜ��n���C#�;�%O�X����y��c�IK=;�����ѱ	�?{FS���TP {�Ȥ�
7+��lόe�(���̟WS��%ͫ T;mh2|����1��i[��Q�-�(�ʠ�>E��ZŶ�+Gp�c��Nps�;����o��O�9��0��:�Ϊ"�oZL� ӈdk�ZyM��ܺ�2��~�����͹�1Ԯ�v3-�~��@�ewͷ�
Эƅ�M��)]��/��f�i����mh�g`C ���5�t����ɧP.�w^���b"��G�X���R�X)�?=T|�(`<_U�G������t� N���o�z�m5�;]�-�w����ZeÞ�oʑ�>q��Lo]�3�qb��|�Yc렼�����y���Mh9��Yv����4r�D�:�����RP�C���`���B�k;X��}�[��Hdf�6į:
��o(���k��b�跑���
j��6�3�Qy[�w�h�*?-n ��6Nڿ�fW��8�������[�`/$=����_8�/�^�_%��l�}
��^�8��u��WQk=���YI��*W�u��i��W�+R��Uێ�R�����T�!�n �Y9d&'��˃
m`��g̊���/M�<>���oxmG�VS �l�`�/!3s!e����
� �ل�O�e�$j��xk"�9<���M�������o�Lɝ��[[�[�7=Í7�A�lҤ�t,��Χ�M$�n!�ǥ�%����²#C�gAb�a�����H�[lc۞T����M��a���7��4(��KmOF20�`�fBc<*ZIq�f�L=���>��4f����|�`_��,vՒ|�2�Q\�Q:H��Jb�lm@����K�c#����*D�O��;j/���ʼ�W�dB����Z����}w��I�^mн���X��:��!��.M�����2�F$�����tv���T������4�˲nƶ���CaWI��-�(����ob�ry����$��|�9�5��Q�Y��s�%*?�}�$ ���3ܸ�8���]�e�"�*��������bb��n��@G��(�[S㞅�~b�?Y����N��j~Ƌ��MU_��&��i(r�o��'q��N�[���Aaߣ��{�Iy# C`ބ?OJb��/e�
���9m�e����Q�T�ǐ�y[@]��Y��)i��V�+��
Y3��ě���Ry>�`ݯDʃ��ոj�p�����]�xc. ��v��^���#����)WݺH��%<���߼":��� ���޳��ɰ��ok��'�a�{���UYҴVuǬ��2���n���3��6$�&���%<	�۹>�!�LCm����m�1��b�-�d5����CBV�E#`e����S}��!����G=��o�Z�A݇�4kɚ2����բD�A���ܯf���c6}7�~�d4���1"qO�}���2fBә�O��|TbX��B�}�ĸI. ݞ�����ѽ'�t���e��b��H�a�|zӪ˞��7q�@1
��n��|1���0(S-�7�wZN@h��֥��n�Etۏ��vgZ7��W��r��#.qVܲ+���@g:�p��$0�ƀ�����:�[(V	e�[����_1��2K��iD<�1�9�/o?g�_��㓣�M�7��m��@��"���Id�'��/��dK��x���%�`��ZQ�ݳ;�jro����hK���~�h��J�F�n;E�dL̫�.Փ>`���ا��N�߯�*i�UZ���FbRp���`Q�س�������=ӏ����?�T.u���bDh��RVAb�K��˜�\����u�"�R�))�T��k�\�"�{A}�:x)|���Y��wt+���������>�ǄWM��O��-����j+� ��d�=���j��V��?9? ���Z���F���f���xF�	r+��(7h������jwT��K�8�y�uC�qN|�&٠��,I>��*�T�n/w�ˌ��S��Ǟ��ۮTԭ�1zjFA��=w"�_=C�>L��Wj���������n�����/i� ��P
æ��B��w(��cP��B��Iu_�O�/6�8�Y�!סr�r�sz��OZ���_�^��!�>��jd��qw�Q������x�����o1]=&�71;$Fn/�����ZƸA�4P�ΎT�'��6l����.���jQH�1�|��$�c�HnŤ�զi��3�FM£��Wiؽfq�/��H-%�B��yg�6`����X��mgo�� ��; �Fv�]�4��<b3�ZY����X�E���7�|�R';�7Nd�De��%֜�Uy��t`��$��M�}�[:)Z���EIx'�� t7N��>��������#[���D����{%�lR��u�c��=���\iyc�b�Y���:o�0o��D�i���	q��I���YJ�		5 ��9ym���}JVl�a,���������x�IS��,�Ѳ�]��4����j�o�T�R��$�M\O�}Bc�P�G�4i��g-@����Fǹ��p!Eˑ�X}�mR8V�gLd,+�}X�Q�c1S�'U��_��VG�%�Ȏ.8��H?����
J��~8�G�gR���m#<F�;����9�b#K�t̪��*w�	��<����Ehf��0SG��f��߆T�[��F+��[�۾�X'�Nפ���o�S�~�p��w�^@�@Q�>�%	��p�����
#��D_��^�wu'|��u�!��ν�M��M�><���~0Y�������̈́���X	�����A:R��{8i�jń#�б�m2I����T����d���l6�TcZP���D��/v�/����W�@���|3�����(Q]B#�z�pw{Z?
c�
�嫍%�������WD��o&Zs��AI3��fD�\����z�Sg��]�a�n��iz��u樂�A�|��`�A�R���Y��w
(�O������ͥ�{j(S����(��H���/-�F���Lui�k�����RG�;rOgÎr�N�����.�(X
���~G!�Kg2'�(��~�Z,p4�הZʕa��a��H~�͢"���^���<L�/�O�hyE!*��̼:/Җ����}i�(N\\�Ƌ���&8�-mw��dA����Z���أ���	��ɅXC�o��n޲L푖���A��s	~���/�B�h�sr#~h���4'I��=m~��j�h�%�l�B���~����Um��=ګ�?�����o�VJj+�S��U�Iw�M�P|@��Gv����S�	?_��I��������&�q���.�݅)�����2���)�������J��0����;{�Ma�C�h�|��71��nmP��@�v$C�$zb�9��Q���xJ$��K(���SF4�A���#�L���v�1�(8>Նu�|()�lW(=�8`>�PS[<{� ���'hҤ���
���k���|:���*��vy��NS���m-d&�2�Xb������7wj~�U!+����������c������^|%M1Ot�����Cf�h���_�V� U�2W�ǉ�,`�_�8+t��8]U�5�t��~��&�T� �L�c�����JH�]A�����)����(�9o�r��q��ͺ�ӧ��60��)�:�)DsU�jg:�	�(T��o�\M�R�`n����8�|�al"�5�<Ҡ���Z;�Z���r𥝬�J�fF*Q��J�K�kt�����B�7t��r��ť���Cꃸ	S�|CF��Y��f�-I�7���)<�M���PD�9ﹰJ��J�0=[���hl�$��SuB���˽�EKw��͉��]6�g��� P4'�OPD�FE��b7>��M�h����B˒ф�%�u��F�r��W�����0ܗZV����3)\��n$3p�7o�ЇM�����lNp3��h)��"3�9?C���1�?�@�w�ƑPz�Dr���ǿ+��^���v��'(
�l����~]p��4��<�>��_+��ȣ	[}����ni*�%�X�)�C_�a�PUS S9xNL�i�i��o�˾3��Ѥ�#T�L����1�4{�o������W���|�FesP�(�oq�����cA�0�@J�F@�[ ���Y����D��Ǳ�L��}R$}q��b���&gG�kO��Sd~K�K& h�#%�-V'��>r��<��k���G���`Z�ʾ-M�6>9�KH�8�H?���]~�kfm�Ba�v���?����v�V���~@8ֻm��8��3��#.
���T<����u��������p�g�S!8|y�	�,��g�x��	�S+��?�_�*S�+���C�_�=�/}�q��"�`Yo��O��v;��Z����4"��x�ݑ��bNUBiu"��f�Zl�����(8j�yj�m����d�eN��Ș ���Zyr����8����BO�8��}z��]b��}ul��4�h	Nym��y6�pˀ��qL:Ҁ���~,�O�;�H-��Y��m�y
%�
<Y�T�ֳ�����`ٕo&�{$YsH!��ˏS~�؊p�������%��w`��=�nyh�V��?uo~�U۩�O5{_[K�Y�hI�dL������I�œo�$���h�Ju{ٵ�A&ڻ!�8��11���t�=�!$$(f��Z�ߠ
B�V4Ҍ�rӑ���5g~�y��=�Eu|^���&@�U�S+�@pj��x#�#I���xz�i��=�+�Z���br��	W!�2BD�Oۡ��AH�!]�q�s�P �܍�I�F��4�+pA��@Z���!�*T �)� z{��Id�7so�����2����F�Mwˤ����>�.)bj����ѣ+
���| ,���4�<�:ep�F�Ź��*F�
�*�s���l��!;OE�Ev�ΐ��7��=�`�C�EVPN
I�X�}f����������"�����H��D���d�F&5'��Q��W#�E���@N�%s�c-�K^"�쟬�}�.�L^���&DH���Wĉ(��pq?S1A���T�|5p���2�ϓ�R�9^��M�����L�V�W>�>�G]���	"��*}��^����KB˛ƍ��
�c�� ��K�����/d%�+5��Q�c�
�B�~~7P@���)rbߝ�߾����Z����z�Ϗ��q������d;�˷���$	��|�}�m�>�s�5בȠ�zx/{D�t���}J�m����ⳛ���B���lH��;��(���C���&3�H�5�I�b���̂�SZ�u�T
�BN�Ǘk�?;J�7
�[[�)�'�4�-�l�Z���9@�:�:D��T�m�`]�
O�,".ѐ�ӗ���̆D+�\*��+\���`zV�PT�/��.��:X���~+��q�,���FÍt�v�����iS+��A;�)�Z����>���/OEP�h��=��3�����߸*�<?6<�B���0���(7�'S���B��,"\����$@Q�N2a����&Tћ��I�N��U¿4J#��&B�:�J(X�v/�ʦ��k�Oċ���L4A߮�}r=�C��1��p-IZ�y��ֻ�o��}�zO6{�]"tzNq̃_� d�H�j��6x����A��3�;,)��{Q|������k�!q�qGO
��c�x)~X�����g�h�9����5��/�R��?ʈ�z��++�*���	�-ǿ�{��?�)��X���]qS����`���bu㧚�nlrLLB�N��J켠�N+��en*K/,�l1����:D��sJ����qgK=��}�G���aQ%�HmI5`dT�=X糧�;��-�����$�jz�`_�_�甸��=�ene�@Tlۣ?a����7;������e��to�_�`4��,�|cC;h��U���

c	����@���|��&��p+4< ���(��gA��d%������X4��qJ�D�k ��OBuWצͮ�Y�.�������)�Y�`/�
Uރ����W��K���El�_���fQo��eɆ�e��fy�,C�e�^��z 6?���l)��Q|I�F@[]FJ]�>��X�pc�s���}EAI���9G�:�*��-#���Ԣ���������5�:g���J]3X�KP0O��^䝨���푒G�!$�6p��iW��⟒}�p����aL�s'������{�ⅇ� �X2�@Sz�])�+�����'���o!��<|��A�*nĶ�>x9A�B�\gǤ:�N�Lv���&8qU?�n�����~�4��x�Ԑ`����\:�N.7Va�d����@\-��2���.�A�oEw.D��.�}�/l]��#�\Q��B�y6!�����6�K摊^z�;�b}]��n�D]	r��F.�ӓ��C��R�POӜ��B��Չ�4݆.��,�'�w�j�EK?
l;�☟a�~m��2<�wB�Ψ��<4M�q���Q-�u�#�����G��0p}�|L��j�jkAҙ#>�H�6\ރm+Z��+����>҈�lE5(� ��L��?��}�'Ќ/��KyP�ɮ�5�[A��&e�b�ӽ�c(�J�_�Vܲ)I�����Ѹ��"�E*��"�^��Z�gLhR��z)nEe�.i%i���&��֥BR|��,���	{�`\k�P����ᥔ|0s��r����u[�Oz�"�����%��Ц����	Bc�a�Ӕ��pe\��'�K|�i���1	�d��Bm�,P�,�9�PW.�'�R�m���^��_&�ntȎ]`��N�	o�:���偕0tQ�qK��݀!&b�>����/�C�O�B��Z��sۙ]�+���¾w��]��^�ER�Yb%�KϹ8=�m"A̧�;Rce�>L��!I����8� Z��C��N���_�ƞFv�G9�>�:vL�j��#��T�B��k�H<�[n�;IP�6B�d��C�I_��Dȯ1)��U�.$���'`�(�>7�c�Q~��r��yl��˧��g-{�IVK�h���OU���.4�OѬij5CY���'�p2�5Ұ��)���>�ӗٓ��ki"��P�^A���~��iЫ�6ϸ�g�"���y��A�����zW��Gw�WQ51�O�H�k�uMxIOߵ^�"6�����1ɭ�X�K7�3�n���g�;�W�������T���J�Џ1�,U:�����Q��ڜ[��;<������fR7oqj{x�U��6�=Y?|E ܎�����#G���יy��h{��i# C������FC��nTܽh뻾i��1Z��Zg�J?M��ue�iH)k'pR���}z�4��TG�t���Pw�����[W>O���@��N]��'��n��l�K�G�l[�֭*��p�9�D<��?�7vS��eXQ~�z �����Q��(���O���|�Ϩ�B$N<�$�~ ��y��0ք[�G�1pC�FAWf�:(�eƉ�)_g�W��:�M�W��8˶5�\�����hZ��\�gG�[��Y�3�F�Iò����	��D?1�)b=�L�q���'�]5��+v�i2N�����i3�e������[E�0j�� ��&"=FT�P)��lB�|
*�KН¥�9�h�/јx��Qukֺc1wS@5��R=q��Q7ud�R��u������{b#��huKXdf��t������%��
�Q���JP����L�}�MҨ�@K0�`�@�9�:����$Y˅��w�$�e�[�g���O�������$pX4n�B����zU���%;n��~�)�5����F�������D=�9bQ\�P�n�e1�aB���,�[���ċ͵z����C�^|�ٱ)�4 !Z�:�3��л+�"���{($�ˠ7+�ǥ��X�듲��e���qM�������u�Q`�:[FfI���m��o7!�c��`?b5~�Ε�Y	�Hx�؝�#�	Xk�P���)�Ph1��$�|��\$�.r
H�K�T�>���D�jԈ�@�
��D��R9��5fM�Q��L��T���Z��Rq5[J�:Y#�!I����@����@�.;�!sD��I=���%uzM���S�>�\9��O��e��@/�f��>P@�,�K��:i���/ � VL���N�4͑\ѳ�����&���5�|T�gr��*����uf|�r'���h��b~��z��J�����y`q���Q�H&Ó#��j�
5��l���۝�򈥇p��B�K�7)��M����e1����΅�@5��'ú�f����Ug�T�ɜf���䙩cnSF���xCQL��Z�!�nr�/D#�"�/�01s$��(=>Qԅ��t�~@W��S}ϭ�"U�l�fkr�Nݕ��Sȫ#~�a�T��a�<(1
!����!��aܙ�dRNR���A�q�9�IfDc<�~�u�-t-�˒``)�5��T�EԐФ`��!�T���Q�M�^Q����*G��}�����n�	�\���1
>� ]��:�v�YcY�(�����;N�x��g��%�:��(!�M��j�����~.䥎�:N#R욷O��Elq��k�"���[���T�U��:6�M�3���(a�A�`�e����M8aB3�qR&Q8m�K�i�乒�jR�(�X�\L��ٺ��S!d��_4^y�L7u}A�t[�0|��qb��~BB.	��}�[)�6�K�T��!G���`��-:���y�Y�O�^&=�r��J^���6�v�Ռ$�� �M%h��Z�dOF�w&w6��Z,�3<O��v�+dF�iן�s5gyHv�|0�, [�è�jP��K�-��d���h�c ��(.\��׹���a��2�+�F?�.�p!�7���i@"}��}=^��0e��)1���
H��wQ2��^VC����(�M�L��� ���Db��ˇ�0#��o�{�~E�_�mľ�khO>��*�3�O�Nmac�u�A���%;��l�:�`7��CӪ2'�v�d�$&O��2;�TC>F�c̈����f����$
X��"��F�q1싂w��p���d ���#(�7��r��rE��f�ۚ�)�L:]��͖<�ݦ�����D�_U˽�/$�f1�I��;ʇ��[vl�����u�=��g�I�#��s� �N,%
�x^�DC�o�=�.�Y�#����ޝ1�S>��n��§�u�}����c���b܍��7���v���a�{�ⱏm���.��VQ�Ϗ��e��"z��8 JR��~�����3,U���@�e� ���
0i��<%�Ƙ�����ت�S��aR���S�u�}H��Μ�)
1B_�'��L��b�M��o�hQ"B�a��CUb�X<m�W���S~�ҬP�LmABb�����(�M���47⥢w��ɀ0#@c��Q��M8>��W�f���٢����}�P7�0m�F(	Ky?�����R1�XZ~<Cv!s�0�5N�Y^u{k����$�i� y�8��)�A`Qci�f�9n��9V-���7j+���RĒ���4Le��2Jlu0�NF
1��B��Ű�:��!��r8�FR�X/B*�A�v.!��7,�Lh�۱�G�D�)�����j۪�`���R��`f�,=^��an� ���	�l������[=X&?t�����]��m\	M�����7"�q���?`��!Co�3�o] ?���<�)JF�y�Z����k�Z��5B���@����(�'s.=ɐM3&��%�a�of��R����#���ﺲ]��{I�2�f:\�96ۜu����� �WS��E}�r��<^=�=�T�� ��(ṬO��ٔ�����f���~�m;�$�{98�ｻ����G���i?'�����غ�fX`�>�6l.Z.� ��Į�̌'%������,�n�reT$��k$���[�)���Z�ʣq��7�ω%ᢕr�1�@Ua說ӕ^��W:2���|b�^��O)~c�;(R?�WZ;�
�Gҕ�+[0��Y�L.~�o���y2A?42)	>��?���=����vSgdƒ�O_�f0��o��˰t*m�@��5M��U}i��r�ВZ�7�S3�c���䯖e���H��v4V�
�Lf��@����i����P���sO��q��[��8��[)׮Ε�?�,���Q׎���^��o0�y�4Ȃ?yV�&�v߳e�Дr��Z�h0�SY�-:$TX�b?stgW]GW��U���&�HRJ4E$�ZP�b�����ݡUߘ�vMa�/N��3u���::Z+�KA��|��T:m"�y2Z�#�l��p�{�E�ც]:�jI�_�� ���U�Ow��oC�6A|���{S/��{� �z�v�R��o]���x��M1ˠ�����_����X�t�^q�����{g"��L�]`��P�CQ����Y��#d8Ѧh�/��0�"����{Ah�0��o�wD����cۅ1�i 0+������M����{4^��?��
q��1,ӻ�P` ��+oLQ	p'����w!�ZO,<R����]�=�G�S��^A%�D��q�p�Do�Ƈ-n��c�>�HFtp�⨲��b�¾��}�F�2C��*����O�����(����ֶ!`����aY
�[���[���AO��"�	�(ޮ�
hu|�ԓƭ���x�D��W)X=���Խ�©����@z��^� ��R1ܻUNwv�`T�c��^���w̝  �d�V$���_U�� ����b�Fw~PQz�������b���1=w����9|����q��z��������=7�ǐ��7���&8橎?�|���)<ƈo��Z�r�]�O�K%�h���Te���U9d���-�!��bd%�U�\p�������(�f�"4�+hRߩ���B��̒���=�Dt�K��4V1q��.���*�_a� ��)G�)����Y�Pd
�{�c�ُ�f����/(�:��Z���)�����Y�L��@w�P�~"u}�m��^�p�FP5�����b��)�N��fI�y��iZ\�z�A�_�dV�`���i��]���s�s�8S%pT\��\�|�����5�p�����Z�d�o��O����BeӮ݂���@ВA97�د`y�Z]SE�d9�ή��l*�<���g��V؄�3�`Ｑ�s� ��Na��r��!�{��UΙܵu��T\��-�#���1��4�I��/Oc�}g�vz]9����s���ɪ�qm��E�f׋?GQ�3W���n5tr�����ص0j-�
g� ��ZT L,ǫ2�sB4�Ff͉|��	!��J%=n6*�`�N��Dj�SUg�"�����o<�l�<f"����͸�F7���.���i�j�l�v�m�Z����(=/ӴMZ�GQ�*(��۝�/�%t� EJP�O4�}��@�,C)+=��U3���xy( ��|(J�!7����I���Q"�sR1;�c3�{ y����ف��Ur�b��E%�n!Mr
��O�����w�׌0�\�J���=�A:�ח�a,��K�O�)E����r$
�!R��+�M��T���VBm!�5	���;��r�V�ۆ%�Ŷ�	FPD��O)��	'uJK��Ȓ^h�]f�~�f|���a�Kt:�� �
d�a�F�'B����S�\��<'.�1�䳬Bmb6Z�(Z �0Z����39�M�z��#"o���X�߅h��$��\2Y����S���N�;ki3�����K�a��y��4#�{ᭌkȤZw�J�A�Խ��nU�I�Z!~`�}�TO�?z�d�G>}�6�S��h�VS1��:F?���2�2:�&��jA쁱�<�uD��
��ߡ��`�(˻m�Q��X���'�|C�{��8�&9�&�@j|ֵ����n% Y�oC �J�$~X�}�BG?a"]B	,S�T�^ ��ʂ�y�� V+R�%b��:�τ0V�"�e'@Mc���gWd��y��9���ڤ�+N#�X�ʮ��=�8s9��:]n���%��ڵ��ݯ�Y���g`����e�*#J��HW%�{y�J��4�Č��e��@�x������-��d��Y�|2�V�Z�)�\ R��]Ieo��H;;���au�KEBX���Bu��������n	!!�)[���F���`d'��h�;�Ɓ����A�'~����*;\�ʷ����¾��Co�Yzy�c�I�gLeF�tǭ�{bϾ��r�J�k
;#:��H�d�5@乛������|�R��׵pJ�j���Z�]��?ɪ;#Τv'e���d�h�;�7��if��b;R�Ğjn���#]����zV�0kcf�ˣs��Z}3."�<������1��**�Qߡ!�EO��:�{� %`:#3S�r�Z�R���d=(sX�/�ʐiu#$B���*�O��M�c�#	�FW[|ey�n)��>�3nO�zo��^K9���MZ4<r� mO�=鸹N�D�+tQ1Z�v�
��7�c_������%7Ib���=��:fQI��X�Z9#�|�	���;Z�S7���o�{�?�b��?�x����q������t
�\�ƚ��F�����<�s6���2R޿������'c�(�}���&ru	�m��⠑Y�xK�V񧒗^�f�!�Q;��0��V>��
l��S�Z�,�=���C��h�*�w���+#��+�r9i9������ +s�w��m���?�=�% � ũ#{�`$Wݮ��S�4\��������<כ��ڙ�Xe�=
*M�u1<i1Ȳx$&�O�N�W���(�H%��=SZ@^�c��L�"H��=x] �ʭ����l�&�y�]:��]���R=�R$�̕���C��L��+�龍�N�Z�)a2��Q�[$^����Q�mnCq� N�f���/�t����s*�E�7�W;�<x�[/X�`�H� <+H0?��3�2>׏v�0�/��v���#������u�y1���J�r�c�)�X�nɭ�)���q x��x۔҅���
�����ɵWz߫9��+�Ā�i����8�ݛ��@(�<�Ӧ�5$��UҒO�(�:3������Q���Q�5"��)�n���&��j����4�>F����b�WZ{�j���mj.Գ
��N{s�oY�Ю��!�YE}뾫�-����8d����w)>�C�ě�=!�(J��,�A�}��4��(k�A�ߧNO���i�@ѩt�o���/l���|�-���/�����yBT����"`*��h����e��T|��I���bU���	E���x��z�}M�1��xd|	8��칼s�v #�{�Сx�ȳ����+L���{VWx�%v
� ����װ\���a�����-"�u��y[֜ǓK@H���D9��cJ���U�E���B���f�u���}p�����\��4��i�	Ϲ���"�S	||t�x'8��UCUQ�r�.m�Q��A���0+�6����8���@E,׼E%	��۽�?d�����y6F�a����w�Ԣ�sŖt[B���<�{@������
)��`���@����ݢo�EϦ�VV����M��Ǖ��]Wl4�q����g�����;�*��#�̒h.����ō�=��6�n�w������
����Zk�j�H���{��?e����VK����q0��Į�b�z��-"_��EW4��ܕ2�5q,����A�ģ���xYU����5[�;Qε�N�9]&�H#�Kgw<M5����g#�5xX�s�P���|Ri��R��N{y?H�ђX+잔�a��Hܳ���<2��)_�7����SO	���{����J�rj�X���!R�8��V����iu�Z�G鰙���������p,񂀸�/=����J��9�:~�RBΧ�E��.�1m��f|l9)�ɴ�V���:��~?~�Hg.��)�j�Q�"���#GWEZ�/d?0�^�� 9�8� I��A�en-�y(6��~JJ9����y�F�x�삧�O��{�a���,�%j8r�����Y�b2�ë��#V�5�{>�5�)��:�� ǋM:�kp���6���R��R���H�׭��^�a���̭����%�����T�Ρ���P�(Bg�M>��@d@���B Ѱ�sv4��A���H��В9%�DRS-�
�پb-��RkR�\����B*��_�D<4����D��I�V�49�}����ho�m�4�BN㲯��;*?�t�j�*��j��W�~8ݓW2�̏�kt>��lW�l͌i�hhJ�O��58�|lD}n ���Y�B��J�S�=ɘ��q��%��c#Z{�����C^g�E��Tu�cZ�b�_�'�;u�U����,�uO�V7��T
�����W9Z�ŧ�z�l=��B�_
��oS����q���>'H8�~�"_�؁ː ��K�͛��ӳ(S�"�3'��2/���@��X!�)\�*��i�!�y��ϐ�Y�B�j�:bf�Dkoz��A���C,!�ޱW���f����u�c��a�D�E�`"��8vt(وj���`;�=6�ǖ>�*LD*.?_�ߧ2(�x3�ߠ�Iǃ��bw<�+�G�f*C�.C�C�ߡ�e�!�Jd� �y�(�Tӧ�L[:���	�ԃc&֓���m���-3�~8pƞ^��{�W�4���7�Աe]��ݬ��O�M����M�ŨL�YdK�\� ������5��n*��Z ���:��!s5��`�1b�U~[y��6cPu�N�G���Z���0@l�����a=H�H�O���*����X� ����כ{i!3��3����'"��t�k1��y�;h��˯ԃ�l���lH���F�-2q�*���PgYd�3=�Lmv���U)�q��_���=0�N���l�|��u44i����)��x��N\]ۼ�f/��Ȳ����h슮}(Ñ�RhD��j��S���-�]>W��&G �jj�r���3M3q�����F-_���,kMR��=�M^u��k+×%_�o#���Dy�N�/���`��L���zت������������   (��w1��3��e؆M���8U>�|�֏?IU41�z
%6u���R�`jrR�(���[e�����y��K��x�c�Eo]4A�c.6D�[��Gl����k�g��NUڽƞ���՛.
�l��SH�>�&NL�g,� �^���$��BSr���Z�}��'���a��92d\q�_-l���j�����η	��F'	gP�՟��O`�$��KG�����0�t�["�94*.sIE�?���{���g���_�闰�4����i۰A����U����NA��܌��D��{]$��j)#G�T�Q*�7��׶6D�[�E,	n�K԰S�e&�����TY�w?C`Уe�[z%�.]J���GA��I�8#m���;�.aN��P���W�L1g/ư��+�Rr�1��X85n9�y���	%�%n�S���)�Mk�2�vJZ�}�᧾����Ը�X���_�غz0�%��]�v�E%?�{3���K>�j�oǸ��g)@<��K}������Pr,ՂgJ�en_$������٥�UFm5uJ��ˡ|�ʖ���4o�h��ad:%!_�	�$Ò���.���I�A˻;c�t>�����i[˹=�F^�4ޜ `�pz��Bn�+�4��-�[1J�3ǅ~ct;x<�����|�s�պ�V���uu�ED!W���(
+�-;��a���NHB; %̖X�7��M�}y��p�q�($�j�W�F�D#P�*�Tʰj��8�Y��E���Q.�\da�pWH��N	��H�w��g�ట�!�%��!����Ib�� �[�Ϩ��Sۛ�$l�cU��-�Q=�w�5�����{�:p�]���?|8���+�n���K�\�����I}y\����B�yt_�r����slw��<1'����8'��i�f�k��7h��bN��HJD� Bw�P�1���Knyݫ&�'�q��۸Z s�m�Eߙ�r�sv���������T�!�Ӿ�̼�Px�"Z*��L��2�I��l��]��~ _�
O����>r2Ң���� ���8�������ҝ���N�����ԍj���"��g
r�����)��!_m�-Y:kWNE��ts�:7A����r���� J��'��餑��Kt,��M��CҠ�
���9���%�fXlhԏ��h.�sYr�����.����qj;���~"�|>3=��c�h;	�eC�"�����Bx�.��Ja"�Ӝj���j��ˎF�rX|ϟO}�x��s�Yt�G^D}9??��,4��o���N���u�Mke�OƯ>Ʀpo�#+�^��lչl�ׂ+�5��_�B��5c��Q�8����7�~h��l���4n� ��&X���H �&�Ff�=��N�!� ��mx��߱}5	�d��S�
(ZH�ȼS����Nr+��t;�򄴵���4ɶ�|j�hv��A![�=���eAZp��>�j�V��ܩ&6%`�N��T���W/�2�?����P�(�%oF�6������	�'�h;gg������I�WJ�|A�@Rӣ��=G@3h��I�ҟ;y�2袛*5c�w���o�E�뢮�[u^�${��[!?��*��i-;KI�q�O�u���H�mA�m^X�Ƭ���1@(��_��&�R���wH�x��4�N?�U��B�$=�H[�8�A�"��W�r���ށ�#'VH��]�+�,4�������Q�ِ��J��Hf�ԩ���c�|س^M��D����E��i.��:�l����H�j�<K��Y��+�*[*"�񎵿J��@�4��n}:���4q�u����αjZ���816�w��?Dj7��o��[��b\�o
�A�M�d�-�!T9.��@�f�;�An'��dN��G]I�s�M�p����(�u.ɮ�4Q�8�v�p�):j 
O&��J{d��zaa\Ư>�*�J��K���IR�V.�`TQ�y�(���_��IQ�œ��[��*m7+}��A�5�嶐l;L�����MX-Zg��LB�>�j�B#��kL3E��wk���1�!�x��0~��7�����(s�#y��F�䞗3�[�Ď��K�X���B�!��a�!t�X$e�N�*5Lu!��M5��+U�`��{��7��*�\�ػ�e����f�vE���jʸ�S�9Y��/��1�I/�mK�Ƀ���D7w��0PS5?����o��T2�Q�iN�������"�=#��칹̓	��zL��MOO5���SGO�3�����{�Me|����
,oA��t���*2k����-h��}���K�fM������s�7̲��P_�\KKO�.
穖��"�<]�pɯԉ����mi�&���]M�����^��K�m�������m��qdH��Pe_u�-�����w��1��m�]�Xb6=��s�����ΎM��u�3�äNH��Ob�b;OR�4G���;I��H���^�WN�m��E�H�V����^x�%�}���km�2�qGF���6R����z[�)���6�P��x��v���f��%�~�h�zL�b14���qr�����c��h�� �tL��t�V�B\���ر�j�%�!�?��翮��M�W bv�
�V��b��\��]}ݸ���2H�+A������S?a jwx�~䕂)>��O����������.��j�,�<\1�-�x7	�	�?8�K�6��(�2\(\�%�OR�vBv��~�7O���Mt�Ԙ�X>��yˣ�"�4�h4���&9tV�{|�> �KQG�vx�NqvÁ :��tw`'�aڕ�"@ia�vd��1�dr����mH�&h� e��|���}�ʰ�̓OeoEI��}lt��1(g���v��Q�-Y#��i�[�іO�5�K�A����㌉�L!�ku�yx�̓R4�qYL����|C\
<$Sӓ�)�)��L�= �Y�	�%����,�,?�ȶ{���egˠ�l�&!mN�Vq���֧�i�F�o�	�M�J���gILKo�.l���}ۣ�0Aէ�Rۥ�����dI5���T�-�Ⱦ��H���A.)�o��L=��2�����؋d��Ύ<N��α�oC]�v���gv@O��w	�����%Z>>�=��IF6�����<��B��dՋ�,��{������nC���с�<WV&�z��'s��hp�������8eCd�Q�c`gu%�5Ui+�����H�Jb��Mv��H�04=�5���nf�d�h�B�]0v���%Ƕ̴����K:�%s\8#����2�4nӟ<6�q�!�\�XOZ^�DzU�2$˽��$�(�Tox�V�X�Co79?�ì3��q/�TG�\t���ndBB\=I���&�bj����P���:�I�<��?�}�!��}�9�}��1�џ��9W�	X}�I�/�I�(v<X����u}���?qD� ��4Y$��H��hA#��fB�\�+�/�q�or_������JP��u��q�1�Fn��9��<t�Gw����� A?�~���%����d�mn �{_��CU9ɩ��3�d���]k�Hįeָ'š��l@���'r��.�lH�=�~ց�KԴL��&V��B��� ��.�n���7r'���2�*�͠*������v=@Li��6�K���p?�M�>�T���ENV��5M$@�HI���n�g�Y�M1 o��%���c���H+2�I��j��]I8��D^��5����Kаr��wLKU��o�ϸm��SxV�}���/�[�p�Vr�H-��Փ_�0WBo*#'E��8�{؈��	��_H�p#�<�|+���5���z�\��|
�>N����q��䆗x�L>�x��_�Kg.�<�5���\��3����z�5N�uLV��}���5~�[�|��1�ܐ��(f��^t��AD��0�
��{��^H��y��L���� �ᜅaS)�t�T�����X��HZ��~����O��#Ț�ǥ�i���R�Q�s��u��A��ò2~���l�H�8����z+��U�����Ʈȥ�����7E����
X1���Ѥ�a���u?d�V/6��W��*�/69P�o��%`�'G,��0:R�鷚{&H���c�H�eL���.��[95�L��j'-h�m�p�4γ�����k!�'!���\B��c�����E�v�	�X䕋(Ζ���j/���ۏ��,m!�iI����x���-V��`���>�����n���G��i?U�� y�J7F�P�2��Z�ޅe�s4i��h�n�j�A�Q�2*Aϼ���!?��n{/��1����!6�{ԈR	ݸW�v��$M�N��
/$�7'�+�Qt����{��� ��9�=c���0Ʋ3?ZI���[άT��<��
Q����F�Wѱs%w=�9���\��j;ٰ_��m�p�~h*w��j��?��M�j��7�����R�t�R�9��"�(t�TGX�<Y�	�y3���o�EL�����u$8Ay&����_�z�x��c��=-_r���ŉ��zd�l9��i�;/���.h���3� �ϵ��-����b�?d��@>E&�z�A,!,]��r�uc날	�1.-õt�cs�%��%c1��ihRe��u���΀��G��y���t���9[����B��A�C��ڳM��Wx�����B"k0AI�@���%�it�YUI��	<	����K:S�x��Pl��Y`��ӧ�S0�o��W?�c���)�WP�ǜ܎u�Џ����'h��2�8����HczQ`��=n�)�*�\61��R��]m5��F��O**���)�S��`��x��C��N�}s�L@���{�8���m�*��e'�w�a�:�����`��B�m���A��zI(�S�*#�Cz�s s-)P��t7)�� �������[���wVW	?�n�c�/y�nL���[���iG��/�L��z
E��̖�����
�h[���%�� ?��ur"����=��̶sk�U*�1w]�/��Q|;ܤ%R8�b�C���hh���3voa��Dԟ������Wg4S���Rg��O�վ�ưp@��	�|����һ�Q̰��5��r�;�1Jqj���e:b��"��~yHM	���X��P+j?����������a�I�;i�Wje�;>z�]��M�0�6����a)$�+���X�3
H>�'��_�d��[L�k6��5�/p�- �ZX��=t��Rq{u��`m�P'������Ƙp��J���yM�� ���^w7
�\P-��8��ސ~�?T�m�Y�)�Qm&�����w`�-�����9�����B[����#����Bi\�C����p�-&^f|�#r5��]��_{腀;[�vV]{n�Mo�4�U�G����<���?H�P�7�6&�J��,��(��M=$cm7z�ѷg�.��������I�7-�!�O�ʍ8^5�uW�e��f���仝Tx�����;�A��QɋJr�+��\��w<�}�9�H�C��٭��6=n�d
A�
���9�C�i7��nD��ShMy�e��}��&P�\�h>����i�~n��qBy@�Ƀ7��ta�&|^Q��្��κ��'^T.��<�b��O+1o�/ ��=:A�	^6$z��'&�1�~��	�0`��7Ϋ��� �f�f���&�I�~�y�qdޏQMv����u���T��'�	 �
6�e|�Sh����$v_���-�{ �7p��Vq��t[��@2�מ��*|��<���x��X��`�ѵs/�鎞�IZL
��Lg�Z�:	��*�9õ99"�wL5�!��%W��*���9n*_��~��K�73�/1-X�h�P�U��+�_��^Jm�!�{�����p����b��[�c�>�`MD��6��V#�!IBzf�^e%�nk�0@�8%�k�#���E�����KK����xZ̹!�x��%��gϠ#���ص"�}���-���W���3y�X�c�s
Q�E<S��S	�l� �G�bOl�" �ŋ��}0�ϼ������~t���A�#����t�[���;�!b�a�:��Ԓ��a�d����Q;4����[�6I�	i��1�ٹ����2�44q;{[�Hlۖ�/M^�.�{[+�_*����1W�V 4�	8=W��	�l��v-���,vo�2fЌ�`!9#ؕ��녑�����9]�(e���F|T$��Б�IV��Y��w���M,Xs�T��Cc���I0��� �pZ�x֐�W�ٕ�%����ce�%o!�1�B�~OgpZTG�M�7��j�nz<=S�;/C�rG��g	@�v)���t��Dtz��8Λ�^���R��M��������(�J�{���_*��)��e�ư�$��V�t �V�^E��W5�B�6P"aU`)^|��:D�'�X���
�=�g��Zc|WC�f�!}҉+�8q���;}������)�ww$����4��M3'����h��|�|�NQ&�g��}H����̮l4���)>.���kj�ɷ"��(+�2�v�ʚ�q��w$�aSc�$De��P5������Y�)g$��H��=�{�y�=����t�
6Љ}��H��xo�)1�SR'twh�k5Ml�]��'j`$�Y���?��p�w��u%������Ֆ�'�{H��H\5_y��Sީ��CwÞ꫎�`��B�|�X��y寬���8o)ݟ�&����2��T:����S�����x���t�( c?�z����V����F��8;�����6b�aPJ=���տF"�@��s�$�f9��#xfh���` �M1�;�i�h�p���7����t����I�I+�\%�y2���[.���+J,���L9��Aʊ��8�ojz;o�mF�
�y��zK���;������Bcٸ�e�P�V�uR�t5jz[��,��HN�=���}g+��!h$�p 
��E�Pn�&Jʚ8�Xx!��f�6���mP�^�]e�Ҋ� �'S�~
�N��WpC�k./�|��v�� obʫA����v�'um���AA�؊����Dz{}Ը֦�)�,��������Qvn5�+��I���ܛ��� �*D�o/>Yŧ�Z�T��֥�*�#u�}��qN�"��k���I��o���P�%�fnh���f(#I��TZ��6sh��s18�=J�@�6N��&p��75�	LֹIr�P�Ϡ���5]�V������������������>�c*���#Ҽ��������@�֞�Lx2��s2���a#|4�����%l0\�d'��K���5�>?�V��t���|�P���m�}�}Y����gPx��&I�1<WH�S��:(�@�6Ym��V���j�J�差��ޝ~��'�n	*S�J�=�PE��33rI>����*b�\p�D�I2.�o�)���a r�W�O��(�zC�_K�J�I��}��s��Nn�o���^!�s���� ~�Ra���)˃o������=�~�Mz�)�ɯ�_0�p�ת0Y�����/4Fo��H,��x��|�$ń��Ŗ��z���ͱ���|X&���9$R�b��G�?�k�8����������<�G��m�5���M}F�.C�9�%~8��%�����j*c~��ܑhBd��6����~�M�m����|R�+��:�C�j�?����y��}��o��hj�N��!� �i������Ț�����ƕ��}�w=��I7A��F(uBQ���:�FZ4x��\Z*�F$��!�iH�\'���m����2D�z���d&������.?6�+J�H`�p[��Ξ1�,
:)���f��E��&fo�`�c<i%ⲷ�+��·i����'<7����Λ� �3x��wż-g�4��SZ�F�!uһ���M/$#�rwN��|,� 槩�(n@76���Si1S.��s�c���,�k7�=9�J���s�ݴ���ng���0��Ct(v�zY��D�PΔ��0Wn�Z���6�(��w`G�������戃&ź��U���~��|_�~@�}	��~{؉��~�ʅ�xUt��6��#�F�~*���l���z)��#}&'[� ؀XAP���	\�q���Oi�=���Ί.Vi���7�-w>/��Et�9 ���B�����Ր�j�7D�v��M�Y�/`�"�j0�n@w�y� �V��N��&���Ys��< ��������ټ�ڃ(�V_mɜD(��H� *��+�/�T��Є$]�U���]*���4iF����ˎա�xu��Cd�Ω�^���Ƿ:U��7�vZ�@TD4b<��Рʼ��KP2�7���k"��h��:���������z�d+�*�s0�CQ4%<L���ꐜ��)�0�:<B��5,�a���v�-��<0�� wS�SG���-���#��ʭ�T)�>%�W$H�KUo���[���pwL�I���=��4��⛜	EDԎ���2����ϩy9e`��S�Rl<!���?*���[��ld��%�H�>���9J6�����Fa���`!z�ƃWU�\����z��$Ǯ܍�ڸc��L���DS��V0+ub�@�� N�"tr�n �!K�q�<&��Bm�E.�ih�sB]W,���[W�tP��HHÍ~�"���˧6)�J���B�� �w�� �����4@�4w���B�'�eE�*QU�HmgZkN+�H��!����9��TI[Cn�!�j�H8��?���Ϯĳ�EV�P;�r�(N!����-S8�●� ����G�a�rtZF�ѡ�G��Lv6۽�Sb� ��C��'��X��JI��~u͙\~�W���w��7���X�y�yտ��$2�t�9eR�W�m%�`�U^�s���I1ȟ2���f�hmn����Y+k0���/�/�SQS�a�{���V>m9�#�+��]vP?�mL�j	��v���E*U�a�y�2�'�w�8KƂ����خs�w�k �Y�s,˪4�Ѥ����沍-©Ň��%q���+�PUo���s�q�A�B����_ӳ�0bg�0�+�W�m�*Y�f�FKu��%uncZ=Ȩ�}M��pk޵$�ހ����Y0�Wv��ɂnIRu8���X�Y�s��cVwr������D�ǝ;T�U���!��.ox��aQ#1{R���R�hjQaSد:���Y�T51Dя�kT5��+pƪ�W:ud+���s팁��?�E ���E���ȴwY���v���*$�"w0/HE�2[���n�h�� �7�t6�@�*�≸�Z�}j��j�����Ai5�I��[	G��Y��|9��_�8!�D4��"�v6��`�7L��"s8,���|?�iD���ԇ 1Ћ��v�Ɵ�Se�x�U����h6�0H;�3I�)��dnm�F1SH�5�uɞhk6m}2�h0�_Q`�����92*z���<�;3�#�����d�S��)C�\�2_E�E��+�놩�
���>�c�����/�火��� �(M�u��z�It����N�l�o��Z	��۷\E�I(�טz04Q?�M��ͨ��$�8��8����w-&���9����خ�����-T`�Q��Xq-��]�b�u�G������=T���7��I,�xW]?��Z�b?�O9�@F	�_nKy��� �-{�IT<�^����B�u`�/�4H���w~N �h���ʔZyD �˧�)�y�p�8.4�vU���%���h�;�]�?Z�b�~VZ���wy�2���QzJ:
�����y���7�Si�;��i`���o{���ܻ9@[_Y#�P�9�r�C��K�͊�y�x��^H`���^ݏ��M��9��{���a�,��5E�#�)�k٭���'E�X���Q[��nb����Ǡl�]�b�h�b.h`0u3��l�*�vWد�1�t!>���%+c�Mgz
P����#� s��k( �s�Y�̑����T� !���0FC$�a�*Z�ϫF6�n�����������NEv!�����o*�Z��jD0��v�s���t���A�%���mhn�k��J�,l,I��Fp�!~@Q���B}������;�Z�p�u9��'~�|��nx<���ÿü�k��������\�M��/r}���O�_+a��FE�x��z�9�(��
b�Eё{�pnjt���g�Z�:���͉Hڻg�X�ΐ��dƲ�3�QZ�M�����L��ÙR�Fz�ǻ,J$��"f�u�5�j�Hps~��m>I|���?�I�\�Kܦ�Ufe>Ji�o���x}�m���2���EB�o�F0>S��~��#�b��c���� ��Ob�CYv�6(�!m��wH�&0��������P0c�x��񩷊"��,�5�������;�O�I6��SS�~'��Ԛ��p���Cm񐃝��FA��oؘ�*��+��]�f�Cs6�m[�^�Y�)g�|���g$���J��P��[�sG��p�M���;������μ�� �1S0vT�@/G�w+y�Z��4��;�w�@h���:�ҙ�R��bq�`+凤���"a#��c�@��s�M����D���"��AM��@����Y��'���<;�[�P�j6��*��)�şx5D�T�C5~u��+eMf��?��8��E�=�|�ʤԇ�qOAW�m���%�ʪsU�;2�dG�z�X�7��A!��y�4]��N_���KC:C<����w°������4��d���@���_��|]�����������~4�O�-��b�����fv���(a�$6������#�H0�$�?��$p)�9�Ez(��� )�VM����҇'�Di�bp�؜&�) _�Gb|���X�[Y�y +?b��#\nb�#E���KR�2"Ɓ�$��ה�R�p�<+E�NDr�ܶ�z�H�L`��>U���lf�c�ڃrw�?s���h���F+��2a=<�ì��SE��󹹂���j��sd��ٯ{�@�a��N��z�:��=[/}eZ+O����
T�M�t,���V��0T���꿲Do��.��y�}��B��TR-2�4�>�Ŭ%����֓2��H4���I���X!5��ܹ��	�����(y\Me��)� �+Ǖǅ�.@)1� 8��z�?z�1�n2ʿ
�:���A��q���5��~�	7�m����/n`���`PM!~2f���ɼT��t�~ɇ4���c%��R��������#�q�0Ľ7�l(�"�
����g�d�P�lZ.M&�����r��+���s�����G��h/K��MYv�k"���q�R[TL_��QH?}ܙa�oI����@�GcƇ{�IM���Xphz(NŨ~CG7�k�b�f%���jr�`�n�[J����3$�f�)e0|��˗4߶v� ��X:���9f������Z����&�q�X�kx~K���3OuT�VKD'���45�e7��"{��e5�n��8�$�������˨ =��J5yĚ��5�^~>C��MU�m$!��rJ���%I��da�<ҡ�c�Pg�B�A1"�3�x�6���w�Q�1Z\?W�^��Б�4ɩR�(��ǚ#��ct�jL�U./����]�p7��q� ����N�Z�G8'��R)e��A�Sǻ|
��Qr[�����L�@>��K�$�5Q"�N7��"p����f�e�;�4��v�~N�و���$�2�b�'a
�{�����ː"�_!��"ÞI�ןܫ��]��Mg0�1Iq`s��a�p��o51&5/�7k&�$�I�K��-�R����ӂvg�ķI�����<ou���E0��xɌl�O��b�����8��z��,�+�̂��YR��\CV�z+��_n}f��V��	.E9�"f�:�>f��ô����_�(����d�re�T}�0��j9eV�c��\�n�� !�:�>���6���S�� ��e�,�v�a`���u�lQ��]�
=}f4�ed�~F�#V�H<əY���P�H�yu�٢����O5w6��<�h=�cwM�U���@s��
Mv�4x��@(�ř���X`����ioZe��E�?�4�Q������(��?	��
�0�� �	�Q7�S��C{�~ o3i&������ZT�`�,F�]�L~'P��,U?f�Bɯ�|�^'`#;p�A5�z�&��x+�8~d�ے��}6��B��9_N���_�m���Y˦Ʊm��R� �R1�Y���b�����e�8�քP���P3�>�V������LӔWF��zE�����$G���W1JF8�?�P��S�ܬ�{-�g��"3�邫F��Y�x�F���K� ��䁀� �MO�4_�ص�����.��M�������vu�:�`8�����Q��"e�DǀӾɭ�FҲ�<�����́!O@��>`x��J�(�M�<�M#�b��1c�m�/cL����r<�m�%�aA�CS>�����υ|DB�m��BG����b�����D�v���9��1�P�[�Ub���
_d��Gf[�WH�{�щC��x�0ђ��.���	Hpb�i���N���ݣ��yеP�j��k�#��./s��	�j�����y�w�G~ѭuV=&ǭ�'��/����7g�B��f���[�.��u�K��M���~��λ$�e�l/��jX!x:Y�i%5���0��ea��e%�=
���CTzfՁ�LdN�5c'�cT����p��8%�4PA2�*��f�50�׆I�*:�^E>��I�e�D�H�Bdˁ�]��R(dյ�Z�G�57O����޼�"��� _	P��������Wj
����@ V�pޗӂ��:�\I�����e�,�Ү������Ǯj�"�;Ё�A���-c\�p\�Ɔ�bl,;�#MmF �
�Px�l9�>����G�' ����A��fq��ywA�B3q���yX�z;O�p�` +�T�:Q|������Xdl��9�s�wA��Z�z�5y؆��	deW2���f�eY����u\P~s��<�� �a5�7~�M�&���&�J���#W���FC�)����`ӏ��v]N-���Cɲ��.fm�r��:���f��\6�sGC��p��ȁKEC!����E}��A���j�>�"	E��L��紹�X� [�����gw�٢�Z�\t\s!�4蘽p����+�J���<s-r!�K��b[4TG�Q^!�
�Ÿ�@�Y��h�����]К��Pz3VxC�x#V��N&�VQ���1�pQ���2ڨ �1 z<֜2/`_�4�4<�Gr�f�o\�FA�ՑB�ȵ�f*�*�N:�S^��'|�����/���]ϗc�{���z������7x��"f�ݤ?BQ�T!y���ڤ>Z!�U�����,z�k��o�n�?��o�|��� z������6��H^��k��9d��d���!�^B�>_���§�#4D`��+HO�3�*G?�� [�L���p!�����,���p�n}fVݿ^����@���n�
��l4P��S����G�f��,7ٗ�->��a|.w���Y?�������JڊL�Dre�vB����B��9FPe����o5$�+�@g��YĴ��v����!%uj��K����&��l|A�Y�$�8/�i�e��ܞ_`��x�Q̀~���YP��]����k�N][�c�t���p黋����8h�]�e�唑��#X�3s2ݣڙ�;�����#�2�/�߫t�UE�m2X��%��-��tSCn[K��c��h�W�~��%h.�p�,�O �����p{�J����nz��x!o�HaFa��Rr�F:ȶ�"��ϒ&��}h�=r��*Q"ms	��h9���2٠C�y���,�㮄���8KJi?��4�I_6�pc���6)�ձ=|쉕(�D�8<�$ ��8�K���-��Pg"�2\�����&��"�z��n��dR"�f'3ϴ������$�O�p�:&~��gu��R�"�Å?y�Y���'�������A	���\6'OGO�0���`T���Zi�t�<�/e���w;�	���s^dq�8��PN�{�%!j-�-���1#y�@��P|,P�j�Ԛ��K�e��s��?"�ipho�A}ݼ���"�;���U��\Գ�}"["�7.4�"t���4D�w��I�Mz:�k�R��H{��S_��4�C�&`�
Vj�܅���ה����*+ݙ������ˮ���
ow��K�2����o�6��D�	�����9�ux��Y�3�
`�꬟=u�����0��� +�njU��꓏�'h)���hJU#�����f~�!$\����ߜ
R�jw?���)�m�ܴ�
�3�8��#�
\}/�t�L\�&� �4�(;�j�9+�Kx"���ؠ����ZB�v�"��Q�U-��?��HBG�fx�F�A0/I��MR���9�G�o����o K�xj/����V2gQC�1�s�'!��s�1=C3�J^TCa�BM/FD̝�^�:/'�f��gN��Mnf��.���D��A��Ld��2������6d6>��
��%�">N1���dm�v��,|\@"ȫFh2)�`�/z$�u�1l߹��2R
��I�"�M�t?�>��ƪ%����}�Ug�c�]܁�j�F\�����_�y	�V3:�i���[,^�&\�3~�FJ2b�HL����Wk��鞯�9����Ys�������)c���/���u%؊+	�>�ﻘ�$O�f1T�ƋY��h�����ޤ+���F��2݂ᓤQ�MVJ�hF��-Ą���=O!�= �1G���!3��c�L��o��>�����KSr��2s�	sw��,kCG��E���;g�U�/����O�M���=��1W��>61)+:���]w�G3��|A�u��O>��p'�j#�I�6��8|�!pU]9IX��nx*h7a�w/k�c�U����H���Id/[�d=�?���J�A7'�z���@(��i��W�y�d�~�mOE1s@Ͱ�ҳ�iu��8���B�)@�\�����l�W� ��/݇��{�Į`�v:1E��X�Xp���k���u9Q�1�X���/�8'�\����0�mL�̨Ϻ��Y�F��A�����	�Y��l�+���vc'	�Rw����p�9'�ǒ�3&~��]$Բs�HFz����v��6�0����,2
1V �y���Q��Ō�`r��+D:�G�܌s��;�k�B�&]8���H���2�,2
�S���6�2���SA�s`�f�v�Gi��g�ɓ��N��t�d+K���+���9*��O��i)��Ⱅ�o��P����iL��5��b�	o��}
H�ap&)k��f0\����e�:�4�)�	3�5���ZZ7���`Â���D8�Md�V|������ 	���#�4mL��

�E��SI�Ć�z���<�.�v�p(%�wd�$L������ÿ���"=��fW�fj�΅'�b]/���iŃԠ.f�X�P�K>P)�1r�&�A+gO̿,O�O�B���TF$��S�ݪ��?��pX�����@�%�_��>���Ĳ�~��O��{��M�<Yğ���Q�"��#������������7?�|^�\#��7��80Ko�G�`�S�t¸8��R��,ʈ�M7�d�)4�ˤмd��xYQ�XTu�u�&SY�2ϫh�S�3�~����*
f?�c���C	O]с�{��E�Q���gǸqn ��FVw����*|��~�l��
ƈy��ê��a�H����.0˦70�����(���L��F�r���?cƋdN�a/Y���~�@�4��'���e��c�o�d�6f�@��ӏ��aF+�~zȒR�U�5�d���]���m��l:��8k0�e�̎��r=o�]?��^�d��{� �0^�zx��X��:o=u�q3��ʾ �b#�J7�ͷNj�/�lj�K���j?�n*�G��;-�+w� ���� �{�q��	pk���u'����T��Ew��'����SVdu�J�F�������x��'Gm�4tw�\����l�{56��"�`��y$�ɐ��.Ùӫu��^v_0�~�{E8e�H�H�݀�
N�	"R��Z�"yl��{�[ޱg�ISL��_ i��-��9��m��܄ ����l����`�u���+B0�.H�z��N ��T��~�P�W���N�&��w�9|͛�b�:'�7.ʜ�9����`���� �9�T����Z�wX��	
�Y�>�]���[Ǣ���5
���g�x;X���ߚ`N�L,6!�7g�#@�o�@��A��e�(V��ɴI�P"y�Q�~����Il�)��\�-9b`z}�i��G�E�7P]wJ�b������eq�&}�n�xM�r��ל��|�?��iџ���>��0d�j+]s1��2\��T��M���7�?�C����I2��R�5
f/�d�<�!^�?3�����K�P��>B"�Oz"�fU|��}1��oO����Ï{�L�y=ybt�I����_�L��^tS(��B4)K&b�#@��"7�D���:j�f���F�w�K�@l��w��uꤲ؎�8�[�XaVSDL�L`��_��bS�U�7�IR���wB}S��`�E�R� h!�E�E�B��������9��ՔiN��'YU��H�	���! 
-f��w-��H���!��=��C�)�E�V�%�CTـ{n{���A�e���gy@>5����C�'ڛw�Ӿ�&��@�\M����U� -�����/� ��׺[����\	g̃�c(c���� 0��S��+�EB���JTa1N؃F�:gG�x���k:���.8��jm�/��^6�n�r~�T��H�7��.t��
��ᨋ�7Ɓ�[g�D?xu����J���J<��r �	�� &����V�zD��4�~"�e��z労���:��?�2�x���Z
�Wi�P��5:���[i�i�ಾ�'i��9�T�TJ�bV���m��7��Cq�Dn�1�ϡ�x����ڔ5���_շ�Te�(6V?�)�`�/���`�KF6��
S8�j���E�Uc�8]NWII�^T�4���5�P�s ������K�93�k��l��<�A��%\�_E�h0�ux�}z��d�l���硏*j�t�m�h$dY�Yr�`"/�Ԉ��Q�ú����#�$\��l�k���N�7�ߙsrv�5�Oyn�D
�ۿw�]�o��d68�q	�(�JK��6?�`��ž/�HQ�
y=���dL\FL��������V�W
�Ig�l�ة��價&��f�T�5xv9bh��ޏnR�@z��;z��P�[���ê֒|��@F���%���^�����U�s�o^ǫ�b�p����(A�-�u=�|��r<� ��&}� D2����ᵍ�Q}R���G�a�=��!�r�zZ���J(8���~��g*ܧ�]�K~\aJ�o<`�`��qO�%��lj��sI��DY�ǜ�ؼ 26���Q���Vj�BT��M�A��'�,�1�?�lĺ0���UD�~N�r��� ��S;�&ח0
F�`�Q�6}�ї�+)�a�~7�*!3�� a�U�5�U=�-����B��@*W7{5Ғo�y��)��2�=w��Mj����t	�/ wQ��GKت˿�y�w�/���>��qV4'PfS�YCe����7�'���2m�x�L��{˶�w7���ӻ>�K+�&��#��g�/�}��T�t%A�a�~˕�����_$����>�2��Hݖ��k����9�w݂<Y���k�uz�&�G�/�O��=T9�Vne�:SL!������`��*�;���C{pw�"*�>\��H��Ӛ*�a2s0P�[o��̠�;����߼���jP�Q`b�@G��Q��,�SӬiU�Q�:Zi����x������^���G�Mu�v_N�{ͥ��=�2m^t%��AIѴ(�	 ~����%�Ԭ*�Y�a��.qF-rF�\\�P���z�<�?;P��$�Z�!���&:��H�1��MS
��\��:/�b6gZ���n�(th-�h��ڂ��؁6��ճYu�S��{.p}aO�y�.B��Ћ>3�����i�ڈ�ȞV��g	���[o`�z���
H?�L�a�'�?$�M���"ߢVD�8q[��!k=�a���-)݁���:�dtU�iұO����w�`d���k��ZKߏ�̸I��0�;|<3'_�)���ciA OT�AA뇫��--"	��g�n��m]D��<�����?��9��XZbT\�m�ڽB�����s}N@jF��S�_S�\�-�Bϭ�N$�
�K����+�3�T߼3:\y�y��O@��]�j�K-�d�WZ8uD:&�o�h����^8�#�X��l��F~�1,r8E�H<�~V���:��h���j07 z3ʕyx*#�rc�UmW(��;x��^Ʉ�Ӄ��ᶮn?�gj���-�6�:}&�kB���^��8��jx�P4X����R �O�l8ua���bE/Z��.0�������W���뾚wx� Gw%Xq�'ƌY�-�Ef���B3<6?�x���1g�E���"�L���K���\��7"�}�]pC1c��V�a ţ3x�x\�:���ɇQ�C��Iݍ��]��{8�vё|����1�-%XۧR���_)�%�p��G�mE���<(SƸ#���w���)P}���3|'5ph�崐��P�p�}[U��,���n��Y_���(���}ĕ��7�s;��HΧ
0��c8SP���r����%d�ߦ�N쟈������p.�7q{W3_�餐����a�w=�^=�Js�QxOD�'�A��M� $�E�='#�fx���5ca��0�촹�[o��}����q]��JZݞ��Ċ���%�'w�3k��DT�]�H��E�*���nc�Uù\�ēQF5��m�!������P:��0Ԇ���!h5��q�BM�	�:�(��e�H��[_��7L��Iܢ-Ԇ���#
GˉBr@��B'O[r%Q|C������ט��g��g��غ���P�yW��i�5��XG�Yh��B�>Μ��|����Zb��uH�8��<0eS�B=��JN��Qr,����m̱L[T;B�r
��K!��As���{�M0��v��; �,~����bZ���,�We`U��Uc������ԕ�D1�A�G�$bH�
uz���_%#cK`׿k��(:���]i�r��rh�����$d��MՎ\��Dt������Y&�]�	�����q���H���M�A~:ֵU(�w[���OnA��O��W����� ���dH9�6���U�uz7�0����G�������������;��m��P��wE'�7�J�_q��N#�$Y�:�a�If�2�IB�@cO���}43]�����Db4�����,7�(l�݅2`���c�z2j����7έ�2���#6�n���y�ܙ�غ�zzS�hg�E�d��ySУ�_U��Ȃ�pՔsiK��t��<���Ȑ>{0��|n�F�$�\�τ�=��x�{.,Vժ�;)��=���Ȣ�w\b^û�_�xX�<C�Q5���9k -����m���({�v��%`��DjX���j<�'�3��P�[�}ݒ���Ե,���2��(���ݱ)���}.�į��������"ܻ�^���ݜ謫�H.h>�g�"ѹ�  G);�]�p��4�T�>6��ᑍ�'o��d�v���k������ۥ�CK���w�>Al�8��-w��c�� ��\�P�h�$�k��Q��AT��L�3燌)O]��N����?P�1�����3����أ	�]�1�p�<,���q��k�zDpOv�tE%Վ5�|�$�����%�t��,���S"u(,���I#J4S�n����8���6_���)��_v�Zx;bR�����h���Vy8+d���De������L�D*�ƴ&m"�5\�#��ˀm�c�����)��킙����f��s_	A��Ð��x�����s�uJ*���	*���1�_��+�ݸo�Wz魬��Z&�ȕ\3����6�A6� ��uH���8?yߖ%��i ����\�An��3n(c�[,���()��5��e�������Zi�ȉ
݀�'?��V��3��L0�a)�!�>���1���oZ+h~aB���U��d����{X1������C�Pg�4a���&=A�s�{"E���e�s"�]�/�?C*��D�V:��B���^Hsw����3�?6=�����T�_���}�+;�br��./xt�CdWe����g��h�d1�j�+x�#�*E;!��>S/�����ǜ�E�J���:U�7�����$᠍��0%���?�_�|5���Ȍ�j-y��H�ţH��+�ՠtP]5!�&�XX�����ab4�����|U@pN�&�L��č;��G�9�hdȀ%8�{������s]R�����f�5�[�s�e�e�6�
�t0���Z�f=W����Kwμ�U�����T-uK�3F��2�'`��2��8�.�.�Վ,�c׷�MS�r|r`���a�a+Y�Im�4���n��o�@ȜM��5V��c�z�
ad�\k��Fb��P���bn�A|�ֶ8��,�%:n�\4���e>���qI�y���Ɛc�uF�)���`~.�0��_϶Cӄ.�@���燞���&u3d�$:��y�x��3�r��Zo�;`���Yx��w�6�����-�РgH }�0��ʃR&�X�'�^�@��&�怅n1�d1�}���ϑ����t����:�����8����a����o��˽�+�ۣg�1�}��*�|Բ�F�v�A늌��d�v$y60��h�0���OAn\��^������-���������`��Պ%�@�y�jǯ���T[��R��zo�\c�z	I߻�ho��0@8�Pz=�H9iw�n$��,e"�����4f����U����ϟ;��Z�6y��)�.0f�g�ת��t�����6 ��F ���z�ն	���\&.}�2{��G�%N�2�&��L��ɝ�܃�G��p�B�<��R-WΔH�1��+� Vo!���k��C��9�U���0r�RlԸ�}/*bf��)̺ܤ3��>D�{�n��#�����bN���R��b��+�Bi��G�sl��䷡�E?���u&�l���3�q��g"Gw��8�a����20�◃L?x%e���!s���ѭ�dj���k���i&B�		4eo�!������E���J煉cwbju5+Q($�e�+H����ən�@�O�)���>"n}|z���e;up����FEs���=EH6#���Ty'�
�
����ST8?ү��=~8�� �=a���h��zI���2'�Wb.��P w�Y{dR��2�������.Ty|Iυ����QHR��e`;�㊯��x0	7��d��a`%D�v���5wBJ����E@����M�S�<�}?���4e�<%q�4�j�I<<Qu�A]6��6 �UWJ!�EQ1T)p`WltR �د�A��@T��B&7����]�SЖϑt�)�Ň��y�ʢ�L=���K� �W��C���3�|�c�coW���U���)D�r�_��X�'&ʵ(
�K�o�)�lv���JVV���n�9�b��y%�tm�G��W� ���u2���k��f8!��dl��E����z��<f '���IV��([���S?�z�[ڣ�_X�vOr��r��,=���]O�Cf�|�HV��z���H���⅙��2���Uy%���,�2�w6��~�Sl;��I3�a[�E8����t**����ַM/�V���k�@��'P�ǙN,2f��v���KY���{y��Z�3l3>�����EMI˖���S��=�5�3��S�nѧc�Dط)˴���%yN.S�NX�@F��ro�W��k��\F��?Y�+��˵H�"J��{WE�%�o���R�{��Z��$g�~�&��9"9�>,d�pɨ�qk_�>U�%>V��-�����c���=o��;�Gn��Q�i��s[m��$��3�.7���l����� ԇ�Y�0L�X �D#�����.���W�%{���(ӍՌU�����]��l���6�I�������db�^�f�����;ȊK���kR_����� �m9�8Ւq�*f&��9y��;Y S�Ž5:�LݼJ{|�#��hߎ��ދE��%*�m�M)��l�N�G�[�M�[V{��Ԧy�O/�~����|c%�j��ɩp�.���m����QR��}�1������U� @��B��dw�fEy�����@Fz�do�u�32@����Ҝˁ�h�dZ�&���qlٰ��c���cb)8����Ꝍ2Xuʭu�S:l���˷�:�m�̃����z���z��9g�PN[E"��T��M;:��Mm[H�h�#����+twc
9�K�=`��R@_���֏!mw2���c�f��Lm�iX��Ԡ���u���?g��@11L� 4$�_K �[&�BӦ����3P�ɍf���g���k��B񡌿>�]S{E��ٸE�䤠(7"*��z�S�_���̐���+_k<3̼���o���bbYvG�R�,$�qX٘Mxr��4TK�8�-�5�Ѽ��G��P��iC/<2F�����Ģc\�|��d�/�=����Gv��re�,N�ou�ЋB	���$LO��qfvX���/z��r�\����s Y|��~��Ҽ�=�RX���Wv*�T�b��L�6�U�,TT��|BJ��&ȿ�@����wm�O�Sq4%��kc� ��,̖���y����ΰ�}�v�^g��>������pK�)� ���ޛ��r#�^�4	����i����%Ҧ���68�q�]I�/����	��w���+��D�~��8L�D%��`�S�\Aӷ��������
��3�������qܾѿv2�|�]�!{qQ͗p{�~ 2e�;�v�{#r�B.դAC5N�U ����|j��;a�+V�UK$�<c��3�,M������Fʟ?�n<���Eo�2�ك6A��L~MQ�Z��l�a�IRB0I�@�ۨp٧��1޻���qp?m��S���E���aOG�j��c��1��Av��~�O�^`����xh�9>-G'>M0F
�g�fa�!kB����h�D��R�`��lry�����R�"wI=^ܥf�� �@�ul9:w,��4�3Ae`3���ʳ��>%�L���9C:1}�Q��Xʚ˭�m.P�'n�T�;HL~0�bėu������ ��xx*��6�&�h�u=�K
I(XS)͓�H�|w�]�2n1ά�R\�B7�����ކ��z`���ż8E��OuO�=جS����d_����q��Ɂ��^��X���^�00�7��O��ƙ	p�uC5�������M�\t�8DVh��P�A��)�tUj��|��+��{zB�҂s�w�KM	LD��#<à�Z}�/��a����=�1�"M�q�8��"��RC�ꌕ!��?��h�Θ�WɌJ�+�2iI_M{�����$xLȇQKff.4XZ�]"r���>d����(�)|MM��3W"�SR��!�_t�Aa%L���v|��X�][��ڪK�Z �&r��+	��<�:g{K�szD�
D�y(�>욢ږ%��r#6_�z:�u4�Ia3��]%@�H<���������?������[_(��l������LVmb��jL(���.8�T��YGW3��L��P�3�?���`A$|�}��i�\�$EA51���]�i�s��2n���[�>���(_��]���U ��{��|VĞW��U7}Y�EBd^�FQ#��p���;(��޵ܜ���c>���dq��ڄkL�����D����jh�XZ���YzB��ٯP͑��'��yJT�Է������I���G�J���bO��a�8�ټʐ��T-�R�F�`�q���ߚ�8�?�k�&�)?�C&�W��Fz}M�.7�l��~��0�m٥�=.m�55�m����!�T��Bm���u����y�\��P��;���I����f�Hҗ����3O�$T�2��D��j��9�Bs���!6��+FB�4ȹO4.&�j��mS���B��,]���!�~FS�$�Ŏ�Fh���7.ķ��h�o5-N��oo@��n��(����\N����נ�Xa�0�{+�Ĉ'�鶢�T�"<������s�+�	ܙ�0ie���I��I/r�$�gh��>,�q�-��⾫ $;�p��3Y9�V �>�S�1�pHpʒ̇�F@�	���˺|���B��ƸKg��@(Ŏ����g����4ީ�x-
�g �͋��UY[�{G�Tr���Sh~1���;Ƥ�+�p�ύ�;|5J���	�xy7���n%Ma���=����u8���d�{��
>0���
��uD1�~:�<�Ii�[�=��]k�Jgv���~Ia�f����9���u���E��l���J6�s�����*�]<x��0�φq��t���+�;\�Y��� ��θIV󿞆��kl`�|/�IO`��|k�+�m�x#�+5K_��ŀ`ܑ>�2������b���V.��i[u�D#2��딘\!+fz�Sif�}-^���^�u�'#�l+�8W�vn�I���1��0߼Z�����\ɼu�D��m��\��i��G�EN��TbkI�,l�$�\��~�^��gùG�(�,&
][��jpl��Qa�H�>�<�W-���v�36� �u���I�fl$��CEc��}=��O-PHۥ'��$P.���2k`b:�0��XT?k��g��4%gw�0�{�����aG�,�y�N�-ɟ�P!�=�(���|��qz��kP�!�d���\no�	�� �Sp��PlF�~�s���N�����Oд��Ч�K�}����O���؎+fb/���"h�3dY<S�~1y��sgʨ
�a�m�o61c7�h�[�m�D,�&Ú�h��k&�Z2�_��m�C�P��.wFUI�%9�'��k/��T[�����~'��9����2�X�Ė����������-��?����T��UW�d4U�}���TS���?���_ !+Fs\�P2=21��ʦ^��țcQӶd\���/���3xE(lZ�F�t�i��:��?�z� �9D��ǻ�NC�1�����D�p�6(uf�b�j,t��')0Z��E�V���Oe�*�{�Z>�~�/�_��DS��a�oD�"~� hC	w�[����7�U�˚����y�E<^sd��ۓ�@��10�0�F���f�)�ߌ@���X��,p�~��Z�@f��D��H"dP�NK i���u��3U�0'v����������5�3]n�o�&	���	�J\�e4^��{���c�H�@:��u���qTt�hf� д�� �&>��\��?<� .��HQ[�}��F��J*�>{,�F�Unm��.��F�|�t��B�:J�*$�y)�;�
����s��*�'��hN��E��bF
�uo������������e���伡��fVsW���=�U�we�z� �:�U ˋ)gP�k	������8
Q݃Հ�㘹9���>{���K���4y�{�%�Laԛd-i��3����BV��B~O[
 T�Y��_�L.�d�۽��(��ǋ?\yZ?7X{k��ן�ľ`w�{��y�C�Í��[��;�b��`&����B4�×��;�G�U���%��>��� ����-�c	���	e��z�H}<��д�װf�o��b�L����FUk�H�d�����%[���r]��'�^�%��-V��2��"�K�:�v�� ֗��}�9XhH�O���Or��z�d�eF��E*��h z�lhw�ãy��X�Bt�`��}N��J�
��qd�ķe��k�����~�h����v�<��{G#�(�3"#=�e�qM�̅�@�6��.3�H���k��Χb�ֵjP�};���A
#u[�CG��~��6�n����T�ڨ�͗Ѥ��%��q-r;�&]*��TP���;��H���+��<��xA%��-_~W�F��ضhi�UjS�]t�D�X�bt��>�w.Ƒ����aXr�dhB�!J�u�>���%�8Z���>*�'-�9�J�%qb{���%�	�H�����]�7��M]�8���VQ��L�o�i|��?����d��3���9�J!#G
�'�D���L�ߌ�"2<�m�)�v�a���ѻ�G���Sl���?tv�+�[K�l������Z�^]A�|7���Q�#&=���Ai5���� pS��%�»	W����gXoU��އw��:w��?�7�Iˣ�,���oϕ��ͯɓ0
���%j��HZ���߫�}S��Fek�&P��W.��ɡn]{b�6�Q S�lI��u
=yEhg��a�?�873���&�eȕhRM�:����һ%�L \�_�"S5!���k��gC�9�k���!R/��#��k�Z���A-�eQ��� �w<�]=+�s���`sl�B(2ʷ
���i�-)M����Լ	��Us���0��.�~��X�ލ�G-{�rjIA3��ēZ��7���su]��/���l=��G�Z�O:m
�;�J�vgMы{`c����|O��MX�������;�Q�q��ά� �'[� �߿�-��
t,|y��z��k�bצFz�vq����o�-$�um�(HU~��BEy�'l��IR8f�^O�"]�����v)��nH�pV*�~�����s�'�t�K<�����2�o�lQ���)��D��t �j�4'7T
2{D� tN"3���@� ��p�3繽�G����v��TEw�����Y&�'��OB�y�d"6���P3�iƱv�Ry�������E�8�Al�>1���n��&�F�w��l���_"��}�go�k�ݓ=��g0W���AZ�%F�����td;!B��!p^c�h�h!^�����^�%��l��d����f!)��i�eoҎ��uPt�^�4$3����*X�[v��a 7{�@��oT�M��������o��1��TH��Sp���M�`��C�h���Nؤ��K�����`���Hc;�~^�S;K��?����C&���(dV�İ����1-|a��Z븮?�IQ�]+'_WA�:�./|�-o_��P���.:KY��t�W�R�LY�M���#d�6���ǷɅ�$ͮ�~�'ٴ�+�˸�� �T}�`3�`O�EЁ���J]9��?�`.Ҩ�^�g�e]��)8�Zʹ؎S�G�.�S��󛟙yt�?j@A�ʌY�xg��Z������%˼\������eaP��]���׻9�1��Q=)�{�ʵ�]��`]�J�_Ka�#-b���H�w���P��	}�������9_R�ڋ*��%O@v��BmcEjAwph�w�Ra�h����òc�%O�}�o�K*����q./�C���SBi�4��Xk�$�������&�N��'\�Aˁ*��@��J��5����G�xѓ�T�/c�䫢�b���2_L�!H��i��Ӷ�!8���4�����L��I����(� �M(����[�Rrհ����TI��6X](�[̖�ltcxPu^
��|M*r7�����<�4ߢ�=�_�m�G�1�a�7�,�ɝ�I���q���[A�w#��HN����j���Ƅ�ܪ>��q����K�5]���