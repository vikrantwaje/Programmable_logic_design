��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�y�D�/ֶB$��Y
Z���E��[�@��T���&ڗ/��H���b��.Ͼ����KClL>��DD���7��h���O�+��j�B�xP��FS�s����IE}��o>nxo�vPg�I�\������Ev,���N�x*�Sr��6��:t�_Z�	kz�f�u�@��ϫ�؊
B�!%:=��tPi���0�$Ŧ�X�+XKZZ*J�� d������a_�u}QV��{�Y��y�'�5�6�ЫtO�!��I�����,US3��o���-����SQܴ��<}t�Z|��!/�Y�䲑��ǓU9�9��w�r>x0R[
A��-.X��2J�Ï1��G�$o/��A���a��ԥm��[��!>�e���{��4��^��o$z���*��h����'B�E]�9F�ʵ
�IԦy��&Y���a�!�3]D�L0N0Zvg���s���S	��nGg�A�4��r_YQتS'P4�u>7L��s��c�Q��[�4?u�zE��|�F���OqE�����h��&�L�'FI��^4Wɚ%�;�owб*�)�[�onv#���-�5�۫���1�}|#���݉ �����4gr�m(��ZIǔ0�FM�
���d?��O�����t���̎>��v!lH'(H�z����R�X�f-;�Gt����P�~a��N������V����%�d���#gas2�A§������@�+����-�v��%�S۾ݱw�z�v��e��A��$	��9m�����~�#�@q��?��R�"�Ԗl�a�ʣ\�T��F�j�4u�o��U:��<,���1q`PZ�<�"M1��Z�Fp�M�1g��9ƖP�S��X'E�ߝlg�8�O��;u����ѭ�ϵ�+w�k<��>IMB�7�I�ꯠF�	�?��),{��	)�>�S{�o%����u�:�B`R��0�s&��[;Q�#�NMb+��ܗ&3���� ���@����'�Z��?��
;�mE��������&�R�ƺp3|^34��}Kq��uܢ����x�����_k�@���LU1Ȭ'N��,3�nË4��.iG�%��n����nĚ��6���r���94m,x��툘��T7���U[���%#�aݎa͠��k�#ƯX��ׇ�Qqc�$���5V]�J ���a5�~���v��I�\,i�SD���:��v�I7�5�o���`������� D�?�@S�S��#���f�/ZcO"��J�����pN[֔�ut�?+ �ѢJ��SQ=��Xy3N-�T~/%vl�,~�ض|��x�@�nb�wUB��K�IЩc�^��U+���.��}�O��%v׶f?%�^	�����z�b��x�Qϙm��8A~�w�O���OQ�~+�_��ّ���R	�[(v��i�QTqj#P1�=���Oy���5T�,֮ʡ&+�ЖD��	�}���9]]�e�?Kp�G���c�g�ܰL�O�0`�����F��h��FO�	�U�X�I�7�B
�ҥ)�ӄ���v��*n�>e�]ٲG���|1VzU�y����DD^3����AC�W1�a�2u_M�B�y���ꁈ'/ĉ����j
����<G����N�!S�.����jOM�ț�,a?��v���v���^�Y����=�F�ᝉAO��C9��ڸ�:��9�ISy<n��c`�S�p.�����ds��g�c�:��ТLb��0V=�*n������g4~/3�����*J̵4Q�Z+*V�Hm�)7��
������O��mS^
������%]}���Sgi�(�����C��{/1O��I��+�\?Ԛ+Km�!�j�20�N�4��=�Xs�ti��A?F�ߞbe[F_��r{fVs�S��W_2�C���b9 �������/] Ta��蓈H ��mW�H�6�2a���X�﬙~�F!=�"�!����H澋�i�:�sJ/S������S�M�|�_0��-��NH+��|&c����T�*J��+y0U���;�|ԐL��A�Q3;(���Wo�  �QfT�͙���|����w}$�����3)�(t��,�c�=>"s����������V�]���V�B�/�`$�@�M�[�
�O�f�'�&Q5����wF5�Ww|�p�������^�����!�F�ջ�v�O0Q�G���%�����:Q��r:���U��a����\y��;��"O�t���+��?2�&m|��%f�N�5���J'~�SdO+>��Ф�7�O�3FDP;7���i���R;���p��I���V�Mt�xoE��>�5�Wq(�̊�Q��<��(��	�ϐbj�����4+�WLp5�:���=X�����n� ���f/�������ˮ�8øʟ�;�1ۗxQ��	�&�_߃��!$vZ���*��[��Ψ�I��M��nͪ|�,��:�m\k���~~���*%Z���O+��Um|�\�?~	�wTDJ����)R�F5�k&���y�<+����أDz\�� T�oH{�'�[4	���_�]`MG]��*nZ���}����4��tߜ-�D�[���q"���@X�r;kM����8�@2�<ɱ�=N5IF��"�>�Į�j�1��ϟ3# 鏢�
��8�Y�N8�^R���*9�)3F/ZXF�	6J��IcB��[�j >��NR�Zs
�����di�K��(��#�H�6  1�}U�����ڼ��8�w���߯$�{����gƙ</�c��K� ,�z_יH]��j�0%,
�=�AΤn�lp���'�>�5WZ��q�X�/���'��2�V$"���ǂ�i��/�m%}�ѽ�����6!c�|��R���Elu�ǳ��:Y�䊓�ߠ�k����_�X���z}+:=�#`���^}�0����AU�z>�L�
h�X=�!)������g��A?G�Y\�0�����R�y��x�*�aD7���:���uD�#UC=^�e2$Д5g�MH���Et�S��c���|���|��Lp��#��Y�2����ڱ�`�'��4��\4�j)(��|�2���l�s,�(���DGog@[,��jK8�^�u�}��}��D
���� z�'7w*G�}F�q?UL7�@�m�w���5����GC(C;!b���'���]��r�a,x���1L]t�h����o�(%�d���"Coʙ x�sq.�V�iU.f�(K�	Z�˔��)J�xH�`�m\����K-cd��x�56�3�dN��b���2�_ܠ���F�dD�E/�SY\�*��=ǣx�/�gXz_�c%��D">��?�<F�]ӧ�hB\���6��m��8��&���^��ؐ������D��0�v���_��m�������_�h�8�g|�^�	]�7�Y���CE��A	yz����=o4�y5�VX	eT�V@�(#fWnek�R��S4�Lz�����w������x("+�Q���.�q5�RQK
�r$��r����zQq8r$Z߹�P-���Z�9�,X��k=��0x�����f�W^m��)62l�)'g��̄�tCh�=B�C����\�|�ĻE�뱸� t)'�i��-��u�Is����x�;���P:�dc9�7)Ҵs$w�&���4ƫ�;8/�oB`6p��qd�����fb�Pݹο�<	\&�U���#�fe�y�:��޵�s��O�|tX�o��Å-��'�uf&u��^}N�Up�c�Ԏ��~#��k������3(�*˨�%5�8�@s7YCl�}�ԻЭ�m���rT����	��D�n���&U
d��dQ w�D��h�4FB�.<��Y��$/�(����8�U
�y��Ϋh�r98��2�rM�|�1������9�T�vi��2v��E���lM�v�Vy�ru��vk9"$� �;mL,q���~%��v5cG�޳�T����ׄ���F�!�#�p�vi�q|���J-X�bQ�/R���E:k��$z��M)mUw��k��Q[-�����<Պ�u\>N��x�}i�*�7f��#'i���R^�,��%�$4�ܜ*�!����DBi���G��$Zv���ʖt*�$ٜ;aV�.l^��1ڑ�o8�L�ɞl��W��+lB�'^syT�)��(�/).���,Ϣ�3�����.�?f��I�4��^��O�����#���xFT�)&Ì��v2b��{�x���D���H�.��2����s�MB��}��L��y���l��(�J��<�mP
�if���BIe�$
�8|x	�� R��3+�8b3�lE8[� �=�ɯ��
���0q��5����$�1�+M�ɍ9��Z�w�~#�V��E�{�Č�Q���&��#��[a8��z�%>H�~Ԙ��m��@b��a/�"��˟�� XM:��i���#�8xm���}��,M�����n3%�{كa��NZy}�*���M�I��A��6�"F�! �~�E���������|�'�Ƞ��BqcF�1Vi�� �I_��le$*
�y�g>P�9]����[��Q*�|��Zt�j�7���P#�H���o����P�:6��v �Z*�����{�E�Z�BX�2s,�+Д(6�'���Z.��!vXm&l؅)�%6D��ʫ},���`�v��v^�)J�>�d�}�0�z�Q��)Qw��;e�h�{zq@*�D�u��.� �`��~�Aǜ�t�dz�ľ��6B���k��"`,�/;�j�/ �P�8����6�	\�~��᛺&�>6U�>K&<om!�lj�3/��%Z�6�v?��Xj2��v����^�70�-����r�Z�L�������hH�X=�SE��'(���M/�=��^�r��C��MnLu_��Uʫ��V�\?��ht-M�֙F:��Pm�c��FU�s��Ȑ���^[���ӻ�6��=�`< m����n����s]Ȟ��p��� ���>�,�;��eF۱qp�)�D !Z����^�|p|	9l	�,@�W� Rn���lŨ���X���s��VJ�O#S�bG��f/��!tD�e�h6��-Ow�N�3�F-�� ���R���:��N���hC��M�xU�^�`O�zظQwYvBc���dj+�N�p]^���3N����)2�O����!� ��u�5pG�s�ab�<*���/��+60��[g�q.X��?����x`Z� V�+l�7�gK�m�ʥͶ����Hd��~�)g���8!��0ǎ�S��ۥ��6>tp<�F��}�5�LN�5[�M�N�v3Y�jrW��_�x"��� �6~�̊8�����Ӵ�&����:�������m�@v�w�����p��D���ܥM���%������y��fR����p�{��س�6q��cSМ�Ӓg�3~}8Z!�p'������`���! )� 
�Դ"Ԍ� ;�5�fh���Iq�͍�d���I\D3��4J��|Pdr$2^g��w�?��9J�R�K��R@�3��%)_�ATm-<��n�-�ئ������~S���(6��{��e�Q&����w�:J�ض�;��t���O7������P�<Gf0�16�����#���k���Ϣ�Y_Q]�`I�1��:r�ݐLi)_ͲG����@6-��� �X���� f'7l]�Ak�Jw�M���x9|�KpE�j/����g�PM^*J�p~�j�!`R���.�?<29v�`��,e5Y�^D���B�
q��?Ór�ЪӪ�I�K s[���=���z�u#-���:x��l:�EHMA��7��/��p(�<`���ƕ-X쳉C���+�J[��:���-�����b��r;XKbE���	W��/s%p��A�~����B�?9P@��u��sV\L�l:�ۻQ��bN~o`Y@��.��X���>��^2ԏ	w�Q�:���\���^>3C$]N��襛3�PL��0� ��>{��{D�dT�&�d9<	�U]�Y��6��OĀ�/�-��y�����]��R���t
�+_,��(W��c�5A.ߢ;mJ��K��5H����]�/;�Q��Sd.y�-��)ϵ�'��!n_�Wr�����n٢O����*��N�Fxٟ��ȳڇ*/���Z�����?:\��@�r6x���������B&e�j�F4t�-G}��R��Tdߟ؋�%[��!�Ho���[�uU���C�Ǜ}H ��#��o��gI;̘	�V��J��&�:���'w*:�7�QU�7�Q���^�5"��zB�)vU���[�xX�]9r���~�	������[��"=��$�S��ȡ>�>���Y`�/��(T2�����~�F���	�_�A��� a>sX5'�H
�"�U��w�if�ynj�HX�˱ua�C��
v���6��N����)p~g� *f��!�J�xI������R�tͣH����	'��l�þ����:�0X�ތ�����Ђ���;�z���l��/�NU���a�Gp��;�R���IеY�1?I�W��RN��U��MF�v0���+Ȥ�]%��,���dN���<��I��"�)�F�F�R���b6Pt��k���nd���u�_?a-W&�Ş�>����i>+�L��qԶ_]�/o�� ��Tn�hUF��3rK9m0�N^*S8�dɕ�(�>6��ʲ<KY�
�ո����,���b����lȜ�?g-SS Q��Z��v��<V�%F���c��	����T��G=�#�"x9�O$�n�\��C�ib��ri�{�
�$�h[�B.��0���2�vN�+av�e�,\>��٣[iae�[�#��T#E5�/���w�\���k}g1��fWDU��$�����P���t��MP�-c�'�_�	�x�"����]m����MX� Jp]`a�Q�T r�-�~c���ܜU1 ���J�hOE�ּ�v�d�/<���Nj> ��r]������47����9U��MYU  �N�x��<���A���x ��|���~8��~=bw���7�l�;M�ȡ�oՙS�"@���7�7�yV740��eU��AFm|uНdJ��4�U�݄j�о�m;��U�M/ҫE��E��Z�7���Μ_O5�e\n��J*@��$�0'���Jo���֪\�]�
�m�Y��`f�=�ٗԍ���!�Z�ǢB����	~��{��њ ma	��e^����"U�JⰑ�]�ٌ&p|��0:-72L�ew��0��G�&v	�,;f�M��η�F�f�(&��T����$XS�ꊣ��0zB�m�y���4��6y^*}F�n;өs[�ER�/6�Ke�z�[�Y�b�X뾅2h[�����.��� ��䖸	��Tg��7)dב0R��Oo!Z����8��ע �9�>-Ġ�o%��G��m�$�|ǈP:Bi����W�e}	9�B=����?;�M!a8̻+A�rn-��J�:=��#.�\˻xp��lu�4�G@�T�7��ۦ�J�9�!x�!������mv���Ի�����B�t?W�t�[S�eJEW�Y�Ȗ�b���{��`6�.��T�!T��j��P ͑���&<���D9¹UG��o��Ӡ��1�v�Vn�]"^��p�Ix['y67��f�iI - ��J�#/�Wܗ�%aD)ڠ�DpKK�̤�:U6k���ٲ1�R����#�����,�T���*u`
��hidQA�⅖ l%��0�g:��0��X2�=j<Ci՚��(�� ��#�5o�c��4��Ls~gi��(M�Z��ם��'���q���Qt}���S�X�-�xAcc]��W��/n��$k���� �X����"��R��-?�[b ���+=��MZW�E�����ȅܳT`M�]p8M����+Qzz�'�u�'J�f���O���mp����f��/��e;�,^c��u���K�q����2�ڔ�5J/&�)l�GXSo��<�f8⠄�e��/7s��ȌE2<�-n��}6���i�Ф5?)�g�F��F�u?[rã�Yo�yM�� U^�N�hEg�ܠ�,:|�:��m|����,����8ө�2Zt�<�k5�塂��\ظ��"�Ǆ���lX�^��p�?�P�8'����M��x��o�#!�)�O����S$ԟ�#=�����Y*�V��' �_�-6&�ggܧ�����`b4�J9�e��v�0�RY"�*�ج�ՓKODՑ����d�:6S������$u9�Ő�,�����9bV��G!��%�:��!	j~며&:5�v̄|
]ݟ�B!E�v�!*� kf8�t�Y��z���m����<��h:ce��;
����
�?�F�����R\�n�>G6���b����b���N��T�L j��O�����y��5�w��>���	؂$�9Y��Y�i��Ȃ�F7$��B��mC 4%OTEX��|T�`�}cH�Z"�P(��c5��ۈH�����.�k����A%������I
�7s�D�ξ������4\���t|�8b�x�x��*ПDąh��P�^ g��?���y�E޷��D�d�e���F7�O�%ՠ��/��d�Ѫ�p\r��]�w~�����G�qU��?�A=_�̀	K�.�����iZ��?�- W��ۖ�[|#�'���>\�7��,��dمr~B�(ﶩn�2E�\�2�SQ�P�t����GM�Y�2���"e�#�4���ï�>��C���<o�4U��6�&��Wy�`��"1���(�1]"w&`f�1~zS����ݱ�#h:3��Z�.�'<ōM2�ݠuiSRly��ϲ����6��g!Z<����Z$�-0��D�d����u��b�&ܦ7�G�W!���g�Z9���� ��_Z����+�k�δ��S#/Z�~.���P��uS��7Z�q��@mӰ�����`"�+�ί�]K�����A����S\*�Î�*�Ū�7���DcͰ�g;�D$Z+���ew�`;�!>�ّڬnY�Β��<��fu��sj�;�Y:�C�0��ܱ��-4�.w&`�N)��Ǎ~?E�m4o�Ǵjܑ��!�GJ�]kb��CYTf�ػ�Ʀ��b�o�O���8�nϽF١���~a�Y�s���8�;��0˩�y��0+�[B
�@`r|��
S�Q=�/�3']&�}lC���oP���l���^!v� Q�>������dSX�d��#�N�5�ဧ������j��$��@\�0��{:Ş������/~�
[�{�^M/��O�`��E���kvS���!�K���+^��#q5O�f�ٟ�d#�Q���S�R:b�ni�*Y���A�I� ~�b��?i�l��s��!r_��}q
��7v�/�"�9�:�7�~
�6D����W�sF�&���\�~�A���0nO�磻��������a��w��Td���'�m�΋���9T��=6+��P��8�tj� Cdp-�T��!�G\b2����흦{d�Du��{Kj~ͧ1L5�-��~�w��ar�g�0 ٙ^�jO�#�+B2,t����pQ��p�M��p����K'�QB[_~y(K5ʾB�����L�.@jɾp �愠�x9�v5(��0�XM/o�ww�-�%�!�"GX�ʘ'�ʋ��ک�W��\weu;���9��	������*��3̊dm�{V�v�Na���1 ������G����. ��/m���������"�w[lz!�?�E��c���d��>��6#޼L�y����&��/���&�r���f#9��/S}4�^�ɨ?��'���6h3Οf���(:oɲGw���E)}��=��H'��%
��n���ߥw/nM�vI�O��O^�%�g~����"�H�#��v�������Lb�(C~'��,�B����Y��i���Pv»d�D�-i!E"��m��95�l�[Ю���d1>'lS4�KmӇ}`,b��U _�y��,w��s��\�d��SE�,��èDp=����3���HZ���S�\aKm��8m�O�yt�ԯ(���
�wn�I�;E��^@o�}�p�Xg�F�BY0[�_OI+�	���?N�1��M�R��A$����Y<n�~�`�)͠�1D��ı�~i�Peu>�%���\^�#XNm$6���'8d��i0Ìq�7؍%+�sNuMcd8��w�ӷ^r��[�x��y�5��n�3��Բ�	���c�@��e����nP��Г�8 ն�֘����V	fC�hvWL_pe�3��BpmKӚv�.�z��l_[�s���ɮ�Q������00B���#�1y 8�|^�N��D/{I��N��(�D�!�g9#�M�:�!��2db��Y�Z�[Q�75w���.��$w�tF���֏���v���2٣�׸S]b!L�Fp�����now�1ckV9Zi[=Ya9z��R�,�t���Z�xS���?Y;>��NßW��k���}h�P��s!�cJ�h��ؚݹ���$��#G�Ѱ�АQ�K�G�������o�^Iv�l�}�������&&����9�f� �j�U�,�z}�˦� Aʺ�Q��Q3��|���̈�?�6�cHŒ9�Kp��(�g�!���F�������Eg
������L�"���� ��+��P���Wo��2WVp��'/ﳴ��r����$!W�pF�$Z�;����!Wڥe�Y�@�Y�'�B�q���|��&�/'�[ i��$���l�b��*p8��t�LG�F"��O�D�#��0���[Ҥ&�Q��3�=�eϰ��4v�"KY���l��2�1f58J�c���T܂�P+�}�U`��z���:ĉ�� w�M̰
���$�^E��t"��.T?4��d� ���l+�Gi{\[��z�G�a)T�Q�u����mM;�P���_ջ~����A��[���w�09�z�|�,o!Ŕ�Ńќ�*:\H����f=�*��X�j=����'xgjߒ�Nۅ(���N��(^_k"E&��G�0x:q�S��8���#��-!I��K.���
e�����RХ�1(��$N7��;�=W�Q�� 	V�(�j[4Ar��9zt����7�rc�������9��Q穘�_!{J�g��ί��7��Y�6Q�׬��JD�vWoV]K���ѥ���L�?%��O<{��+\�F�vy�����Ԅ%<Yw�)��Po�F婀Ƥ���5�4�5��c\X�0b��Z�ti~L�������3���5L�C���?H�QW�-��"d�#[�?���@�-[m+�Nyn;�!<*m�?�6�:�yie�,OL�V"�\�x)0�-��� �&�z:l�Wpۮ�;�\~�KD�>�h��������t��Wj^a(q�zc�l�ð`��`������>_X���N����bk�.uh��&). �CR�ȔZ �[l�7W ��t,��1>?X�c۬K���qD�m�@��{~�7�,��M�� ���]=DI�_�����sU�e0^q~��W\:{/��(c �m�1� ����v��H���� ��W8ׂB�`_ fc��U�r蟞����>):z؁	���k�]���}B���7��]%����7H����9���]DH��CRl�+�g��iP���9
d�.���.5B)bN͇ x�y�}Z�g8^``Z�� l�唩u����Uځ��t�P�VCg�1)���	�o��>�&`��<��wAy���6,R�q����/�7z�AJ���\� ֯o1qo���੢���d}�}� ������Y�e�u���r$*E��+�O ��U+5�Bg�f?v�1�W�h{!����v�$���L�̪�������7���n~�z�8�^��RW�k/C%D�����|����(Q�@b�Lq�Y���.oK��^��W�8�=}̃�}�gn��>��@i��o��"�(�d@܋�+��ZϬ�����
J��e�b�:��Cڭ�� ��qD��"��_bj��i{�|��X9���"�LPK�Z�W�^�><��s��"ՙk�1�N��T!�Y��Hv�|L�)f�����F0��G瞖.&u��2�~K���O�h�������	�����^$D�T,pҙ_���m���e�lѸ8�m�� A�Ȁ\m�_��������n5z?��I����+3��ճۄp!�V�����=�Hd1�_Ņ<�ѳ��jf<~ʍB9pֲ��j��?f[t�T�b��
��F)�R5�!���6��_U���_Mmt�G˻�