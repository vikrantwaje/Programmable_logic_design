��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?��
��$>��f��"��kΰ�O-�Ϝ%���<�P��;ȵ1��_�N���"k�����u�Ax�l�h���x���7|̡������39�B��븽��96�`C���E�@u7_F�%2������B-*��^�̌x�H���D�������Wp_��y]"�����x^��i̬Pp����5���'H!�j��)3�=�����[L��il���9mnUsc(�#ƇTQ�B|h/�긱��_�n�_^f���?�)=�h�e��Ayj��r{��ӕ�)f�W�J�l��W�1O	�n���,\s\Q�bf�Mt�����%���eH,�?�6/�E�l
��ۭ��2D���>�k�c-�_���s������ �C���{y�n^)1j(W=d9߹T4;,Tاl>]�2+4<9-�|�et�m�R0v�T�ɑ��JN��$�?�tܾ��K`\^��&��vvtJ8d��\0lzL.��-W(��j������=	����7\@��P0�w�5-����?E�?P����2��{�S���P��>k���[����w�'�VJ ��K���j��Y�V����R瘗L�\^���Y;o;��su��	�$e�U�D :��ֹh���O�C*������nKrׯ��~}�TM-�����z�q���3��|�]��J���
����Ё�Vp�耤�-W��ƃ��8��X�Si���=r#r9��!����NN ���9�
������'��uD�Y.Ҟ��6/S����b�g\���I�����8�)%�E�*�[�Z̜(h�jޫ�۔�φR����p5!Y�Z٦��1Sǅ��N>��%ssUW��S&/u��.�b ?/\��~���"�qܽ��'i�t�r�!����ћ[���#�𻟠��S��)��r��r�D���>O9��@���1�E쿅6`��9@5|0��|ec,%0�<+ �L���,��ӓ���n���2����x��_�h�%
sj��������xI���^�Wj��y"��L��jǨ�-���|�]ˀ��p����=�� G9O)!tʦ�"�,��}z�u�#�>P�(tmDeK/8��
�:?yEi��ؼ�B�Pu�n���pN�s/�� �r��c�GV��eCl�x��������!R���t\�j%�bΛ����;x'�o� �[Q\E�zp-RƇFhgW��5�GO2��4��O�M��x�CJ�'�GěƯ�˥�a��b��E��)����W}�M���n��/񤨒�%+]lL�% �F�Q-�K�*���zq��D�ǳX��R�=Il�1.1�H��������|YA�Nw�y��ώ�x̵�4����﫧�k����p�:�9��]��fG���7��|�"Qp�4��6�_��Z+,��5x��S͕�>�� w~����
B���)�i/:_0
}���ܒ��U��\/'����?#�=g~j��eM04�e��|E��>߮���$D�XT��ñK��Mj<�`<�Tyt~p���p�fs�fK�~���==w �߮Ba#݈��������$�.)j��M�	��#�G� 4-ok���+���ZeT�9�0��,J�FT�Y��K��q:\,��L�ni[��C �Z��c��x')|����Y���=� >R9������;SS�B���ԛ̛�>�r��r�B��6��\�Qc{V~�����RCO6�W�w���( ����F¬����"GN�i���Ј�/�e� �6 ���v%��/�]��2_�~	������ʾ �M�y���"�E���Q��}�u�x�:"�{`p�g�a�2��}=oTGK꟰�����<�؛j������\�`k���v�3��r`�>hM��pj�֪��*+MJ��y�� ��'��'!���7�<×K	G7��b�7�G�����Nށ$��8S��GR�J/��T�A��B��6��]`���j�g��+��(�|M�1.�f��B�7d0����*�qo�K�n�22w�q͡~�9#��̸�NK�D
�����J
��eX/�r��*pJ�cw�e�8!ݷ?l����4��p�4��a."�83��l5C����I��kOckp}ذ� �i��Zaj��H��X��^�V�4�>�4)<�I*�/ʆ �n�r:�jU�c�F:�KY(T�8p]��	{p�S��2ak�ge���W����?�(&!a��5���-/�����^�w�:��