��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&��|�Ύ=>D�v������h�O���X�8��������e�F�;�-�JQnK���+�V����ٵ�o���J�������<��W���i"�F���
���t��K�3��R;��U����X���gu#kpA�,ߗ�����Q#c��"�[S+���}�_ݞD���b�H�����0|�
nEb�6�����,p�ѯFwRc��\����n���j��s�Wv�W��������C�8�BJ�.���8Æ\�w:LΈ�}	�*"�b-��l\�=+��Wf�L�� ��[�������hx{i�V��,��z��f�Ӹ�6�Oxeq�@�O,*�� =ؿt"?�̡)Zځˈ�?���=U�����iJp»�';����d��ȅAw_���D��χţu��Рq��^V_�}�c�S2�Q�dZ�ə��Bu�5�Wg-�������Vu}L%/>��`xO9 ��`� իx �{���ڟ�O%����'�q*H���8�В m0�9�Z��F��Ǚ�<=WN�t�Qr�c�z����k/�,�����Q�N{͕� ���ge�0��iW�nsPCh�\`�ý�VaK\w����?�aI�����Æn��l��/���ex�Q����7}�,��`�����A�)iu�f��S��O?�� eF̵�w��f���-gR�$;��&u}�0��@�C��t̨,�'X�PHO�Ln"I�K,�{�
Ȯ��AQ[�|�ܓ�E��q�����U�Zd6�=E�)_�����nU���n��*g��3q�߅;X>ݜ`�Z�e��*����2��曍`m�O��˦?=�
�YS���b`
�p�A�Lc*�XoR��U�⫢*�a_y�a�l2��3�(hIw�􅝗��`z�,Q�`�o}#���i���l,2���3S'�����M��RC�Յ��~��[�DɌ��S�~܌bܷ�T�#���k��c{�������58D��R�x-Zv�,��86�)+,`��X6@��l�9"`��tP��J�͕N��I�� v@����������.�Gy�Q��ě|�:���t��D^��~��k���P������hw�����(��@�@��
r�z��@  ��拌���['ۗ	M��BQX���7g�'�q՚�"=N�����=Rqt"l�%iD�jՍY6Q�r*g���^�ֻb�_O��I/䅱�w�J)��R�wG���n���۫2#9�������u�t��6ͷ�|��d@d���'(�Rhk�9g[u��u�̠��:o�Yf S(?�+h�F.U�g�.�Ld����mw�&Jq�Ү��8��/R#���j�
8����(~�T���>�,|�
��	��ݹ"LgShZh��0� sJeY���Ց�5�(E�����ĺF~�- ��-��b���+�n�Q�A��ͷ,N[��[�R�w�h�S 1�	����/(�wf�/Mb6�MTP�%�)���sqV��鹇X�'m

&L:m>��:J�^�;N{?F�_� ��Ũ�qN�6��d�sQ����a�r�#5��u�&7�͙Y[�0�Iv�2�4�q���\M`��C/��r��qv��RǱ�\:�u(]zz���R�`�ķɆ����������/�t�v�����3N�`����C��5�Y����N�V*���n��Z��Ø�~\����I �-�JU��W��!��?{i�p��DVk��P����Đ�M�g���%ַ�H�`���S\j7^���x^��o[Z�n'��G&|��֛{re8���:�w���� :����R]l��H}/��	��]��7^�����k4�������i�� 劣��JQ�  �Y��V�P�r�⻦~̾M����SP"����ÑdR }l�w����ۇ��Qp�J�H�&��u�!(]%[�����8�6�q�J�(�9�8ѕy���A!$j�Cc�1}�3��`p�i۫Zƫ���H�&`N�a�W��;g1�?��h�@	6S��3>�Ϭ��GLv�z���iz���p���.&�¿�x�mD�Ȋ6�)�{��$�s�s��B,h�����V�|L��	$�5�O�`�̵�,�3��!v86^�T��sB{� o
h�y)�/$�f��ە��M��뒟���;-r:'l�Ze�D˻�W�c��v�y9n6Q_3��c�Z�Z��Y���뇓n7�խ�_����l����;Ԡlh�C����)����Ň�5�鄐�4ה�P����	��(֖4� �Bn*����Bs���jƧ/�)w]=4�qD��--��2Գxom�5�^r�� �p�(�,l);���C���-�< f�v�u�*{#ޯ�|@�2\mC��n�����(���HuL��e߼O�պ�k�w�~u&�<�fC��ի��Ex����cxX?���sB�eƩ���D�P̩�U�����0�׳+#��w����� �`�/�;�=��/���"m JM�=_��"�w��حu�7pԈ���_���)E�G�m�:��
y������w����=i �M"0-��.��a��H+ai�!'�>�&'/�O5l���S�TU�R�U׀�t�D�Vߣv��M�Z&NҏJ�V���X�U³Lq[s�AU�{��>fKi!Bu>lN,��T�(O#̠gR�0p���5(x��ԦC����@��q�j%�qC�=*H�f%�����P�(�b��\8�bU�#u�s����j��d�8ː��_��� ŕ��nN�ZSMi9~]����zç�h�ᄘ.�����;��`VFc?����f'��b���+�L�d `���$	��Wf�H�oG�P�k0hj1m��Dv������|�M����Z�8��#&�5�T	q?�$L�]���
5�k��U��8 p�ɞ��QC/Dk��=yT��J=r�!�ʊ�&hcX�΂����[l����K�n��J�%,����^-�6���h���kx��ٍ����s��P �7�H�����]=[��Ӷn��5a�����������)��������l�g��]���׿�[��s9���>��:A�*�u/�~k����$mi����j[a]�Ko�v�G��*��%\h�)%O:�7�V�Xc�8\�u�(W��}*�D�qRGY��SU�0�G�)�v�_	�T؋K������X�X�խ��vi��I�x洭��e���	+���%@-\�R垑Q�t�E���)^�!�t8
m���m����3$6����q?�t4�,/� ��D�H��X%�̥R#�4K�ǹ�"**S���]�_�,+_ă�
M�m���,�WY>5:��߲!������*����@l
�����J�Ҥ �fw�!qs��i/0ԓV��ꗝq������2	��!9&��z2�c�Mm��/b�H��q�/�����e�Eqۯ��&Tw�[s���+�gʣ�[:ſUz��a��Ì�B.I�+���3�ɮI$��ژk���'�Nr)B
��O��j�4T�����l\�׍�Fʂ�H>N��43�tV��L�I����/�U����JI[��ۥK��k
*��wI0�Ot�3R�ʇ$8�D��E��\�'h	�q�d:�Jp,I�l��m��\U6�c�Mۚ�@Z	%�8~6������A�`\dV����Hu��@���4į���P�H	����]݋�Wy�1��ɶ��4B���4���e��?6b�
�_%�@1�z�򪊉p�J@_�{��a�ѓ�M�ʿq�Ӻ��
�i��W�:	�K��0�$�B��q�'��y��!�	Jt.-�k�)�	\�Co?��	-\s���{�9��=Гg������@Y�dq8v�iX��#3����B<�p�pw�t�S�Vs��Tv-�m�� ��KK����M/�5�e�ʇ�!�r��d��)�j��r�����,m��oρ�E拍Wk��Q��h~	�F7ĩy> �S��/�Q�b�~	����5 �%�����闆���9�K��}(��� Q�B.�e��C��ѹ����z	��'QVM j"|�A���F�k�d���,z�n}�+��V���a׽��L��7���<�
�K�~��֐�&��F�?��V)f���Q,�����
6b�Q��a`���:�_�ʚ�7˯(U��T;}y��	��d����{��Y�v7�~��|u����N|:���/���]Q�K
�l�[3�-@�K�� �<o�\ԼB�4gjK%mT���p�[۬�s�����V �8�2,�l�o����X�ec��Og�*ީH�Bv�@�4,�W{�����Bi��	��x��{a�y��o�+��H�����;ӫ(�����Tθt�̯Y8šѾ䫼���%�<i�6�\���DX�u����s�7	��CП��t/U*�Ggr�v��{R��B��P_BQ��L���!U��j�!���e�ӌZ�:���� ���u�ZO�o0A����g�ƺ][l��l��ir���z��Vn�g�S&�� _�:}�\�:tg�%b4}xj@��|X�QQk�T�,c�p8�DRA��.��gӅ��
dof��&��&3�{`?}(�(m���| f�*�/����yF%�]��]�h�Y�ܮQ	.�lN;��lVE���ԛ��ܻ�G����݄3 ��I�p(x�tPFc ��tJ�rq[�I� ����o�rΕo�(EwEi���A�]�����	w�$軛�^4$Ǐ��b��W����,�;�y)���nZ\ ӻ$�oRn2��Q��p�0Й���L(��Y~4�/�Dm�=S>������IN�u��a�gz��;��um� f�����6T)Cm��ľ���m[վO�� '�� ���mŢ���oN�Y�?����rI�� /�\csP�����+u�.�T�G}{ohv-nPy�D�����o�!�)N��G�Y�;��`Vŉg&�g.?�qr�YQ*T��T�u]'���پ�1c�p��+����
����hg�Qr��
���,��Є�.�;Y������-[�7uEfv����/C�4���3I��W�5/�N��af�b3<��]|g�w��&O���RB׀�d�9h3��(k�J�p#�O��+^s�0KhI��d�o.�C5p[�@���%v
~�/�`�WF�����E��]0l���<@�J���j����u�岖�l�iX�����;$�*&`nu+��&|rPXj���Oƌ:,+2��(�|Đ1ۮ�256Pe4F]�;�{��Ȕ����$,^�iQ�?<���-��5'�ļFȕ�!��	u̒�k� �j�0o�1�UR�?�-�J'gWAF��2ڐs����rj�1/�~'�۴0NwM\�)�Lflt%4a�Lq~(��^�l7��E������Z�p��	�zPy���W�Ɣ�Ί ��P-�W�N*bO���a�ឰ�Gvq%�����I#G=�æ�s�1����9�%��Qrv�|R��Rh���<e(�m�2_N�su�!��y���:{��N]�7b��ڟbܘ��}��;����ن�]	�њ�GW���ɹ�;��d���^�ٵ�C���H'���I���1X��B,��t;��{(��k�D ZC�(OA���BM��â1�4�ٗ�G���M�<�vù�?�}H5�vV@ߏ�^췦 |�Pź`�m��3ɣ�R7��ēVEԘ�����f��mO�.��7�=��[���h���~hM��G;@_���|�����1\YJU|Dy�K~�;�Sj4I������8�ȧ�2�ne/�-{����֕�1>	��zF���
�� *ԑ��Y���{�]Q��1T.g����i�S-T,ɝuOgf]se��B���%m�[��^n���
_$j.��ٵ��@�!hvq���4����P[B�-���b'aZN���&�.������&gJߣ�sǍ��L��Q`���͓t�Y9���ժp�Cw�����ge�|O�Ѥɗ}�H'������q�%/*�:o^j�KU��w�D���h� ����v'{�h��&M�������r�~�?g8��O�4)lK�@z�x���}_CH�����O����x�$�o�ZV~�"Z�h3�v:n\ Ґ�Zv�JI��`��#�O �$]�O�� g��.w�c�:F�P�p�K�$�i
v���-o�$�$u�v��E���K}�O؀(Z`�>��O&��W��l�3E��)����/��t&��9B�f�-Ph]�s�@~��8�f��RAG�5 �>��;]/"�{f���y:��bҪ>�t�'\��c�;��X =}����<�v>�[m���Ѳ�&�J�K!8�^4�+.h���}޳4ivtdn�le�`ܝfbs�]�mM�T���lƪY��U_�H	��^t�jr�N5��w͋�ͫ�|jiVr�M���q�����Ɯ2�:�a�S�V7�oQ`o33� ֫GW~�SlS]Z�
LaF*CI<�wf�HI�H��� \�v�5j�xW�<iu������Q��0�v=G�}rt�{'!�/��V�0�a�(x\4��g�u�,��/DG���D���3r�O�ay�kOӍy�%������X��r����Q�S��my8ҫ�>zk�r�\���X�k���2������?V��� �,�9�?f9_�H�O�ƄT;q��>�X�D٥��o��w��B9o�
��r�7G�׶ΞQ�W\���l���>�U�	���E$�@v�)��̷+���_p���J����z���W�	3=�|V"Hh̦���K.t�l�ۥ+,������G�9�3l�+�3Z�`����
-ENa����"K[�І߄	��#G}�g-��⥕���gd��G�G���3\�V�to���=�uˊ%�'8��z���OXG��b>aН����Ղ[T��؟'z۽��-�J�i����Ǧ���H��Ǩ@{S y�s�~%��T��f��5q
4���m�;K�H��75�ˊӿ�GT@?^�	�<��,�C�E���j<�ʛ;*���N[�2����������T?��\j����OrF���ǔ#�ͤ���_�����y� +/!�h=��b�:p.��Vx��Y���u�9���Ok����ȇq��N=h��F�дFs�cz�E&�Y��&�u�j�9������!�b���ԠDӊXo��S�������Ut5_ {����J��r/�#�wH�������O�U��דey��l�M�č;���T���w��*�-�S�fq*�C��+S��x°�Q�.,#,���cQ?���/:-�ٍh2����L�r�j�~�L��w$6Gm���@ݩ��o9(
nC� /�t�(;Sto;F&�KZ���֤���Ks� �6*�����U>6��ϗ(�p���|�v)�����c��q4�E-5��0�ُg���q=����7�Pj��lM4��BѾ�<*y�Y����f0^���t��Y��m�J�2P���26���gʭ���|�%�^��Xa��&^淜[��_�k���½�i�ڭh�]�(w��S,62$a����Q��,:T��HN��r�ks����T��q?|�%�^	,ͽK��ڄN�� ;�����7��|GA17{-�(�"�F/�A�iH�7!n�	����F�'{���F�������q�W�u}[pR��94����</ld"���(b�ajz�����b�������8������b>/������eo
�ĥ@�~��U�ɒC��4RS����}�Z�^K�G9��F9�����
�������j�R�n�dEA�F�qsyUf��|�<)E��+�G1)�9}T�3'���2t`�I��~X��q�5%��]�G�u�o�<�C]W=CU�p���m�@�_�����^:�~��SL��܁a�yw���U��?�qǬ����JCg��m��0AK�����Z��m���<��@�f;�j��Ю��H�qH�Is����殴�,�s��Z7�u�9o�[��a|C��a��9�е���	 m�}�a�K�e���� 3���H��������HSn7Av6[혳u0d[��g~;�dZ �LI"c���A�Kh�m�+�lp�4of�%�4O��������9X���C�߃�>�æ���n�����u��F�����GZ���\	����N6e���f�~�����S�X�"���H�� ۅ2���x�ݻ�C�A�t{�$�gк���݊K�G���uT���W�,/[�[h2,,%7	�:��O >��0���v�`Wv��涸�$��?$�q�lW������6W����?��Vޫ�|8\�g�W]wGOb�wgq�������F��"��/dQ���䎚m���߫9�Z?ى��?7�U$�/8���6N�[?K8Y@����jm��?ܙ���� 맴�^�SKM�9(.�J#��f��^��� ����X;#�����~U|P���Q�������_�3	��`�"���#>s��~y�a�Ъk����^n�Z�j�{˹H�J�E��z�^A�;�o���q�#�\�F�ئXo0{��&�J��O$Xk-9 sbØ�'G�$7@>�+�὿bOfg�~�ct�6�&(�ǥS���o#���u�`���G�i�]����@K#��>��o��~��q�ʤ��3�'�&��M�8d�f���J��*�Z�a^B��B�EiF����^�J��Ҵf�y_�ݯ#�˜z_�'TeG/�k"k��o�U��)��Jw��
܌�ЃR%��*�����̧f�r�}/8MK�9S��t/�q�L@z���k��u5�\TQ��4n��M<�\&�ՁZ�b��8������D�;_ �},�M�IO2}��\���|��*�BR/P	E!�#J�>f�eQ}�7�"��*��)��_����E��f+��|c�.c�E�F���680���L��o(�pW�wL��
��Q�bLY�$���Ĩ�ғ�5@�����cU�]'&X���$�A8g��&N��!��P�K5���k.��K�z�[q�ܪMj��-b=ot@����W�+@$���T�Z9}�����f(��
��>p�\vPB�U���#�����0�Rph����>��`���5��O�#z�A2��_Gu�x��=������ns��Щ���UB=Ѱs��B�Ps�W��P��OokC�X�QOG*��?7g��"l�^���Ȩ#�)�AE��[_��i��$R�W�>?�ː���Vx��2��PVh-O�\=���5@�>:�'����b���}�� u�r�FLʪP���y�W�VC���~F���T}R.��yW���o�|�ӈ!���8
r,7)��|�����H"��޹ș?+t]�*ylo_{�)o�H��o5�z >Jm�B-� ��Vu͵�m�'TT�B�6Pv$�O��uk��p6g�����^�	�؂k��H�ڑu'h)���2��֒�f$��$��ݏ�B���fO�am���/����w�b��1�$NXS��5,ݧ=�>!�8i������,"vl\�2�N
'@f��/%�.�SR�B���h��]!�9햼j�d�z�@��xc���e��,��R�'%�#@�ↀ�l�����dbG��D��yX�ڗ�H	tO�P�|�?N�4o�ߏ�F�3ꞙ��
3�M�����Ek|9���-4Y�{w��Nm(�7ؑ��2��s���+)j�DO�׎�����r򣝷����q=C>O�p�����bh[BGUt��C�:�9�D=�gq��ά0���F���^�9��7aJ}���̫PnPl��>C'���B_м�[�}���L�����@�>�V-��G�������������;��4�,�g	�3���� ª�D.�7&�b�f�7��ʛ��iS��Maw��20}�H]��������V~��u����B����I�Ѡ1�ϥdh޳����
�Ȱ�F����I��ގ��pW��G�q����5Nj�YHT	���CI,�y�2㕮zS�����S�n��� 	R�&�F�$�H �O�eE|8N�nX��������"G�V>w.ݛچK�s��t�U7�)'�+�U�`�[a�}��O���/T���v�"~IJ�Bc��o�e�_1'dQ+�ϵx��2j�cք�*�`A��I=-�OʌU 
t���i5���wڵ?�+�#%BE庡�_E��
�F������R���N�
+z痐��U�]��>Mܿ�k�g�s��������S#��Y��"�!�>�����ߌ�i0,h�f/t��ń��O�pV�f����Qc���a8��E]�1��
��̯/N��P5�&�1l'�%X�^l*)f5ɋ���OV�>��܏hR�F\�����v��JD�B�x̂��,o��E�(^*�����CgE\��:�Ex�O�+}�"]�<lcޛ|݇D*��Ls��0ҳmq��R�d�y\h��5S��������*�}� /*j"�7;�Wޭ�����iY�̖d��n���0��@+��MN�%�	���w�jQ��yAd��ślK�����	�Dz�~�p���s�D]6;"�j?ϣ���{�%O�4�o-jF�5kTe����P�巖}��,l����Zg��H����+�`��Jj�St�?�+�12
�� �궕����=�Xt��s������)y�^��-6 ȏ;��7�D�{��	����qє��+����R��.#�v6J���T�ǈ0y��<8�.��IWElmyu�W\��b�6{��6����#h�;[&
[� I�V]|��G <w��Uh����.f������r�/1�޳-ĳ�Hc�$�(���1�"
�̥;O/i��"�ܦMoKV;d���:�ׅJ�:C�{�"��ņ9%G���8��<+�����V��}����n�\�9q�K��~[8��s���2��B1���e��m���x����R�y�<�i���pv����0�J���5��Fs�r��@���z�t�kَz.!~�S�y�4>�Q�6��m�]z�7���Ŋ ;:=��j}���*�5�y���1`� �+d�Ѕ�I�:%'����K9~��a�[�x�;rN��e�춇�����k9��<�D�]f���a�9��e���{��OH-��I���SlYH��F��85�.�uQ�k|D_�������Y�_����g1[�@G�����Һ�w��k���m��b籩]ϊ���o��m�aGX�)�U���;� sc�m+#����]!+�	���c������(,�0!~����s�����z�pCZ�l��c`)*��I�+Ә^d�W���Y<$JC�l9&s��A1�\Mak@]'7�}�K[�}����+��Xg�mE�<�5�t?�9�xAOI����:�-�J�X���yWҨ��@㈐�$ {��Bo���%�볡�I�w���<Qm�L��\Y�Z5��_N �<r�?�_*>�����a[	D�p���֜����#wqLf�5o��������c�U�	4FMGH1'fDj�1e��FCu�l����C�j��ale�g�L �^�9��NV#�<6B�-n�L��y��S��4�n����>Ğ����0&�h��k>���3���������	��/��kk���lFt��Uk�G�]�RR� �b��"��^6��-�n�a#%��2{��Q���5���\ �\�Q�q�FU�%
..��FFC�釭'�(#b\�P������d�*���&/��8<5[��I���zо.��H�9iQ�yz��b�:~t�crQ�쳟{M�sGN�Ɩ�#-�0=�����U�ʘ����*nmi�����9�Z3�����bL,S��c��˿9��i��Xc�K��qL�\m��1\.wjڪ[�׏=��Vl��ivse�d*�I��Ꝟ�-�M"ۚ��M�wI�P�ҨN�8���_��(K��5�j�&L���S��T��CW\\�	�`�-��M>s������b6��x�|*�v:������r���@�5�/�Ю	g�u�\����������z]e$u�-�C��>oÜyU�$*�i��Q���۵��Fn ����h�w(aY�'{&Fۯ�N�J�#�H�~�4�����D�nL�'b�Lpgx�!�H�!,2���7�V�as[�K�/�'����X37��	 _����km��@i�;2h�X�_��q>���<���,.|'��|���ӡ�+K�{7�`��P�����/5��~��3C9�
9���� H��%�U�*�.d�#�^���VW�sf��௵;�Ġ�d��6��d�֫�@Iצ�d a]7�����b!���z���<�'�+Na~����%X�f����V���춚��F_컂�ܽ��^q{e�𷅄��nq|����:�sKq������{���p���z �z,ђ<�'3ý��a�(9�rZ9컓�G�W�{]�j�]��E�MS�K.[~��#�$B�j�Gƕ���$O�J �@�/*ڨ��	�V�y�	v��Ԭ.���5�&����V�<;c��Nٺ�u�w���m�*:TW����]�9$�F2�VV�+C���).	�[~�$�%�����i+Yz[�P�m�3E^2����vڴ��4s,<��p��xø���.% !�Jy"���-N�^�%t���SԼ�I��RY�̿����&�7��_�lK�F:�>K�~U��'p���H�cn@�V�$F�#���s�l��f��@lBNB$>2���fպ�_��Y$�����bڔ��~!.��ѯ&�Vj�d�r=��Gd������a�����|�*�G�P��E��*i����$G��$c�0��<�_�jR/ϻ�$�?p��&8�6��u�c�Ӌ:�b� �	���L��%��a#�����ɧ�T�CG���F!{P�9�f>.+W]��/���:|�]�,d:ֺ�8F���\Y ��{|'�ҐC�n_��>C�/�Ȍ{WH�~�!b�,P���`�K=��w�|���hC��n�N2cx�
1�p�h����z���s��dr��G��N,���1���y7����+y�.��x;{7T4��@��7�j���0g���	�u}�/P;�E�>(�����Ɉ�^��d�-��ٙ�0���
;��a�;�o��#�����/�Rq���d�
{���|��#A�l-�Cٱ1t��`��+!����	���ک���v8ۚ(տ�3�L�-�;�NB�1(��v]���ꕕ��o��m�영h�UC+!f��^>V ځ4$���3 3�iL�ey�:ܙb�,R�UQ��W��?�>^ޤp��j+�S6y�>p
����nU�z�g��Ť`�nw�@���ԐU����d Q�y|H�^˂������*�Qߧ��ƕf�m?!l�� w�������q}3z�P���
���ѹ�1�������ce41�W;[ �&�+�W�k%:��V�;|��R������Ƅ�K��Ž�]���[�P�*T�_Q�G�Msb7�lzy��r���������>_�VA�g		�yE�G:���>6����)̀�8̡O�@�!|�;(%�{�};;��=�;�<�d��&U�}���F~�.�tNw���:�<`�˧���	�BϿ涊�'�|DGp���q>�|{�Jy-�O�����NS����������|���׌��Ί�qz��C��^u�+�#�	8?cIα�4�xY�x\H�U=��=�h�O[R%$44���zۿ�E�Z���Ȁ/�L��:`˕̓��I�9����CO ��tH���`	�GTGG)�Qf�Z���@P� �C9%g��x������>Aw*�	WV2"�w"�Xm�鿓Vg����WR�����"�y�G��V�t�m��y�&1ém��쯁d�L�}P] .�6��h���XyL����FS�g43[g�/c]�=����|r'׸P��j���F��£^�w]���!���vb�&�Dߣgw�2:���8pK���0{�A.a�EHy���pf�Ӻ�Ls���:r��z��ʰ�aW�Fei�R,v���yt�ؖw<�خo�U��||Y�����|XO�$7���9�����Pc��Gf����2���5�g�(rӟ&���
}1��x1`a�|Z/��ܴ���b�%�NY�ږ��'���?�h�9�]X{YU�
�az�{� �O�M}���'T���.�
toe�o�D��#�o�(���f��Čz
��_��9.O4���CW1�D���/����P� b7F	w���G_1.#/|b&G�8~�/���^s>Q�y7Sa��,Y9?�"@��#�TW�G�ѺX�����K��^rȝ!*�LGEU%2�AM�Ͳ>�j���`�^~|���3C�D���N���ѫhc$��g�"���$9��?/-�;����I[x07w�TN�	]�u��Z��bWX�o!/m�|�o��/��$��n#�9H.�;qw*���w���?VR��?�~�A��P��Ak��H�r0{'6�"�঄�J�<N��AujYh��T[�V�>ww�^Af2H�+6�>
Z��E" ;�k�b��#���)�;,-Je����e�&m��/�����_	��*����a����7��	A�13p#h�Tc%�!MAR�y�.Ơ�D;��eW�pi�`����:"Z�ϝZ=7�o� ު�%`��	��J���cs��pn�\��Gs)Q�Zh˞E+�D:��N��Ɍ�F�4��[����]t��k\��y��`3S �s:'�gyC0�yR�5J6�y�[�
iĽ2?��ٷ��Y���ی��z<w� �V�����>���x�U��8�x�-H���Tg���P���-�9i�t
bl�S"�)H.�3���S��؜�����r�GQ���	�N�׌K���[%=���;B�So��7Sۖ}s,�>�5�>0ߨ�ʝ�G&�>&��3�]iA5?�~�A�&?�8"���L��O���<O"�h�+bp�R1�psQF�5ɞ�I>K#icH�������0%����ɶ�#�������{�q�}~�J@b̻!�+�q�c�&��)�Z�4�V��G-�h�py0�@���b�@���}";��mʊ��0��>��G7���?�]'c����-��H�����Dy�G��`%���,���k��+��ކR�������)5)�s�,J���m�8t����D���o�i/Y�ʩF����o��9;%�� :��D9��y>3b*�l�s��ܕ�<	�?��Q����7ƨ{5Z��c,w�pC����]�\���4����LXv�����ɍ����nd%C:i��6�?��
��@,��?��~ ��D����o�0s���bR�8`/��R#$����Θ�ܻ��m�.��K���O��S��|�K�k�"��zm7N���khN۾��TY�p�'��3n�l�axKb)��H}��D�8w�	��¹��F����Pz���e]����K�B�2w׎v�V����Z5sIza�R��mPv4��Q�H;��!����n]�˷\˄��JS��\���fJ#�ܦ�eq���@�"^�0��+d	��`v�@�qǻ�N�F9�oX����Dc�S�X0��}f�&P�rC1���Tg�Z����'D��X��,��,1��L�����((�am�����X��U12y���8��"��3Z50����mF��[�H1�H7���I��Zm pv�}�D�&��+�8�K������i&ĳm%�M�/x�3���VV6S�R��ۺ7}a���4�@���<'��'�x�ZKش�M8"��<��3�6��p�����+�+1;կ5E�*L12�'�X�idS���~6�a�č8q�����`�xc�Tg��ݻNdv���q�ѹ�)e�噄wzN���5.4�;%z��P,��/�kB'�k���ˡ�s1����2�g�2��>1�2T1v��4�L������CB1�� Ա�ED��^�񤦙 � �V��@C������p���X��`��og�eRݤ�G׹N)��/���{! ��^�2��,d����h�~<�{��#(���|�@L��Hl�N��������g�	]�O�+u��U`�m�w��R��ՓrNO�~C0�f��ʩ���9}�XߜO��]���L�X�X`�`�关���B����q�>�$c%zH�9~Z�j������<��|��&��5��M���mE��P?�/��H��L��ש5�F��g��3Ѫ>��L^�͉��j����n�^����h��r����m��+񞇀���B>m,�K�>����~��٭�qS*��X%��I��c�om��%�T�z�����M�n�9tlnUυ�b8ALe���~E'�dY�fM6m�a�)�Nm��<q9��y,%���fr�5���?�71�fk�/���o�������U��ՠ-�6|����.!uGy^T=(�r����{|4؃$��f�)MX����c�!:�I#`�=����pK�S����������y	j�<G~"/�
��㦫½�Xt���)�����Sß��׎�nK�Ք�6��֟�tV|c�;�W�yg���U�6uG��dI�	m8�@
��E=��|�L��ԗ�3<�U#:�F�#[��*�n��9`�=��N=��_!6�w����VB@��x����ЅD�lC� ��)q�f�^K?��>#G��� ���C���tY!h.��	ۄى�>c��D���7���Ұ8����P_:(�?T����-x��P���k�����>@X�nk��k��=)m�J��O2b�;�Z�Q������0]�����Re��.� t�XlH�IC��ԏ ���~�u	+�g�}���:5�ѶZs���ur�)�<�܈Ѫ�Z,�<��B�US�����+<�~Hj�$�&A`>e��7��8�Mx���6o�ܭ�j�ҏ��ۼT����p�s�^p��$@f����e���@	���(W�1-����ڶ��0Q��(~�ܐ�N"`h�����v3�>ꦻ��2�m�t��z����lu-R�����&]yۡ@��)]���b�Q���\tM���d�lWv�fܤ�.�&�kC���'�e��D)c�������C����e�f�ap���'�C?P�2��]<�W*��V�H�h��776��K@��ZU�*�·�_��G�M�Ճ(�T��)S�׃;q��`P,�̧�\�����iXLȮ��`M���%�KJ�
����x�z��V���a)t�LZ� ��bdQ�&���ɜ�����{�Mz`�����D�ޡ@F� W�p-_����=�|��]��i$ܕ,�q�߲c7Z��E/y�둲)D}�����Trw��$��0�P�#Z�L��ɤr�։�F\��D���&*6@H5��I<.�����n*��a�ȃ�ŵ�/�VNa
��߱��=��J�e{��ֲ��{�� F���*.ў��ti&h������T�;8<�{��CH>ñ�<[�vX��/�$�@{�,;���<��u�X�h���vegM�})���	�bx5����tW��$�(��M��3<���/	+<�<_�P�ұ�ύ��EpTtxΞ�d��fv��I���C�-�/5�(���A�4�R�~��=�6ۓ�^~5�5��3;�%���9�"�3X��W xW Sl�G��.3�"���W�.#?�'H��mR�b�#Q4�-���Q:$�^P���b���n�g�Z�0Lc�1S�~"��L檾<�%��i�<���[N��h��Ӡw�h��e�F��І^Ie�-�.75H�{U�1�~�!;���Ŋ�5D��;���?x��a��x���s��i`�o�f����G>�u�d�W�����)G�{4�)m�l-�nL��_���a�����\�H�=�8�C�0;�*By����Y�C7��U�q��3�Z��P�}�������6-�����~�v��o���XW�Z>��w��4��\qG�[���3;��2��é�7T*_���ho`ܤ��q�ڗ�V�����3h���W�v��|ް�`���9߆�Y��7y��`"~ٯ���vೕ��lG�{Ŋk�Iu� T�x����$��7BF�)L.��f�;���h��sE��_�S�bu�<K�����p�0`�Lӓ-sKĈ��n�25u�;o�h1yf]�5kG��s�B^��b��#�FQ-	��!�#A�x^˨��T�H��'P����i�[��9��Ai�@_kO��D�g{�Ɓ��^Floۨi^<�Ʊ�9πq#5��ҥl�{�0�T�]n��ʈĽ񘵐�˳���kBW���U9���9�*��Ͻ!��q&�k�~��n�B�m��c�1���˭�w�;>q���ƝR���}&��	�Ak��nD4n�����r�1Z��Zʁ�@�m�E2���Vg���޽.x�z�F%Z��˄(,)@�T� �xX��`�'�|_������ĉ7�u��V0�C}����Gp��I�	�Q�M��T��h�NU�:*`�6HFgyo�/�İ��Z�tC�7w:�D�#��B���[K.ړ'C����\�k�7�燦�������f�wqΟ���>�r	��ʟ�"�C�C�|�!���� B�v����BeD��=b�Nv孽iF<28�����2��z��H;|U&-��2��w�"S�����i�ɿM0q�Q~���H���\���k��_6�V�OPׇ���Ί��3����"��t}��K>9�����j��/z��M*#D�s�ӆ9c���KS��yo�b� �]�k��:h>�!�~��wb��-�:��$��k���������2�f�`�A�訽\x�7��n��h_tu
�:��Ϡ��/��5ay�q-G��	HTdV/�����.]�ۍ*ڵY�_�u���ih�Z/�p\�t�A�*Z�����^Nrx-Sb��L���F��Z� ��v�?����T&�����ũi{sД^����i+>�sQ8����sZ8#�4j�[I[����g�������f �!@~��j^g��tݎ�qf����m�lo�0�L���bH<E1P@�R=��yk�]�4 ��)�O�����J@Vqsϫ�Q@�"K������4�gm{��B��ٙ�ݞ���š9�P��?�h"��"�	���}������֓d��~�us����������(Ywǥ4J.����H�ս�@�O����r9��b��LdkK*� HS9��bi�Μ�eo�7|3v6ΛO��\����<�8��������s|������I�S0	�@>`Iel6�	����f�,�}>򉪣�Ρ9�n�_�k����0|��h%�#��۰�z?$�)n��m�Vh!��e�FՓ'��)���2_���v�$�������s3�J+��:̗'�w9�	��e:���y9x+�z�����"R`�/���$����4P:�Wn�d�%�nc����Y�E�r�(���"���X���#�;&��ONB&vw�z�P�l�:=�c���d���E��'&�xA%���o9�V:8�����_�w���$	ٽ77�GY��c�������u�ƅ_��c�);�����g���׬�N+�X�I�m�H�g�4��\���alZ�k���)ts��$�tKj����I����J�L�Wg,���(l ����	��;�`+�?A׽`5��'Tv�b��6O���8��HuA9�`�o03 ���I���2�JX{�r]�h���{ݱݢ�5�۴��$��m<}���;�a�;���ʧ��ʆ���]X�e#�Ͱ��B��C�.�d���J�y�gk���1��.Ψ�:�2,#a�߉ýp�g~T��{)�ѻ� �mh�pV���5<Ǫ7���j�R2�,$��gX�m_�c姼�_	vs��NE���H�"��V(��_
rO;�d\�=�;Lvq��{;���`R�@�/OZ!L�S� G�)6�vO^�V�Vl	��k�6�I4k*��sɡ8Qg��)ϙ5��~X�f'\U���L���\*�p�?"�U� B|�J�ҝ6����� �N|���C+d�팼fy��YC,����s���Ԫ^M�NI ���L�@��Ǥ���;�YEJ�fKq��+���-4����wA����pC��=BȌ��^�F^�m��d`��\rT{,���>��~0�
g�x�`R��e�	���o��'�ߝM�=6M�+X�N��ai��E�FӠވLT���������O! h�^��U����g�vl� 7`���s7�����r2q�C�?ĻK�d-����&���u�R�A`�o��2���7|f��ܤ����{����9��܂�2�f��Z*�P�|]���Jt�K�9�
�iq���N�~A�-T����5������U���S�b(^xR/�U�['3�,u�j "X��"U��:g��߀
o�_ؖ!��p(3K"X"e�W�O,|� ������?�����R��D(Ԉ���o��$VG邐��m=/�)R�s�����=�%�F`��k�'�У�E~��h�T�ŭp��U�֛�y�����z$E'�Ń�m���;~d�1yv�:�����{U5��;�(2�G�C�.����{�%;��W�`�
E3w�4��K�wo�k��G�WWx"�{P�&�8�q����U�㒣�A���?`P�Գ��K�]��v��ǭT��E��y��������rgo�G"������t�~�T H�$B{ھ�sj��m�ۇ�JMLY��bH�H�8�
�wj�4�,[�2�KѤ۬r�.`��C�޽V�x��Ruq�ƈqiK	�^�'� ��ީ(� =�{�d��~�jg��t��F�N����WZLdD
[�}BwW6 %g�W(l����f-� ��	�����;d5��Js%`8����|\�>��0]D���1�#�9��d5"�sec�e�!J�+���{�&)&�~�����mn���A���a|zKN�
�ix|��^F"��Nu�m(	�ّ.i/���W��b�m��3�{d�9K9�p���@^�H��!���[�5ΞQ1fi��Z,���]B�[��DI��D���5���,�a�8���΃��dJ�q��N��8��<����\ޑ���
c���W���l�R>a�eC�1&gc0E��*H��!8��&�{��:���;q_��#s�H��1�=-D��i�FY�$��4�8c�(��z���/�x�$ ��{���7{bϠC,��$r���3�Af�4��=����#1��RYg������Z�k�����d���~5an��_�!��x5D�8"�B�W���ɓ����r�$(9�}�1X�?H����u��h�d��x^q�b�b�b�9\�*�y@�]d�����ȉʆ�~���w�ZE?i�ú@3z�/��H�q-<<�M��Y2:�\�P��cHpR�WB�4��&ݟqZ����ń���Q�|������J��0�"�_Uſ�P��"��~�%��#֥�9��� �P�q�i-�9"��x�v�i�����ˊ�(��ҴY��dHhQ��<a�/�G��Փh���Qӌ��يh��4�j�i,Y����\ p+`��5�di�#Cqt��Y�L�ԣ�t0f�}�|��Fʍ�C8[�S� �KlӨ7}�[�^�MU.{�$+�qt��q[���uP;W�V ����5�0�byoa����V74�(D�L��E�}"����(�e��'8�s\D�����t[���)���l��LF������E