��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛�����ҩv�[r�H�b���x���������yU��߼��FKw��Td>	����5�3hH��������W���I��(��}�7V��J�?`�,Fа �F��YV��b	 ���5��G��r>`��)��]�jϞ�3=��sa�O;�qH������!mi�����d��������DM�:$y�����{PeC;�PϤ�l�X�%���B�����$9��V���0Æ�"�Z"G���ؠ�x�� N�)��_]&���9
ynX�k�͍�f�/M��~�.?�C�>6�-��V��u)ͩ�#���  ��a>(w 8����
s���
���R���<��I��5��Ū��Hwh[8�n,tğ/��9��w�����!$���^��@����,_*�w��+o�V���vǙ����/Ϋm�h�0��E�k7][ddqt	��J�|�mB���)��?F�`�I +��s�$;� ����(�X�����/�{E�mu�^����!�Dɳ�IwlO+�$�\t\g�*�-:�Z_��JއT���D\Gݣ~�q��_�#��F�$�فE��j\NP��R�l_�P���(M�`�
�+���x�}֡b��d�����Ӝp,W����*�l�Wi��.��c�܏��a���6]��v(t�͖�C�%ʚ��]���l�je�_|�pY5�]Ƈ��
��l)-P��z<1�Ԥ����!�U�q�ЅM�R�f���5��r���j%SL�J����V�"Q�=��e1p�d�݁���A�N�� ?T"A�Q������}�����s���U�@�a��k;�R��Z��g�t�s�V�0R&׎��۟K����mq�i���n(�z c�^�$�2�,as3$剴j2\��{�-�M��}�R�Qvg���_ڬ�%����r�6�C&�����9*���X_���زU��)/���1M�.��mL9�/ם���Ш?zͼ�(LI����y<w�5?VO^6��2�/�AnG�qthb=�s�=x0��u�-�T���O�����@%y�#��i'����{�x��M�����Ӊ��a��:���)�u|o;8��c��l@W�C37��[��%�wS��^�Ep�$ФG����M�����H�:y�e���7�x���16pol��_u5�[%��?ץ�
�σ,�"ڛThw���%�ȱ�g�J^��O�����D�I�d<���U��݁���N1uC�7\�R��^���̎��j�_����;S��J�;2�x����jB�1�lq>͔�i����F���b����[�ׇ���NS$��縉�+��@!�J���?~i6�ֻ��������R
�� �6 &����HC���~ɫkgk���K@y�!�����m� ����V��|�/���4͏L,�5�׀޵��S+��W�����T%��<YnZBQ2�S.�� r�%E�����7Hyf'�e����%��h���p�j�b񴴜�?1�T�Ui�s�x�EeFI
nW�yA���\�ZSG D�==���{��Ǣ�䇜�ho^V0��oo�*E��X��7R�~S/[����� ��Oy��tp�-�<���!�-�|���<&L
�����ve��4�2��L���n�F��[��iB�38=`��u�'�sx{%x�6`l1�MK`.��V�7��u�z+vS�]����1>ig��:5�0z�=��xK	�W�M_��k.�W����ߎ� [��t*Y�̒V�bBN�*y��lE>�����mˉZ	���46D���v�����sU��uz��b|�J�?FH��� �ܓ��vo��� V�2E0[��V���yNYBL��OEt+�٦����+g��ξG�a����yĹm�uK�wN�TYQ��s�ݵ����ul�f��'K�ݤI	�v�1*�}�������D�G&���:8�r��7����@���%�ec^�4���$l累�J�:剕1�%��m�>�>Y������D�,`����Tzg�rhF��0#��3
�Q�2�N��CJ��2�}�(�E"�ȹI�V`\���=��q��>!�r\�V�	�b�ck�`�!c-�����w�P�_*OQ�Ȅ�"L��$�xȚ/��$!�'V�ղ�
��6�B�u�`�!?�P�̺y��;U������,��a��~���dn�Q}�AIbG:{�D%�O�u�ZPP���t�V�<�jB�"�
���YG����=�{�O�o�c5�ǰ��/�]���Y>��w�BS�l��W�@#�E�bc�7�C]*�	o#��
�@�wQ�7�H��e����OÎ[f'���[1p�~!���o�WXL��!f.K0���W�`	x֒��`-���!��4��Wau9���u��?B�U��יq-�(k� }��Oh�|���������� �?�����R�Xf煁�/�W� �B5-��غ�Wf��]�=˶��Vn�f�Kw��W���!����Kǩ����\�����Ⱥ!|_y���o1�Rt��Ua��v<��E�b�<�ܔ;��JX�rvV\<�!n�6|��Iu�:�bݶ��t��BsMg���ag~�q�㈕rz��u�[��6�q�=UT��_��~�~Z�mK�i�1��� ȗ��[�逊�Y&�R�lY��Z��t�P�u�A��������s�|�� �C����{`~S0 LiX���Z���_�0�b����}�d"F��#����B㿣������|��<9jV�
�!p����n��Ѯ�`>7�����ܷ��ܮN��7ex���Z�p���L
�E}�|�e����6��e>]?��j;uwJ^ʮ�̫���08�h������ƿ�u�yu���N���Q��cR�78�֎�&�g5�c�*�B��9۳��|����+�goV߷D������T~�!�j3�5I��	c�"��w�
���!�'�r;�(��g�U~p+��V�S����и���W,�gި��Eë���,��WsXʙ�6nW�*�U1>�w$�D���~d�@��g~��al�~��Q`�@�y�@��1R�1B�	��`AT�� �h�]ga���Nv}��g�ނ���B��jֿD�Ia�}>�a�?���C�UrN�d�Qx��?����8���\�}I\Uņ,%��Fgv2��O$GI�F�Vm�M,EQ�t������jnZx�kB֎�.)��V����/��}�M��d�bT�Ҥè�5y�SE��5�v%��u�����OJ�dis�Lu�f�4� dz/P�r�h�s�V���-:!�kV���U��⠕�H���<��gz�̕,C�� Fd0�>|dv�6�HOwB.�5d'G ]�э�F'��S �#��K|B2t�Q���?��V�:��Bk�;<��ff�7HJ�}�'��ҙ�C ҈�ῧ�pw�Q$)��J��sXƏ�[���S��&q�g+I�f�_�˝�GO�%!X-��������QS���%��	ĦYݸ�z��v�D"~鶞���Fk$Y�{hO��Ąv�jz�hM`ek�����w��o"͜��E�z��<���Wx�Ҳ�$�<B�g���S��?�I�X�k�s����9j0��}c��� :���W-�h������9�r�k�B)��|�b��Σ)�Yҕ0��,�ʔaɆ�~>��֜ ��$HK����?����l�A���F1ɐ!A��FS/p�u>��A�[����6��3j�ï
�E��t��Omĭ����Z�7e�W�-��/<~{_k{X,�Eˬ���yf� �x�?�=�K��XS����{�87V�����3)M��i
a�����VZ	�9%c�tι9�/��쀖^i��w؄�~Ky��4=)�UT�#��1�v+[~D�g��Z�$����V���"Q>���8>�J�lb^MXz�͞M��[�'a�W;����=�0*J���v��T��q�����e��Vr�E��쬼M,�Z��<d����0�0�\�V��%�!�`��;��^��=Z_�p��J*5 �/�@�?�}� ض�N���(:��G%~{�oI�!�"��'��������7C<���~�<��zc
���#B����[�9��}�X�Ť�-�6B^�&�����7�Dn\�ªh/!�؉$������DV>�P>c�?�O�ش֞�9^:3LGqf��F���0�eӓ�`&��2���[7�ʂ>���5ۤ���=���3}8s�p�w�i�C��l�ܕ�W`�����Br����2���,��Pn��FVl܅�qva����G���_���_¥�H�X(;���n.����Jc�S<Hߪ�C<��rO�)����i�Q��bf��h����,�Q#�Rc�ߟ��JQ��	����n4قe��\�"c��΄_��ef*��LPN'�F�:{!Ha�Wy n�Ξ�l�}�gW܄})$㻛?B�D��Baw��0j�!�
�����[�����Wvn�e����������г��+���皥0�'(-�g�иv�Xf�d6dZVQ��2���$��;��O�����p�B3�Վ�\�[��w��Ӣ�*�7���\Q�%`U�&6����ٝ��VS��ﴟ0����N��� �Q�T��`����P���,\���T���BĴ;L"�Vg��ؾK��/����u;ԈU^N?Qӱ%mT����A�+��4�_��5;I���u�<컗=�Զ�gQ߸#E��gb����������1�%W2o�t3ڏ�?AW56���M
�m$j��֪��r$4	�|��<����wY!�����;GG�i� ���������`a�eZ�TA$lի&��*��� T���ZH)��Uep�:��\ܽ�&�8q!b:s$�::�AFN$�Dw���v���/�3T��L�S�!Z�K� g��ǐ�y��1�����OL��Ykm[ή�������i�x�H'�!�s̜W��@%}���Bc1��F��mC�U�袅�)�.�J����ۗ�������s|D���}<�*��޶%\/	�Fu������k>���-�A��׺���f���9Q��>�+Gl t(��[�`&��5㯦�]����%~@
ݕ����,�O�&~i?~��y	Χ�:n� ؍�=n�]G��4��U���KN�z���y��7��!i�6�H�3u��b��������?�4?DĎ���h%��ZX�+�4�g|��;vk�6M\���do�Nu�I�����❬����[�G���L�!��ͳ�W�c�q�Y�1=R c���[���Uj��sK�,�o�]o��mh�trvչ
�E���g)�R2B��N�_���k�5ݯqXՉQ���zf�|�Vx���e�j�?L\vU�W��ć�U�T.?Q�`������o`~�No�3&*\Y}h�f;X�(k�Z��,v��u�
����S@�<KZ��U�+�h��F6Zڑ~��@f/ %(:����8y�:�^h͞�*8e��Z"+0����O8dof����2��8 �U��2�ܵ^�rn~�ګ.E�!�^G;��&�ib���9:{y�gOR�������ʅa��b�bh��c8h�dj
,�Ɯ����}jN��V��)#��|#��4�V�T�J��^?-X���W?�0侎vC�K$豐xr��51�$�.2�X�$�rsf�����5k&���5�z���Bl>2�:�6uU�Y�%�r��1�Z�HH���.|�����	9�R��,6�O���m��cO�잩����el>i* `xi�/�ոr�c��K�����Ђpu�hQ�f��txM*(�y���}bݙ�����1B�颬\1* :�+���)���uR�g�ߟ�ͺ��7 �$�UW^��y�"NW�����`_�� �kmsL6�\+�sr�
U�����\�C�H��_��%�&�B�B�b�g�Nhi1U9~E��ܜ���b�BY�,:mӑy�;لxKۓUNA
?��o{ȶLW���p:b��M�-��{�s��%���3�
)�+�Oq���~����)S!�Ba�)��C<�p���f�C�!a�vr������4%Dk4�i<����{˟<K��R5r�΄�gt0���;�Y#"���C���9#�9��kO�QqN�T�����R��?��K�D+����3�=�Y���+��C��R��o+�&��'��32Y"K�(5LJ2ڬ��gī@r����g�Գ���.�uq�J�ќ���(�b���k��!h�9�*i���
�D�N��t���bUO�ǐ��*�;;�'u���{Mx��^i-�}�����V��k��q���e���R��wS"�r�qÔu�D��"�.!i�����D�ĽUO����RA��P�<��=��,X�~q%=�*eS.�����G��wuG�2J�/�OX� ���5��E���=&ܩ�	K�~�#5M�E��d�D�8�����A�X�{m4E��74����*<Q�(��ǖ���A�%4�$E���M>
A; ��_|⮗:����)jţ�y�&���߻yc��E�-���A[?���g7��fԴP;  ��8�΄n_���`Ic��ߴ���aT����L��"������>0�}�jaN8VYi)���Ҋ��u�C�;\&w�����x٦��<� �c~�T���D�O�ĊrӘ�E8^�׫�?��Ds�4���9`-Vx�����#��!H���)^��;� ��k���� ��vҊ��<h��w�����%�l�s��DU��I�B��+����ΎD��6�>!S+@�I���� �0��.�>.�4���*�,M�|�󭮧���\=-:�5��ޙ8�w J*/�	�Ä։ޢ���TQe+�_�{h�S
�M���d�^�I��/N	�k�G�6��/N�����|ʗF,�Õ�8�x�����D󪨆y�A�.�wh�*��EP�+��75�[�3
yي	�|1�)f �+^����ߎ?�Nk��(7�r�����
}c4�g��`Nn%�,ܫw��ݺ��5�;�v"��2{�͡?�y��_���:Y�ߏ��<�}C�(x��A`0c� �(��{��vm���G@����1 �pzkK�@CIB#ϘT��e�<�&���5X�[� ���5]�miV��E�f�^a�eyg������t�t~7��}����H�?�ӄ^�K��[��:YD��n��خ��?�����e��9�PJu��'��ޕ��=HB�sJ,>���O�c<X�'��_��r���:rk�<�UкI��8f�1�{����H� ���x�ګeϚO���	�&aҬ������õ̕��0u���pX�zl>��◖!\ſ��(�{���)��X������m��a��&EUR5�u�s�30 ���� �|��}|��9���]ʼ��X�#�6I�!��d'�%���c"~�ƎQ�kcM-M)eٳjJ*&]��
��X�2%du�@��x�]I���l,����K��X 7�xoA�7������2�h=�w���;3�0���-�t��$�߯��<�#V�:ߋQҙ�5��j��Ԁ�
`�3�H�����<�o����I`��U=�L�f��H��Rׇ���$���3�ZH=����=���:�gƲ�LP��k����,�~r�l*\�{��͗��u��6�a��r};�Q3�Z�m�]%��o=�;�6�0f�����i��ӓ��_G��|�,�Nx�2�=9�4j6�=�����>���@����Lm*�:cS>�pW�����n!+Q��=�e�pt ���d#�ӝ�ƙ+�Foͯ�8V��'���v43����1�%э��r�i�];�٭&�W���Hg<G��fH��@��M��O�+	.��!��d>{��gVTs&��Q6g[���I�K���W���Tr�n"d���JY�=E�v��<~�E/#u�[�c�UY=�%��@4)�F�R�oB��,��T���R\ΰ����n9�	W�e�ˌȨMl(ľ�`�`�ͩ�% ����^����C;������K����݋ڷ��C�r�C�}�8��K����oK6�|�.i"�f�� a��1�y��3�,O�`=�]�����_�[�v�㔤
]��p��-�%��ڌ�U���D/�Un��T�y�瘍��٭G ���v����7s��,�xn#PK}����'�0� � .��\;|����թ�����a��S�1�H��3m,N�Z��pwcB�BW�"g"���$v�3�x�%e�@�r:-%�|�:����+��y�zUH�Ƈ�C(�uN�U�9�F/=,jl��
JDB���^.b!���oÙ�ۦNՓv�DL��v}�is4�٧^��{��!���Ց^���|�.fwoE੼iX-��\��c�H��l�(�\�����%=3�B�a�7( ���@jΘ:�@�����2��/d%�������F ���C�������Y(�oI�{����I:�w��VL ��W����4��|ǍD�̈�\zBf�0Ҷ�Q�f��-����^a\
Қ������H])���+:z��$]'s��50Q�6-����Wo�zi5��̃���y2ֳ����Q��H@�׽�� mbAR���w>DbZZX�Ѽ?=���p�	���F��aN�������p;��af�f��A@:G��52˱���/���I�~I%�B��w!�=o%=�p��˹$6��oE�{l�1��C�M��&|CaI�D��~j��k=����?���AN^J�����N�<� �Pp���eݜ㍎HR�ҤIN�ͪ�4���i�/Dj�K���6#�^� <�~К���-���rc��6=Ȧ� ���[��}�t���!�5�����.��bџ�?��Ɵ�FF�ʰ��\6��:��+F��ɧ��ꌀ��@�vզ��i*���hVM]��Y����׃z|u�?��x?�q��ժ�]�ޚ�b��87D���5�\�F�q�!�`�f���:��4�:X�;!�����*���a��D3��	)��nL̈́�Mj�h���pd,I�&:;��j��3�aC]R��xd�B�)�0�; �	�L�K����`�~E0?#��LBL�Iw��>�q<N'8c1-o����op��ۅ/i�CdX>�폍� jNy�<V�pX�8~�f#�1�T� �p�rI�s�K��� 8��)A�*����qAWB7f�!80��c#���*jb6�R=��y(Pω���>\͕�ĳ^�!H�@���Ś]6�as6�L�W�N'���'ap��#�Ix�-�ܐ.�����O6<��j;0�F�{v��CB��%8EՐV����5�()̲�X	�ɧxs��~I8�Q$��gHi��~g�����&E#'��ぬSY�_.�_��8�U?aai��'�u����n��U*|�jE�?��#|ۏ䢢1[_�������Tj�?2w�Q�-Qa�ʍ��S�7�'3mA=�T^��d%e�i����� Q��ZA�HU�q�I�D��k�v��}0|B��c��a���`�Jl�;��q�_�n�t_NƠ��[���==~�}��Zs-	�����sK0�B�Vlz�?I�ݹV�tM�m j���'��s>�0}�r���\S���������7�]S��*m���\i;�h:��|uv�F=$J/v�(W%����<��<�2�~�H����j��m��8C�|]�RKy!?p���� ���(���j��/Y[,4=%�k����m�Pk��06�KQ��N���\-*�J��{kA��V�#�=:�Ф_d-4�FS����}8᳦�q�^��x&<ʠ��=DH�X�E�AFG�t,|X�8X�?6j�I��t�2��a1�jd-�_M���%`P��&���{D�. F�8��)\r�����B_�,���V����s�A��KF��iE�Y�1r�u��n�(@�����d��ڑ���΍#��I�,�Lpt�������m_�w�D5+�Jk&�;x����o
q�#����"ִ�;�O�V��[)����p�TQꞳI��s�ކ�/ ,U�w<�m��Є,�]�m?ڏ��u� �c���nJt�J����&D�
̕�����Y��:���-��A{?[�G[x��m_�8�KWngY�b�&;�yU��"���}7�<��E�:VUU�����s�a����]j���hL�l~�'6�G�l<.��8��D��&������ய��k�	�@�ҥ���; �h���P���NG����;�L���9Ԑ��!�k1P��>��АTy��)�w~���#�h��$Yx���ͯ�q��]9OV2��9Y���(�(�i��Bpm��n����%�o�xm/�C�2?uN��bg�y��L��7HD�X�s���6O�.��=]��f��Qn#�<?F�@��+W�PlNMe�'���.L>���<�{p���^2����Y�����Z���:K{D<<�Q"�x�+{��4�y[ I�����M|̪�/��F͗9,%���'�57��K��40��<��ˑg��M1�R=�30v�u��&������[e}w,�ˀ�rV��4��6#Ja��U�e�k�i� pj'���aRq�J�M#Ԉ���L��Y+W�=�����9�H����o�3�t��	�{���h�U
����e�,��M��V��_7~�!N{�F����b��~+v4�K^��_0��ݜ��i����y���Û���[�K8v���;ztz��I8�����Ӧ�pJ��ݽw�Du�ףr"1���L��I�%%'�`M/��S�6���F*�+}�x��+��1�,KF�N9� 2�~�:ic�=�*�;�����~(�N
����������ju�+3���O�sSGK�b�ר��[���?z�zc-���	�fɀ_���ֺ#���n�z}�3��d󄘘���'���+F�b2:F�J�g���.��E�T���q��A����X��@
4ݭX�(�e�)Ȱ���y2YX�b��]���F~`9���%YX�D���M�'w������b�������vex���=	7�Hu�!{r�����kR�yQF~G��Ӡ�=��4DaT��q�^����#���_@��c��b�!zˈ��]�P�%b�C��f+�&�u�4�k�k��igi��.c�yIkl�����C��ض���R�Y�d6����EgȳW����2�,&���k^��?	֬A�}�0`Xe���,5�VIPgh��=}]����ź}N1x�D%���P�u1�r��/^�<ǺJ�,5黾��lp�%(c����!b�7*1w7�R��W	u�c���d޿+.������� W!�a��Ń�c���ۘ)4A_?%��ap2?+����}���eqAg8�A�l<A�gH�9�w3�;�`�*}�R9'���|���T��������� F�P�I�����5s�-[����8iX@ó���ܗ-ʉ:p0c}���z�`:r���D�wW<�$*�,��I��2:(�fR�����U��SY��ī���}�a�r���~n��}_??l�D�Q������akml��m���U�4������ۇN:E
|��W��*ҿ��Ժ��șuYb5�@^B���RC��N��|q�
���"E��~Js�]Tc܌]9�Z��)�J�C�"+5�g�z�*K�����>�/��b��g�e;Y�ڟ|%@q��A�NI�q���E]C�����t1H\
���E�� 2c�T����6�d�d�� ���߁g;�>�d)s�5$���>��o#�/��7e�*��i��
��S�U��W'���Z�8���C���`�_R�d���+׏��������E�Lc����'�	�����E5���/�'P珇�Z 5=�1���>��Rf�fvk��S	#�q���,2�
��*Ui]�FP,�EXK�TuU�ѽz) �����v֊���o����[6K5��Ջ�D�%@x��nTZ�}������w���`��A\���j1�2|�iܽ)Ӓ��刄��g(�����b\Nu�w��<S_�l\"�X4:�����:&Ҧ��8���5[��%�7�"��%����=�p�`��(�R�[wT6x4���u5�YMc#�&�Bi���i���\-�K�\d�d?[�����;��U�F*�%��n��`�KJ�ےCw���P�~c����PS�&�D�����z�ݜQ�u4��Ы�|��.v�GFEmc�ʴ98����E:�oj���X��C�d��ɬm}��5���l�S_��ܶ�^�M;�%����+c���M���r�Ȉ���}Z	�Z�2TN `zgp�$q�:��8#��5F�+�N�.�'�%6�1��re�U`�W:PV��c/��Z�Z�Nr;��WH~[�Gegl�.q�dC�е>�vk��:V���q0�$5Ol	n"kg�B@�"�?�u�D�6��4s	�47�a�����3�$�Gq!�S4�.	�A?����>V�D��'�&2L^;4�X�s�D��h����=������~�1ٚ!
ڙ�:�%_���#�<�|��N���X=��R�ؐR<�z�j�~ӻJ(�
p�M:r��^KI�(� 0^Up�~Ӌ),�"c #�����nE*:ȷ�I:f��5/v�u�w��0^ɼ�h�=u�K1"�\$qOats�+���&����[S�%Y��uG�M�q�I����(A���ϐe������&�_W'�^���0z�uT�!lC �fΉ�,�If��g��/���ݨ�Т����^^�K����Á��qP*���$3 Z� ��'Q�5����e�q��	��[DsU7�/��X[��ي��i�*�-$͙iS���y��PE*�4�x��x�i����5�}����
s�hb�3�����P(�P������If�xg���E��4H���\�*�L��%]��T,��>�W�~9�L!��^#��Z� ϕw�G�EZ������g|F���1M�3�`A�x��ْj�>G�񏅒���rm�R|g�)�%}�c�(�̦��C�I�\�7O±��2���7"@Kc�e�c�}]N��B͖ju�R��!1��MA�2�o>9re)�uՉ��OG�wNp����һ���x��4탊���VVx�+2-���OB?=�����q��|�;�T��x}����Jae�Z�Rk�7��h-�t��m��=@�G��z˻�l����Z���z�-o�71�Q� *QҮ�'�65콟�b:�����A� O��,�*� �;S}>}ӵ����FMu���R۲3��Z*Z�2³����l'�YQ� �N@�O�۞4G|��%�1�3m?��bxW���G*XQ���h+��	��80��l./�M����dl��~����6��\{���Jӕ�u�`J�w}��̶7�q�o��� �h��p���+�~�����G׆���
��ּ�Q��1*R���-@��`�vF�>y7(�>���L�VFQ�`�=;B�6�唛����k_�Q�89�f�GS���{_A�3}l&
���E+I�+�P�q�9Qg�%�+�d�c]t40��؃<	}�[�
��	�j�����ήD�Ggxjp�����l0_�����'k�_���ۛs~g���c��'�>pv��Ǿ(�n>�����B0��/Y�ξ
��xw�7oG���X@-2��Gt�I̗���H<�42��� �  ��Ƿ@��{��	=������
��Ř�z��[�.�Z�V&jb�ic����`[T�<�
v����?�*�i�8�l�=�(KzÂ�T9�h�u��ۯ_"-�#�͌�&	����}�sF>0j����L���}�����o��7�A��ǩ9nPY�]���x�Y�U^���ǆ�X5���\�:��] �0���n�^I��/��
���e���YB�h�Jw�M ����TOT7+�;O�Gn̾q���KP��o�0e��J쌂�S���B�MҺJ�EլĹ�����\I��۸陚j}n_��v\�4a���;.>#D�/J�81�֧S$�Ϟ�J��9b6r�� �bKTqѫ��k!�K��e�������1b7@`�eWn	Lݴ��q�b|��sd>���I�6ŴoX�{�q`�*����nP��olSD���OLM~���4�w��jj�;��rE'T�?��ς}�ا��η���a#��u�����>oq�e�iӠ{�PQ�\B6���\O���3}����QV���OJ�d�/�DjP
�oC>����U���������8+H�*+���qנ��4�'HW��ҭ��B����rp��"���G�9;�X�3\qh�~�i<j:�"<Ѳm�,ř���6�0��B�y�$�����]�I�{�t}�e׮�DtI����p�E��haڪ��M��ΑF��}At?{u��	n�!�p^���P��&�꾋���_���`��Wq?���lG3����mZqCl.t���f\��!�j���Ό���F
�kJ ��~�=K�,V߹pk1����3�cn0ӯ�K�~"ހ�.\�6����Uv�����S���=�I���s�:��M0B��-�n$��,��VI���G�?	`^D7U5����Y���K�v��B��L�E���B���!%�~͌C���x����1jc�N���J�iW����QC��|"��a9�B�I_Y񎊭�xG6���ٜd���bw	�ch����Pdcծ
��ir���n��dA8F�~�E��#린�~��q:t�bݝ�O)N�up�u=l>gjh����m�{�cG;ɰ�  ��v�8�Ds�
��.cn�@)= ���,F�(����:�IZ�v\�e6��<�Ɲ%���Eڊ����u�f�|UFm��Z:b��n���� �4�������KK�
��!�]^��|K���6͸a�1�&��Ҟ=kdqF��U'hMM
8
|rX��H ������?�{W Q{.�s�.�Ќ���E�J��lt��VD�x�RO�V@t��S��j��d5�ZaI+P��v�P�l�[��$�%06�g��^u���ݔQ�՜}dE�f�ǽ���O��m q���3oҔ	^]�Z�),��f�.�rğ��C>�BC����b��JQ�ωb�I����K�|�}v���>�O�nf�E���	��@�Z����D�KD�q|I�X'Y������^#d��$v�Cq���-�@�MA)�� �G I��URr'�#RA�a�����9��x����5�/W�~.�O6��bU�l�p;��v��K�c�?�-P�HA�^[u����J�V��<8��7����Z$���fv�,��I���yq���n�IԄ�u�]�R�D(n�*@�E�}fcJOi��W�E�#��������C+�9��[ȼ@9�ͣ#���ِ)8�sn���ca(����Dӏ�BJ���J"��C���Bz�L���;���lUS�-s��rxPDd�~���]���Qk��ƖHg�gO�D�ؒmx�E���6�k6u������d��yr9�/��j5}t2pѠ�qΩ0� ��M�����t������կ-!�C"k�g$��A�c�z������4����B�^�����͹�q��9^�Ae�Q�z����X3�9M��N�O�b�\���K]���a��V_�">3�.eF8�����X��z�U���B<s�´S��m��<�4��㣊�&��L�/硲��-4A� u �����YN�F�:���x9��BC�?4�0�^<
���J�M�S^=b���ǳ�h�Ui�	ݞϳ��˝v�#r��ed�Y13�.9CeP�'�f��B�4W�����*D#Vǝe)���ܱ��^)XO�Oy���`g,�1(�����P5���v����o���6\�.~�:p�ji��-��&[�$���iz����7�G�<���Ā�����=Wc������N����:���n|�o!�7��폚�������z�}��N �6�:8':s��# �+Jj)H�|:��~�N�z���-�^+u�����/��^m��8j�!�_{��b�Y�^�ǉ�O��s.�Tu��ޭc��H�*Yɟ�aHlS��<�}��,	t޷Bަsuݒ*N:k�?����K-�¹߫���7?\�L�|*�����F�(� d=|\�`"d����I�/]��y��O��?�>��@�7�y�r�qS�������?l�R�_'u��n:���������rة�,odW;�Ú�A�bg/ �9j�!��5���w��VRTo��I��7]5���]�M�}�u/�����^?��w"\lЮ(-���ԹI�� 2,C�e��KlT|���F?G(�@pA�l�dNIU�H��\��n��G�)Ν��e�w/8��:�Jf�kٗ���^\E������ڙ�H�u6)@Q�ߪkB�: ���������@���J+���>ڰS�/<O�}w��c#Jn��n-Z7M`�q���Xa�Uǂ�M�||~�z_�EK�b���~wg�/֐� ��eﳉ� z�Z� U�%��8�q�34��LK��]���J.SXA�Y	r�e�t(��*��㞝��U�����E�4��A�VǸzl�#�M��!�������Q����r��-��SAl�Lp={��>�</�=Q:T�s�0���&�/?!���!T��5.}t�����ڙzT�v��s�
���v��i�m�/l�����
��l��oᭈ&�Ni优{���Qִ��9�3����vV6X�R��oy�6�h�kƍ�� 5%w���na�7#���w�����u��k9�|U������Kì�,�sg�ߡ��$0q�>�v�%� Ú�ӓM��>B�[��w��	d�@P��~4�z&
��Lu`q�$�X�fʏ�e��[�C�I��+ϔ��UR�}$�	�@(#�A��U�^6:.YIy��Ÿ�XΉnŽ�u�\L����ۓ�����R|$\`��d5�5$=�C�Ƅ(�w�E�Աޖxo^~)�lXP�u&�3N��s,���P�M&CHj�4&�/��+0�v�L:�3\�5���m+�t���Z&�W]a����Tmb�c!���-�p�c8�m�ovg���B��,�6�)���3��	C�t� w̿�F�&Lo��1�g�,l~��Ez����� *�D��X���,��ڕ��?��v9��^���Qڝ9�$���%y~��V��v���]6��Q/�A�w1vw-[F�"y�Q�� ~R�,�7�����F�ąх�bq~')J>�$���O}z�Aa�N^��)��S����&���/��]��2Q�)��Zb���s-B缽������ܾ6���3�#1�s'�J7?��*5��d�c��/;����>u�_�^F�;�.̰���5�?H�J�'���`�צ ��T-M�r5����ra~R�Ѐ�m㔯_�Υ��Ge���:�Ԙj�߾�r����9H��y�6��cwD`Y�늁�*�9�ri/�3���$n��!���t慠Ңw/���,���K�
���T/�:?��y�+�d(n;����w��C=Z|�k��"��:�� �G��\�򼀶�BΉ&:��_ܢ��]e�~��VL3
E	�2���R��
�"_��Ű��M1$w��/^�9	������1��x'���}}o0�#s�zĄ�)Ϛ�.�VI#q'���̘7���~y1M�OF�
�O��V�RVA��k1��J��%	��)L
�TEݽ�E ����S�N�3�NZ��ȱ)��%]������>>������9 �x�6���٧ЃE.K	i��e7���&���m*���] �� �y�Q�j&�K��y--r�S�S�/�p�����E%kD���c��:_�p�Al40Y_�'3��O�8D��O^2����ف�( L�E�q_�:UXP��u�ѵt�:�����"�K����(���4�Q�v[1v�z,�N{��m�L5��1��E��� ��D�'���K�0��L��_�0S<rK,���<B	�%)�����lG��ݩ敲j�<!%l	h��N����§��W�vsKjݓ����WN֌cC�[������0S'Z�;�T�~`V^���F�I�����,U1��W��Ɉ1ß���5�M�<���o'���<(2AaY�x����?;�WD#���ܲ\�r��X���Ʋ����!
���M}�x�!͟�^J<��#�����K�X~������wc��EA��{�)�R��Q�"2��H���T���?�
���;�{��R�*�gr�4�ma�;h��2,�F��Ϳ®-���trK��5��$���&�G���e��a0�U��d��ܻ���-hgy�#��e��離i����4�*�������k-`��-X4r��M� O}i��YP��{��]���G�AN��_��\i��8�(+$[:��(��u�7 �b��"���<:����t���'b�g�b��+S��*�![��A"���ğfN<��d�㞬��&My5؍�}�1#�;�a8��c
���^b=�6#.]cT��6̈́	�޵λ�$�\:6��_����k!���
&���
�^q�^�a�	)󖖻c~u�\��i��K�J��ê���Y_bE�2���O�^�,�;�T�r�P	�m�����lF������2�aP��ό�t��Cd�9�:8!@G�j���s��
�g^~�5IGq��	Ӄ	���$�t[9{�m	;zYeI��ppփuWc���d?E�-�����d#��!�Ll�+[��<0.;%0���: �>zs�l��I�n�c��qfMf�c��:�,�B&�����nQ�?C�?��S법	��@��2�7��>K�x��û���m��1��S]��*��X87AKyvd�ҩ�z­[}�G,�_LA� oX+?]�ga��9G\S��V5��>0�φ"3�٭G�u���<����4 �ϕ��ɪ��p�i���N����7�c��b�r��gө�j%�P,��l���?'�W~Sml��p��Ġ���A�oZVԊ%����|�d��?J�6b���Fw<O��/_�=���f������0�kv��I🗇*����׈�O/�3�PlDyz�.��XK���s���܁S��lS��b�<�_��ϭ�?��2e?�A0�hM[.84�D6�k��h����Y��)���s�G��'�ab-p�Lo��7H0D��-f"́�����{�۪�K��ɗ��+�g{~M�/di�c;�}>lA�<�	�����B���{�A�>�Nm�9�����О`A!�;&N�	��0l_���h8X�腕&T7�4��b�1%B�A�����xR�6XO|��l�N����.c�ؔ�hG��X[�+4����^����c��-��Wkx��0��3Pf���uU��ĵ���hSOXz�V2=&�s5�;��O��A���W�]�G(m(��I��Y�B����-���L����� �W���a��'r:�B�E!gNL.a�B��6�ʆw����Ъ���W�_��<���\gJ����z�;l��zO���Ԍĳv��ɹg��]�2ɢ&�*[�fH���h���YYgr��5��Q��[/��i^#u��Q������=4a�r`���k�>�����ʩWi5��Owb_N���~H;�����N�T4XYS��X��s��;e�)ͦO��>n�$���4Ћ�,�D��&�m���\���g��B]��ƺ��ՠM��u������p���8<6�����+����\vb~�>��������Ø��<n��,N`蜲���x�m�	��c���L�͵H�����T�F{;�
����r��HZN˼z�_wH�bg4)Xd͗�7���%�g(>+R�*�9�\t�j���E<4��}�'��u����پۣQ0����R����&�{�6��?)�D�ː�2��B��@�N^5�9;��767r�@Q��+7g���N����\�gܷ��]�������eYU
k�f���� ���*Bm��|���`1��ͱ�����������;�c�8�6H�Fp���M�:#��B�
#���oH1�N&ެ����Y��J-�%��M�'����@zT���C���ve.f�:kEg`�hF�^p6��	NC�O��ػ�.�hM��s8ťt4�,�cp�p�B	@Y9�%�P�[��c�����-&���Q�&kU=a�X�)SY� ����6C.�@W�yܝo~�ZM���4����l	{�����ڄ7 �Xf�)��-Hs�
��ט��t�B���d���r��T�ǂ�E��8j����b?�5�����(�M�e^�
�	U9�QBx;����9�bk&��- �o��[�{���H��|�x���$�w�esH�x�o�EO��S+��S�r���~�ea1� �:�H��j��԰�W
w����ԫ���59wgo��IK������
�5�b(�"-30�/%%��x3��&V�ݼ"�����/aŮ�QN��"�t����
��C�l^s-ך�~�ԅ$����捚���%I����?��?7����A#����ƍ�@U��1���S/ɥ�E���N�0���&���� �)[5�a���߃� ��3��~T񕘒IL�9��E��eH��<}�g'�X�k�, no���/��5y�):��<9���٤E�oպ�ߤ&�LۡNÙ�b��h�����s-��Z�,xOLg����ȋ�*4l,T<NR\pCL]0.�R6�,�.�~L��֮���Rb�詡&���n�ף�ج���N���^�J/�6��t��g��"�_�ΖUX�Pr��Ґ�-��&W!)t�*7����hE��<�XƁ~��1��Jء=L�tD��rXw���>ࡦ�����"��5b}Y}�J�8K��c@-��M�Ou�M�E�|<�����;G�^� I�n���Ȁ# �!u��{g�q�&�&8Ow�#�ŝ�m�p1�j&�C���@h��CZ���L���^n���[^Y�ajA��"�I��������ZJ���}rF��rU�����t����?��{�;�Z�}@�Њ�]�a�  |��o�S�Ɖ$~N�s��3�]0gT��:g:v;m7�0�(����s�t�c(�@��O'���}���f�O�*���9��Z�&�@�<n��BV�8����A�bFxY�w=5 ���яgxl!�#9���xr�P�mq��ux{C@,DE���0�Z�	�We	2���e�򒬤��i�EqA�>�y^O�~]�/��ϐc��z�?�pЯ'��N�����D�����5�k���;t�� mk��Q÷d3�<�&�J��1��9��C� �h��08���?�#��H�X���ម�H��V�kn)k ᥿�f<�n�-4������ǘ�������-';˰��6��@�ъe�$���n��@�dF�����
ǿ.s��A���/;����m���=y�ِ����xt/��#�����xa2�����G?��zZ�cia9��싶%��k�
��e��@� ��TB0��j��]��c��2i_�6i�f��L����U�h�T�:�x�H=�E{|�֎�~r��=@�N���2��	�Lo"�r�_�:�J�]~���KՃ��B�����rK�����%?���$�$��uZ*��'���=���<���"t^XAs��'�Ϩ��g��J��
��M篘\%Xs��RI#�8�#1���a�i�F����Z9��326���\�j
�d��b�)x@Xe�%UA�o�����wG1JS��@�f�{���	_ �TAu� �bѫ���;��2��|7��#��'��N=��uɠɬ���}.@��=`����qp��b@.O���S�㉙�m�賷�J���|�)���@��:���JO=�"ЋFD�ןXa$a�ws�I����#��{�\$���'�8�r��T)��]�����y� x��)d��c�(�b3	�1l[�����w�����?���6��CEPe��r1���;�Oh*? m�d�HS�9���v���#�֊����L�O%�8�� WC`+}�wPFK��
�.Z��Z�2����樞���øb�^�u��CC!.`^B0�z�� Pv���併���mHY���MFR�"?��$�r`0E�w�}gd�4�^�%)�EI�����@�B"�Mܩ ��~=�r\/��U(�q����_W�'�X����\|��|o�<T�Ks��D"8�L\Ɩ��wN��J��H����L��߶]bQ�)���4rB��a�"����86��1�ZM����Y�k�AX���l{ȏ��"��\..õ;E����O��h�\@��n:�����f2���690�+�el���ag��(��/�)ͭ�%^���A,3?Y3�4�
�1��Z����!���e�����bE�3��#�Ɋ�/
݉�i��r���Vvߚ�x�6��8�)�Ь�K	{�Ү��w���
ߕ�/���1g��|�������u�q5JI/B`5�w��������~�������b.ʹ�A��&U��<�>-s��~n��Y%:g~%|2c�ęI�M�@f,�r�|$kڻ��b�k,ɶpr�C�;*�Z<�B����8�����(�����D�t*K9q8>{��ڡ�h{ߘ ��~��Ræ������|���"�.\���|�"��W	��6�$y8���������-��V�T�=3Bx���R��k�2e1d�?ޯ�A:l;
e��&e	uE�9�k4�:�1�x)l�,q�{>�u;��K���Hxy>X�VUxQ~s�[��(*A�0��D�a1G�c��7��.��z�Ŋ ;j��6��_N�䠸�+S��V���� @(��=��"n�v�1F��4�V��2m�[�;��v�96�H���v�5�v�q��(2ml�~u�~�ë�*�W��2��~L��.ct��V߃ .�"I'eEL��DR@���~�`��Hۮ��G}� Rb_Q�o�z�m�H�f�r)�J�O �_^q~m`l˱���g"���;r��6��_�w��� �`9m�mꕮ�^�Ogd5 ������R:�,���./!��dNݏ9j��G2>XWL��6ɰ�UC��?gk���z��":�uL��̿+�3C��®�sh�T r.S(�朷��w�a�g��/��F�]�SlȦ�گM����O�_g�W�:��&����?��c�+�H ɼ���Гy�\??�ޛ����q�-��g�;�l�o��o�c��o���=��M]8�K�PT�a@�J��|�q�3g����nmլ�M��h�eܖ�.���+,�PĞ�~��Y��oIuT��yu�n�e��`�/��q�r�6K<��)������:��3������uUBKL�5H�7$��>f(&g�D=�Z�&{�Y�oâ�l�l-rht�+�[����-C��GdW�H�{ ��oo��_EsgT��c�9f�(�k�����_�L�h}��N^�`�s"�d)��@�����+g?wG'�m��B�L�[�����D!Љ�%��\��'���eu�R)ś:���B%&�@��	�D��[����7ҿ��,C���`p����%�$`$�� 4Q��]*T����4!7����2�^��%?e}&��6Q!��������L�LG�p�/U��r�{W����ן(z�����k0HR ��ۀ���� ӟ��,�=A��^��
��.r���S��]Q��`kþ�!��|d�Wȷ�gl}�h�����9v}�$0׹��rT�yMxsQ�f�Q&.*�ks�-���Sx�α�Ġz<���+A�����׳��%����p"�2Kȥa�~~�����Tb�ڎ#E��"����G8����*A��i�0J�w_C9�۹qo�	�r�QB�cZ��#���l�	��$�R��f�^�Bө��2&yB���a35~���ۏ�[��;��`���̈́+{a�i��/��b�`?S:��i�G9v������h"�_6��/�^�j�ټ��3͞H����ޜ,��!�.���$�P���wFo�����-?���� �}�L���e�x�g@�}Se�@,r�~���{8Z��Q��Ov�S6�Q�熫>#����ֱ�}[X6������i�ɮ�_��69�8>5�������=-F����/l�t ���>^� _UrQhZ��rճc3��Z��/X�T�+�Y���2}XR��^6O��3.;�`lu�����mʒ��l�±y[�,���8$K!	�[��8c��U���'�̶���]/�4�u�'�N8S�h��e���C$�₤�#�9M*��TEbV�7���&��C1A��6�nv��ɻ���@x�a�{/�b�sd���t2��޺�|�s�:s��a�A]��W]��T�Ũ4 �c�5�w���4:���	m�F��b��HM�NQ�TvPcM�O�>�3�p{���*2^�C�v+@�4%���k9��������&\U�fù=����D&���� �U�L�Mz��8%����vG�����2��	~"�b���xUJ�np�����z~�������u�]��-.�$�g�^�O�,߸M}
��2���K�Ύ�ma �O�����"�Y��>~�?:��-�,�M��kW~�������aL!��	iD�;W�J�7�#�@w\
V
��Va��q�3�P� ����4�e�"$CjQ*9��y9\v|o�O�ָXSE�W�|���6gf�i6,�����+��� ����Wƻɽ���e��N�65�R%X�?�=��lB�Fa^�=�~C�Y7���&?i{� �eƂJ
���n��V�^��u�7/h%���gGYCo��?e1O��V�u��U4��t�K?�/-�xX�=�N�d�{����+,"��K9��|��:
�h���q8Ԅ�y��dC��T��6������ϻ|�b d�8eW�w�݄Ĩ��`���!t����jfTT��6A��9�}o^A=o�k:�{p:�2�,��%|M�1N����V� f�]�z��g���6eT�FŅh qm��+��1k�§KSpVy�H�d��� ��{m�iާc���!����w��F��t��4��_~8�=���~�T���_/�|>��*�x��>��������A*.-3P}C����u|j:ۆ��Ҏ+�w������������ųr=ﴮ�?�_��`Wi��o���Rܣ�Q�dJ�Tv�'�9��*xb����=����Ӿ���L���L�g:����!�����p��RV��2��bw������Z�@��܊�^�u����R�*�\�h�8�p�9RgL>#�D%�F5 Z:��$�y��[&�K��Ka� ��R���x�w�:}_����IV|$���<ߍ��=#�L/�Oa6l����h��G2M _�%����kr<���d�P9n���SW�s�^�3RSI��y�����V��9�a�}�`�EQ���_�������V��{h�����A�#d��=�^�V՟K�ا�E����J����R�3|,,�sg�8�=����_����6 ;�~&��t�ki�G:�C�/Q�xJ��5 >8K�ܘݻ���΃�li��y��mX�X�!��=�G��6��8��uؕ@��U���]�&��ܺvƎ��-ɝ�ǿ��[�C��(�faV��r�/��e����"����F&�
0<+K��lJyfl���k�m#�샩�k\��\�E��n�����U�P7U��Ec�>�G}�7���M]	0�R'u�ɻ��uݞg�l���f�k�q���p�����?�-�v���ƭp9ߋ��o�ȕ�=`z�Λ���jUΒ� ,\n�!�{�
�Mq�}�U�����%W�h��".�v/���+o������m�D/�6r<s���
V�Z�-V��鍍]���=�=��q}A��خfJ랷�����? � !��C�I	A0�r�.-A6��Wo�?�D�i4�p\�X*V�������m��n)��I�݊�:F��s��|��`�!��`�_!Q�XC	5�`���GLw�~��>�}=���u���A3�z(�-%�MF��+S8��j� $�K�	!O��(F6v�w��"���120�,�M)0?D�O��)]4%UX�r��G��.�I�ȝ�`;w%cH��s
�>����fq��x������SRYˬ1�S��1���x@ʘ���TH����z�e"��|�R5��ȣҶlMA2����s����v�v+υBr,�6
%�����x�o*F��LTD�^��t�+�t����@��5�#1q�I����K�uhù�Ύ������Ck\��G9�(��H��*4�dV�z��7$?c�J��&���n</�]}1���L�T����|v2�+#���Z�J��&����I؆��=�-�Es����Hsna�VU�A�H˛���P�X�^?�u���eSc>r2����R�^GK�g�����L��	��	L�_S�������C�{5u�(��-1k�!������T{_|.�QG�3�[�D{�9�����je`?�u��!�;��$��UCFG�z��Yy�#n�8m��p�L'qZ�d9����ݠ����9t��]�Y�$~�I�p�M�͖sRn���-�%埝����c��v���f��@���J��w�u����G��T�F��i��}A���0-X��L��i/-�J����S�1�����h���h����{*&��\��4A�B�
��=�N˱�h,����>Bk
n���������q ���+!AS�Z^��_��MHh:�&��uʆ���-ח̢;~��'���+��M�e���o�S�R?o�`����;J�(�Z[��:lo�/x?��^�pz�1V�1 ��>r����槕$�?��r�;�;�����-w�:!�Wn.9���D�Qp��
e˩�x�C��`"�RjBz��DKf43��5���޼���٥�|~q�����+K�X����N�VT��Ѫ�zW��ō�X=�����'	�]K�i�G��TT)_Is�cƆ�7"Lj�U\��	�����{��ڦ�N�Z �/j�d ��g!�Xb�mzml ���/s_�;��)�!�k(�����r����L�����+u�x�t{�g�*_y怽O��
u���"+�Z�	O�����b0��O��ƺK成��\eb:KO�����
-#�L>wh���{����=�T�Y~�AH�����������m�D ���Ν��(�TB�Xy������k�؊#G<R����f�"r�0�� }�_ӫ��n%�)�A��E����)~�" +��KR�~sI��j�/0u�������"[�J�A�7���e�a9�����l�$�Pz� �*0<��#��� �����/�N,(H����sy�2�E�ݴ�yB���{��ˢ\fo!ៀ+����b:i�����L9p��h�7X��j�_��V&ys]E�3~��� %ͩŌ���P4�D� ��vjf�4�œ)���&�.���f���B� ���=�0Y�8_3_Ԅ)��2q�2Q��Z^���|P���2Q�h.qD�kM�R=g9�XzwA}���O�6g�n��,:�'����3f�p�����Kʧ�Vc鶇zsHdiZ�6��+:}P�<r�`[e���������~] {��[$�0��p�'�r
���(��O暋�$����w �2�U "�!@^�2��]�	(=�gYY���C�_�"S�����q�	���HP��u�H2Ն�������=g7�~�s�XA{�[��W5�3}��f�-�jtQ)���[OpZʫb�I\�� ��(�B?�("�<�����сY�/AR���ƴ�����s���|��œ� ����=
J���߄H+�5e*j`!?Ey��a�|����#�ܟ�{�82�[��qt�Uqa��*�=�,-%���T)&��橢�c��D�9���2����d441�.��888.;#����
���v�t��r����!h�a���y����5���5�w�A]�8/��w6_�f��\5j����_�+�	��x���s^K ?�SAN�j� ���nɸ�F�I{Q�t������R~ռR���t� }`{�4�.9:A��0�^V�԰esE3����v4�qD�͖>*���mS�2�e��J=���b���WeS�X���	���*��\�Ȍ����)�p���@�~��_�"�y7JB��}�/���D\�8�u��� _��0���SU=F�?��Ӧn򧸓���������V����S�>)�C��$�ȯL���s]�@WژIUj��*�x:����GqE均��z��`�ť�ͥ(�q�P�����,��1Ahő�l��[$��4.uk�9kT�/;ި;�3%����c���!�C�{'�R��Qa��>}_&h�ޯYiD�5Vr��J)��A���O��N�E*�Si7�*��r�$#�)Z�_�>�@��-p�r	�	���E�b/��^_a5�{Y�R��L�5���_�f�Mz��M���!�Wo�j���^[�6js�m࿴W�H�h���(m�9���m4c����� F<N�bm �s�ϥC������q���w̟$�~N�	�������فXO¾���>t��7Z���� (�6��t��������$����Mf�~�P�͠|��E>�?$t��+�c����:�&������-C���ܿ��k��gzi�9�c =(�%�����E&�9޾��j��C-���t����*�.����l�y�!�;�$:ߦmВ�}t*�P��J��Q���-
=��]�>Q������^���T;;4"V6�@F�4�-�\����l�&��WfK�':J�6���R]�n]r�䐊d~��[n�$!ѩ�c�Lj*0���ԝ�����&�w�D5L{n\�B%�^!�\�T���Z w�T���b��:w��;�jᒂ$�ޙ�HU���|;��l��AJb����~�h�F�ƃ�+�`i�CE�Dx&[iN)��M�cl&[bڄ�|,�dg�}ͥvAL��k�t�;Β�������q����4B��%��?﷑�����\�p�f�E��%�"`B���b�J��T�Ez/n^���)3,��k���3��&�����~�ab��6���#����]�?�_����D�=��rX�ط���.B�|�hz
���(˙aHS�5}ZE�[��?}�cx]V��n�o��i/m�AS�7����'ԏ��[��J񫴪%Eg�MgJ��3t6	i�{�OO�A(�j2����p8��V��I6u�y��eM9����WR^�C�����ě��RIF�Wt�#K��n���^��Cr���ZP��[W�f�T��� ;,b�oϳ:?�s⿞c�%�����%u��W��/T}�m�װ^��!�S����6l�À��)Sdmw��8��>x�p�g�����9B�f��Y��%��Q�"��Bi�Z�@0R*�8�>�jY��1�PZ�T�˼%;+j�BR�%v�i�/�^�Zv�&�>�;��ΰ)}�
�oM&}Ao�	E�F��;��Δ�H�Lxb���(;��������)�F�����c�XM;�M���P����!���qnh��Sc�x7ur��^S�bE֙5�<�#�A�f�������G,����\�T�s�Z۫�&�Z��	;���%_q;"��ӻ�*���S��ʛ�ח�eb݌|I�D�e�3c>��-xg)=�jƌ�c�0��%�i��i3@s �B%گ�	���j&��!O�A��&Z,)������|�l�j�(/�=Ԣ�x� ����gq�9;�up7�0M�K-�#{#�ȖB��aB�a���j��٭v+fl�S�b��WL��V�P�W�l�>�@}��w���E�%C�K�|�	]��������#�GT�F�~�)�6Nz%,���|R����`?�|�_ܐ�5v��ڄ%A�7ߋ\��5�B���a����L�(8�Iz�!X/3,�V]��n99����<|2/,����}2Ҁ��W�)zV�ǚ�WM��1]��x��3v�h���2�PZ�{�z�{_�^Ӳ>Z�r��ծ�D�?\���:鮜�Y�MrF�U�Ƴ6�?�\�����ߜ���ڇH?_VX=��x��'�\-� �;���{�+�F8n�pd��� ���.r���{��󢛎��?[,Q[7@���wzim���z߰�>�*�C-�Bu�.Jo:\DP���\RJsb΋���>�ݰ:D������۶�QZm�з��p��M��
�b��We�5Ϣ�-�$o�M��_V�����j��ةo���{4���)�ѵv�ʮ�������L-59�?&��=~!��V��)+=i�?�?e�)����@����T!y���	�Q=�Zqq�I�].�E5�M$�Z�%d
t�hı���F	��t� �<��>Ch��~S36�u5���7��`�iHMeyY�F��@3������!A���=)_�g���i/9L��Ec���+)�=��V��ř�,��_�~�	�לL���=?�`�]�t�ۮ,�����~-;RP;:��ፃ-<�E�օ7U �d���;���4�!�2e�i+�&�T�.C<W��b��U���!�M_)|���E�Iڥ�M66���8� ���!��ME�s*H�D BJ6u��m�ն)*U6���o�0���uNQ������7�A�x��3� qL��M,RA:����qғ��unMݖ����6)_��%�'����p{k�ˢ��6J$�F=z|ϐs|��U?YS<�O�����
�,�� �(1F}��ٔ?�����Y��^�;f[!4s�Y���s>�n��9oM�T��8�+����Q���+���=�-�����a�i���Q��.]J��J��|f,�&�Ug����i~�Y&����I����(U��f&[]o$˩U�+�a��b�ΫD�U%��K��o^��R��BGk���`|���)YaM�*2g����M���K���d��Lu
3�%c��d����X��3�PJ"�c7hTy~�������+�I!F�7r��ݻ~������k5�\��b})�O��&���͛�>m�8R�}���#4��6o���\�|,�����m�Y70�����k<]�/J/}^(�e֕�^���Laf����Pz���X_τX;���|,�M��Z\���
cAܢ!b��!�����-�P�h�lڶTv1���`��Ӻ���X�o_��PΤH`�� %kj���粒��iPW{"��Ξ����%�j\�k�U���^!�!w/ 4�O�Z�	=|.���ZŊ26ש�J��!�ʑʧ�L�	&׼�#�"�))�.Qa I}�9�V��1�����8���k��u9@�	����_H�STW�>؃!�l�i����`��t�TD���k��0U�IC|f��fCA.G�W~��ۣv���e��d�?�,�GS���W��r"��&|���l
�ߞ���1��i�ј.�F1��*u�s�nN���̽�*8�c<�*ج/͛�G��)�U�S���}/w+ET\��w���yG���\�w_����3�n���	�/��Ȩ�W>�����~�n�H��J�%���-�=q}��v�'�������C�a���p[PL�a����f��3ErD]���Hv�vl|�:��(�u��Ļ���d"m�cZ<�X�a�dq�l�^�0����;VP����'�O�ٮD���Y�N��P8`Ā�;ܻ�w+� ��x�KY�A�u��^�+UQ��H̽���c[l����
6,x�� d�J7�; H���i�g���	zo�N�]��Bޑ���~�[�xh�8�[�#�h4��^�(iǁ��9�q�,ˑ!�
�t:p�o�*冿)b\$�cƙ�?-X��s[#���P�f���ˎ\��~���!:�{��Uk^d|�O]�a�vqsf�J�p+a���������5jHqY39���RV�`v�q�C����!T瑯��Y&D�C�Q�D��0�"�i��bC�F�7���Ѹ,^�����E7)�!N{zs�=�!�zc�j����b�MŃ���X���'��yH���}��S�x�Ü��C�?�Q�)�H:Yq���dJ��R��Z�T�:&v;���)�U����WT���!؎Cr����y��u*uf� Ȟ����cq���sSRT�ir�ق����(��8���s ��3��A�: o�r��4��+q��,�f/*���q<9K�S�R;��y�L߭'��|"��ŏ�P��XL&+Q��+h�[��b7�x��ǵ�u�7'�T��F@l۽����zEKc̼�Gxo���-����"Yh���
Ʌws%�n˸L^E
β�v�"s�7PEQh��$	h
�D�ߘ%<����ﻋ��Gv��J��~��X���{�-q��PcV��.�ȇWK���3r3��._ZQKf@���q�/	��vf_����h[���3;؁�5wE��Qy9�(��Q[�3��=l<�@�$�:�Q��F�/F�6�$A�v1���/�n�}L�YLK� rt(/�RJ��9�G x�����������u�X����U�ӋH�@x�nH�� ��ff�C�H�8���I����-ndŻDX,�A���]�b�}�$p�OxQ@ç{���G"C�F(Q&G����~J���;/��@�L�M�:���$�]�Wb��z�Ʒ�3Q���A��n\$��Q6��t�1����co铯H�r
�W곹�إ�\�~���z�:֧�W%�p!,��)�n����N�6��"��~z��#�}���Q���#��?�����>gvE.k���LF6���j58]�����c��T�H�&c?٣;�X�+�8U~�iw�}���uf~��
����Ӿ?:�?%�e��n�X��.;$�I�6zIol��C@ۉ{�\�%�@~Q�	�C��qoTo�[E�)���GCk�#{\XWue�؄�r�&{P� zk���P:+a�|�Č������N����YK �0;Z��v3H�B�
��G��W?S=e���-BF�
���2�"���	���4��r�W��d 3�Ĉ<���8���\Q�CS����r=G�h ��9�m�q������p����
�����=	G�+؇4n���\�)#ڶ���2�F���Xf^|
o�	J�%;Ae�l�����p��ߨ����b"xx��:���e��>�~���4�w;*'��@o�Z��{�B�9Q0�]s��"�\Ё:G������V���	fӣ��@�ĵ�Lh�<S��B�pK'Wv����<l���̟��j�3C��;J����8��Q���(���#��j�C�<}��|�i��`�������� Ҕ+e���.��]rb�!v��'��%�W�X��V2�fy	v~ߜ��}
�Hj{ڄ>*Kq���@�^�Lu�}5�@�j�>`v]�l�j^׀��ф*��i�.����W#�9��MpsH��#�È���~�2���#��C� �1$�$h׾�Գ�1�:JM����و�����B�7�l����8���	@�T��_�1���fq�Lit�H�27	����'�B�JK\ѳR�{�օ��,(s���u>�L���+��w����w �_)
 �>] �:�g�h��O�Q,!�hp՝����~j<(�z��q�1W�M��]����a�˂t�)C@�qᵔa�o:���:g���u.RU�f=5ଦÝ����)�����s��;��-\%��s*�=+��Ʈ��!B�%@��T(��:��U��&���t�&��g%1n:(�������xS�x.P<���IG�i�B��䍬�5�u��m�o�ieן����|���Lcթ��	��{e?(��*G#����D4#�<�4y�ݩ� X	��]�Un�򄖳�>q����d^��[���J���h�����2��ɵ�2���$���7��"��M���!o�i1v1K�����Z��"��\��cd�u�B��"���/����ݨ�l@�y� �u�S7��$�2�Ktj^��hZ�P�ϱۦ�iC;[၇u���)RR|�X��d�⺷�/���mUxB�<��U�)�t�F��u���Զ,=��p�ݢ�_&���9���D �6�"a���?���m�:̌����0�5�K��_���mH_֤�O���Oۗ�;���N\S_����!�̍qWC���E�� ���K}Q�9��qm�AΩZ6w��jlC m6�{E����}Hu��MB��u��	�?��G.r����,uy�C����� 	���'tb{�Qkl�A,#����*�R�}��D�;Bc7�! ��C�"�����Ĩ��h4��m�ts�t�iT�
�DI�f���IY._sz,t!�7��cp�t����v�1?T��?t���a��q��i�G ��~�ܕ�4����D����2�P �Z�M�c�����F���:����Y6�(���P�������%�g�Yi�i�b�k�j�\> >WX�c[9d2��&�E������逆�9�.k������v�l���oo9Y6�	C#���&�-{�t���iӜ����d#��>5HOyɳ�JH)9af\1B�e�O^g�\�v�#�>��S����hG��а>��=���HOK�}}0�� �����2��d�/��<����h+��V�5�`S�h�W�Y�8�\!��a�!>S��>���g�lV _�Q��m�JI�Ԫ��������.(�HdM}V'8��%�F:`��I�@�H%����^��T���0�s`Ʌ���0�/��m�O�(��/���z�Đ��i� ����y�@>ۜ�O�${�S�Ҏ��	�:25��YC�<ī�Z�_iH,\hY㣆2����]���)���+#}�Wj�ru��cPf}]{�NQyQ䰩cwԉS&�o��~���}bl5�U���b��<�6c�m
���M��8:�0KX��)��|W,j%�ٝBź���J�&-�\�ԁۚ\w\��\��Ic������\-�\
�Ģi���*�OLO�֓o��֨lmւs��8<����կN��_����9Q�e(�#�X:"Q%i���Yf�]�e��9��ޟRL��������'�jC��O"�@-Ԑ��(�Is� Ē�3{쏂���N�u�'�֛6�I8��;����;��*L"��-^	��W�@��P��"���z%�j�f�~�}��S�NN˵hMhc�f��*,��<�/�D �6���f��+%n}�_�6��é�~6�2oL+?5J�뉅4`G(���Ǩ/
�o�!12aS��l���UK�O)��u�����xPN�`h3,\VEa@�&"-&"�onZ�Y���0�4z�BȠ�[�)Iz+��\x�d�����%SԥM��1����[�z�av82 �rW��x����9� ƀ�/�yr
�|����@z_������O.&%7��c����?v>����jd��z��`ⲀR�{K(/0�j���Z�:��=�8�W��@�l2&�j��!w�Wzwn�z������#���c$�#�G��[a[�F�t�����v�y|G�.�ʔ��K��@렗;X�Lc��a��Q+�.��$HN�X�ܽ��2u�ȣ�3t��\Ϊ�;��Gw|Ԭ)Z�|�e"�rSN�>k�NO����q��D�|HT+�x��\,8��VPTZ�>�5�|���	X.�"q*�ϥp`��!�;̹�A���!~�����6�?� "��ug����`g�ԥ?�ߤ�d�
;�{*��wM0}ư?Ob�X�$�{�ٕ>�RU0��c'�}_՘1r3.~�)�Y����J�J/��I�Hǁ ���{#�
n�-v~S��hU�אq�TB�40�ʏ�{�l� �!K],W�"08�2`�R^*�K����?��t��Lg�Җ��%�ݑZ�<ci��MԙQ�	K4ǚ̚˺��$d%\&�`b���BH�<�ڱ�p?Vh]��L�$x�C��x�a�Jtv?���:J�n���SZ����������d��7�pV�d�c�;#F�L"�Dt�Na�
{�?!�1���2P��ᑁ��ӂ;JkB�
�+�v�ȩ����ꉓ���~+)��$�ҍ�t�ы	�-ɬ/�~EL�	�x����X���Hn�-W{z���k����O���_�h�k�Y�o�a9n�������nN���,BG�}#V�I�<:���"�<��MT�7����oF��q{r����y�IZ�B�b=����J:}���A�(	��(F٪U�S�-NS�ЧU�0P.����w'�n�>F�CTa����vPm�߼��,2ܡ��Y����њ��f,�~!J�3Ol���F(���,W�ئb���|}��Nɪ�\y�����*��1�C<��347J��*,�{G`�d�ƓWˣlUQ���}K�hF[�G�UZ�em��!�8�fHEz8��;O�����b@�U���'�~�ǭ������d�+�ga廎���䬆�)�J�x��GM֐w�R8`���3/9j����C��M�a�@Q��{v%�C�~�fS�'p�z�i�K�`ҏ�,M_�8me�U�9���;�z������Ua4�$b��$�b�U���+��(C r�:�fb��oQ~�������f�X��u�Y޳��-�峅bB���Qa{TX��MxE��U)��{��ɦ'o��2��$Z�����r..����+���`s�n�Õm��O �e���gz�@�4�ڔ��E��%��M �i{�2A��i#�����c�t�j���r��m���~���I�߀���r@�i��]���Mn���ہ����2�dVR�Kgej�4�ɡD.&W�������W{�k�oG!��D���%��,T�G���ۊ�T��x��4���u��L��e�h�va2h�Pߚ��!��Й�u�V��pV�,]��C\>'��) ��N���j�1�����%޼�Iat��,���`6o乇��)x~ir�xA�d��0#�,w�%�dX&b�ߪ�#�xc�+!�%���Q�c�&g{�u|���i�_^�]�ߠ������4�K{��uN�8��R�xa�Y�9��?DdLGs*�l��0�H����%���������P%A�*Ґn[�,���Pt�;��?gN<d�z2�Bu$�YЀ+�=�^Y��du�+�5$��3�ȝ�`�*���e.M��8r�?�4f���`
~��ČԘ/'��0�#�j�7��Τ��|�X~.�;Ԣ�d�nP��H �P����=����*�{�/lw@������i��{F�@q�fi��h{���_X*S�e�-�䏓�(Bϩ|m��j���6�����:)��m_~6)OSf�x&�a�7K���nJ^}��5U#D=}?�@�!�D�t�W�ud�Vl0\���:1��N!�U8/���9却&l��%��u�ChSR��u؞�TU"j)�Z�����u�×�~D�;b�D���݊���/S��"'g�zi��/K�ـ�G`.d���p�1>U�Q>��� �Q���7��C�E��M|��C(��$�aJ�Y�ю�=�*�uO4L��#ϒ�9��PJX�	1�co�o2Y�QI��K��vO~���Y}D��W(r;�ݨ//sbN��e�(�}��l%�[�%q'��䍋��Pa��轎t(;FIpz:���՞#c	Jkw�y�J$�ˁ)�@�u�G ��E��F���}�����̗q�r��0>^2�E�*{������@e��?b�Jl��~kh��	��6�
�Iy��S;�@�x��h�&9�9���P��}@ׯmܰ-�2��߅�c�!����mF���D�4��٩Zt�L4��} J�W�����-�|�I+��E�u��vfM���CEhΰ��*�E\ȳbS-�8Qt��ot���-#{5J�9� ���{��}�F"����V�G¶e�]����w�7N���;�ϓ�^Kը�p7�1�����,"7}SXa6)�W�A��}ᛋ<��L��'����ӤWFߪ���v�h��";G\�2�\R�N��cd5�F<X���Ol�Az�a;#p��Ev��X$�`�[��pXqt��r$�'c��ꁆ�
Fd���sc�y}�N�8|���c?au�}|��رؓP�wA����Ni�T�t�/x��=��y&�^r��7���|H�%�ot�y�<y���x6js�(fm��^P+dc�G���C��d�^�4�x���]�0��j�HSX��J��i��P�p�?'�:U5��a�2R�m7����]��8�|�E��f�H2{O�E-~x,D�'��� ��e\geZ
���L%�9"����~2;O�+b��޹'x����6IV�T���y͗޽�Yk���L���F�3�H�4����΄u�?6?.�W�((����B���k��=j��G=���ҙeB>́�jw�1Ӻn�=k���}\��*[yU���!��U �]�Q��%D*7��?맨�5VaD���/����U�H�k�hՌ6��WǑ��g+-^+y҈�%:AYi�:����R��;ư�ǌ�X�A����Z<��M�#�*���D|���Uik���&��{�э% 0
��z9˽ٿF�
ۂ���<��e J�n����^�Gmu�<o�Lg�	ߜ��]��;�]�?�>j{�q&�<(�G����
j<%�#Ia�Ȍ��E<�?=
�@���4��M��6+!��Tu42��O���F���G,���9۝3�8�"� A�$��{�a��*��~��?��Y6Ge,o�BS0E��ho��:\���blo�
�A����Cɟ`1�������5���ٶm-$\���߬B�r�qj���z}�i�ꮈ���l�X���m�ӤlS�6�i��[L�Lن��[�|����-�a˻7)V�Z�(|�P �W�8��;����ɔ0]�6���5~a-�uVd�a z���Nm�Z:͸��H>�^e��2�
�	:j���8��!�qa2� �E��.~@�uQD?���;����hF�-�~��EٙS����i_ph�	���i���s����W��ѣӴ�@��H��X��}�摽����� �)�}]����jW�nb�����Ѻ��Yh7�{����ڗ���EQ�7�sB�~H�f�א o�j�j�X�Y(�W�Ě�%M��a`��(��B��B:�ƚ�)�?���Ugs��Ƅ��^���V_������MJA��܄��H�[��g�V�� ����`��\����:
��mM����$
�O�:��Η�ѵ���XMI��k�{��IA��`ٻ�������i�m���ޝvڈ	��4�W���C�HU�B���&U��.�\��B	 �+z�>7�j�ԈBn��E�>3��@������ۢ .9l?'��I��zL>�"Miv��Åꁣ5�SO�L;$�0ru�����@�\edKC$�l'�G�FHJ�-��4����&=>lN��(&W�fόD��K3o��S��o1D�1�*�j������\"xC�<(�0h|�=���uW䪺g�$�k'I}X�.��� ��G�/��Ѯ�;�o%���f���0��"R_�Z`�h��i���u	��Lq2��%j�6��$��|x�R)��>�Q��A@�e�f�nf}|���l8�'1$�Ûik&nhx�C�+����J�u�FҒ�/�
�90p~�6��nq��Vi��L������Ĭoޮ���;����!y�p<��_�����r5:����ͅ`�ExFvK�q�w�`6�]��9sS��/��11LP��C[8���~*���&k�����:&�	����3� 2w0]�`KrS�ɤ�dU�^�l%�9��9|r( $�8"��>v�"T��t|��e�=��Zt�7��9������L)(��� �xc�v3����9*��q�Z�d�W���r6m\yQ��>v�*�/D�����������SM��2ջ� z7v�Л��z���*�t�ϗEfF� �;*���C2n��xô�LO���E�d�t��clOSf(��\��u�������EGj��H�$����z��[�%�X�6z	B���Y[;�K!�m�G�h����[e�,Z�h.��$t
��#��(g���s��C9���t�#�<$���H��kd;��=5�N��o���qA0��X��*���t���k�ݻ�΅|s���KS$rn�œ��8c@�7\~�J��>δ�x�_A��KtAO�^4�n����Y���s��Z�t�#�Q);EKzU��U|��:�`oS��a�����H�6"ָ���]�N��|��Q���
�;x�N�����Dq�h�j��i6��הr�|NDnq<R�c�D%�=�l'��&dx�ç���  [�sh��*�9nC�~�~��/�E�}�yA��9� ���R�����˥�u[����ըY4�q��n���Yו���E�8�|�n�N[����m݁�=���))��ߗ[f��԰���@�Y�<�[����^���;$���_K�E��:4��V��ե'����k5>A|	Og�� / D�;��~%���i�ٖ�/���qb&���ea��V�I+ch��Ӻ�<�]e���톈Sk�����r�h,g��r;������+�9��Q2�ь�����:U����\�|l�|P%��c��!�ı}��(�i��xc� �!�d[����|�����I�6A�M�E�Z5{w6 �K?y�\�㕙���
��1���d�dL��,��"��2���h�`:� Ic����zĭ~��Z�,�o�kO�X`�nw��'8�j#ɶ���ʚ���\�K�D7;�_(�Y 	�s�.JX
���wSbD�ʛ���#��1}T�C�H���HX��_ޛ+�1���}6�,N�|� E�G��K�> N
rU�$���8ϸ�Z"�H�3)X�u�w�+^��~�ޖ`l<���!T,�˙��m{�~0��$}i��:.%{����i��S��o�e�\���M�.�Q�3?F2�V�x�Ob��ۂ/�Ru��` �|����v(Y�Y�<+�9�����i}i�(�k3���Lο������� �fdeg-?w��c+<u��f�Ζ�|��kh*���3����&fhp'J%���=B����B�����Xbe0ߔ�YSg��P&WGffE�Q�³�v o���W�G	lvQ�{���,���CAd
�������D�^�O�n��lː�?��.5�t�zE��Գ��2;]_�Ө?�
mZ��q�F��ؕ%�*�
7<sE޿*��K����걳�,�m��m�<��(j��doz*L�(���o�҃
��w#���ɯ���(��r���p0�YB�,��< �Xjq��D��b�{��(3E�0�B%��@�a�"��*,{|�D~�u��Mzf�D!j A|RG���5�[�s3j8� �:A&u��T)�-V�^�sƌ����'	��G�F�a�j~�	㱨���rر��٩�:,{�XED|G�r�Ʉ>C�F��ukg�6���L������m���҄�م?��WdI� �7J#7��Q�	E@���W�l��ez�S8���%1=�ID��j����q���!�^���b�n���y�~j�E�&�I
��E���m�h0��9�t=h�+Z���n���Ykv�M�f�S�#��-Sɣg��,:�K}��Z� S�t�SXo}_���Oq�����&0���~T�U��Ҟw�t{���DR�E�,V�n��a�"Ԋ	hs#,��YK�P�ξr���pȕ����`Es���R�2�&��mÿ=JΟ�4R�bHj"���X��3�Nj����fz��eJ�˒s��"����n��0D9\��ܿ�ýn�Mʱ3�A�k2�j�<YGǱ/C��i6C��q\�-�G"$�Q!|3���-.',P��$b�XA��,�ml�l
6�()tգ�Kg�観6�v��@����������F�F�,7��>o�n��s�,b]=�y��̍�6f_} �W��ОB�w�i_�pL�Z�4?�nݎ�j~Ir���v
�)c�'�䁘�{�Ŀs���Ju��Sn�ڮ�O�t ��H4y��'ճ�c��b�%<W4S�!{�5�CbY�����Tϊ������ Ų���y��kF{񑝿F�ڤ"���V� ��W�����~m[��p��{�@�����_�Y��}��'�z�f
z�ځ�m�.����������y/L�`�$P����c���}�7`��YwX��!�?@���z,P;^Cj� ���Ļ��jxFL]�V[�ǽg7f��r+��U�Y�4�����C��?8�O�k�2�4#�o�rP�>�[�>t�Q�3c���
r\1���	c�^R0���Qwj:�8yUC�<l�y�G�>��N�
�#�vU��b[�Pڥ�a���x��`:x�;��a�H>�.(Q�]S%8�G�Q+B"�/���5����ʹ��?�}8�L�?I�����x�s*D�8.�u[I���헩=G F�R��x'e���H��	��B�����}����~�R14�h�K��CQ;˫V�x�>ٓ�p	 _3~A�����e�*Iv�p�dy�U��KK&r�o�4�dO%����S�k䟾p���u�@.�o��J��P���I8r���b.�ϟ�����TH�gg���	���-ܿ#�5�O��-��7&K5�Y16��T����7�+�A�^*���uM.��OP�5�+6��irA
�V�Z�X��t,od��d�pr��),�C�--P�'��Jv����K@Q@�^�Lu�0�R��,�p�t	��v=t]#�HOJ��rCW ռ6�zh0�l��Z�����\�kW�M�F����m�󫋵�Y+�yS&���P6�4��C�4g�9�ca�"�aP��JK�(�����W�ˍ$���hݿ�g��.�k�Ȕޚ\1�|��T�> ��Z�0�2�rԬ0�н�Lg!W����	_�+�2C��3�^
-�[�1dJ>���쓗\~�ͯ�bh[��}s9��Y4:�m�	��J��_��b�0�7��v;���I���-V�p��v��m�O�Qo�\EQJ$c���b�%R"2BH!���k�/�QA+�z�� w9�y#%ۍaS�����:SQ�*SJ�[ng��Ҟ͔P���]AmY��t����N'�2�i�M�a	�<��΍�Bz�O��UI���cG�QTv=P5n����ʚu'-�ʺ��	�������k��k�<q5j�>�����0R���*�Eنk����%�С;��&�5��K�F=ȑ���H���a�h������թ�%�[dד	�꣧!iYg��L�6���9	�@���Gx�͎SC3Sp�X�oLy�D>�Z�G���[�S�A�Y�K"
��2[�N<��C]����V�����Z[�Z$n�6cV���E+ߠ���A@�ʃ똰����W;P�J9�G�彻�`q�s@y�!W�(��T�IJ[�B���,ٯ�jj�t����e�~0��
Q�F�Vᷓ��;�	n"����L����M*��q#�����s%|S��)e3��_h_�>少r� �1����&]ٙĨ����A�q�1}"W������ܿ��n\=ܩ��Z��@+%غg'Vp���sRA4����%��∙"���|t;��c��<�7���侰w���v=���j����vz9��j�U�,M��e�&�X�hSO��l�'��T���w��q�d'JI"t��H���ڐ��t�,�i�t�a`Ym!�b�e��gs�i4d�H�F��n����Z҇�za�C[��K	(r�����%��(�5��x4��<��E��,>>��3��r2�!m @Z�=e�䠘y2��+����p�$�2n�l͛ʫ����R�xy�-��>�$@g�xfʖ�0YD���$|�w��x�#}a�x���-B4;	魯*��}���X$�:l	��Ų�+	X�^�]x�vL� �^�rã`��T8v��H;���;Da]���<jw�ij�b;�u�C�{e�X?�J<��H�H�������m��5פ��r����H��c��ۜ7T_��jc&`���f�j9�-�&v�@8좇_���(Ć���̠���p���7d϶M�<m^���@�6�w^|�1O�bA�+�q+�r1N�s��5�p�Ly�c����:<�J�}պH���6	�i:��j�$�x��@�3Qһ��
$as*��k��o���3�𞂐����[���}Mϳ|�nO��EP߉�?w���G�{��ծ���[۶�$1�<@��dPL����Td
��
'9>?����|���D��=�� �K��s.����*&���&'yC蝻�W=!^2�0F�
-)�|�4e���S��� jCC�v��3Y�8b��W�wW���-���6OnL� ��&��&7ث7/�}&I%���|��w_z��P Iɗ�!=w<�S`�����CƘ�ρ�(����+5�Tk~�9I��HҀ�m�]M�C!��hZ�����:/"gɴ�&
�'�ǟ��c#6��%5S���}Ӂ~S� ��U�#��0���5�~()ޑ�A�y��T�ʋ��%*���~�o��Tl\� 0�IC��ǡf���)f#5Hp�_�f���SJ]��4u��8��m�4-ݙ/�4�0��D�n�f���҅$0.�7!h�4�WH̗S���rh��U��Қģ�~Dk�P8�1NK����BaK�E��(X�,�p@�[�[�#�b�q���O���|�~Kű�5:��eD��	��4O��L�K� �L����d�3�K��Ĺ���4t�Cm��Gz���7�U�F	z���c}����-\)_�0��Y����|s8�΍C�� ~�6̶� �1� 9;ݮ�ht\�ƃL贬�7����z\3��(zPb����?�c��٩�������%���,�l��t��s�.<�%Q=�J��]?O��Cw7�H��	o{o�y�W�A���-O��`L����#NDb|��V�Z�������i�<��e8 Ta�Ȇ6%�旳)b)��q<-���Z~��[I��-;��$�@��#ύ<T����24�K�#�B�����hl┈���@��Rr@������$���P�UaV;H�m ���b�L� g�F�Lts���# 8���y@S�_� @|db�XN���ZO���ș�,Y�K����gJ�4�ܓT�)��6Cڤ	#r I'�^t��<X�L�b@����E��R���o�7������!�:f���;���Q�f�:K�sy�V\S-6���'��������-���S���xҺƛY���x:���M�"<���%�x?w�9F�.����Ӳ��VO"4�Œ��Ps�%y�e�M�pz��<���P���$����K���Qm��������If�)D!4Tc��8���*+G�e�|���KUlJ�m�Z0��ｃ m&���k��H�w��Y�G�ɸ��ԹL��w��-�YGһ\����}Dׇ�T�v_�7� ۔G_�����"|��x}��T[��r6V)����wś3�4��#D'#[,*}�ݫ�J�﹡I2��t����G'��\7���q{�G�{��i)�<���+��%� =���,!�:
]𥙎w����y���kEz�SF�t�"K]���<��O(��9�q��g�ؾӖ���"a�5�>���ל���^ �X�Db���=P������?�j%��D}E�䶕F2���c�-s"�K'�:i�����G�|��
�#_FC"���y��/�I��%	%G�K?�j|D���&�dO���H������3����~l�����o��/S���\�(����C��=�^��Wx���#R���Zzs��Ny� ��N�;4!����a��ʠqf�%-H �J�h�
5��N�ָ_����L����s��#��G��I���.��,��#h���8�#�Ώ��ΫO�w��㼥���$|l`��]y�`�)q���P<��or��������V�['�N�Q�=��6U�k+��H{$wО�ԅw�d�lBg&�����5��S�ͨbS�2g��$M�EӤ\�j^1
w��֕�9�.㊃о,b�@��J�J�z��W�rz��Z�ϵe�5�Y�yڋI�a���uӊ4.wϥ?�m9�Q���FX��: ����q�@�cCMշ�6��>tǄ�M�/	T��?�0B�Z�6F�"�7g�J>]X�kY�
~۩�bH�qL�M�Z��H�L���V��9�m�7�ӲI���U��Y��K�t8���+��ۂ?�Ox�������zui�D�]����	���$�-}�o�0�=��}96�=[�.B=�;TS/dey����̙d��/�֐���ݵ2 �W�ɺ`~\q����
�ϳ��V�Ꝋf�s�E_ޛ"��T�T>�h�Du_�>0ѹ~!�pyZ��gs3c���dX������g�TU�����'��u$��΅��qڅ�#�Q����/�s/�#X��'P޾��F+j��u��8���L�^��(�Y�*���^(#�gI!��Z~�� ���A���1��+�Yئ�������s���*�nK#��)���m���rb�jeYO���0��R��4�,�:UA�[���Ԛ)M��z`F��c�ڞ�����V�˔b��v�x!�a�چ�X���D�g;]"��㷙�߻q�1�P���*c�Z �doD汚؊���r"䈦��>�J��?)�x�E�%��E�+?�-�q�����œ���	�76g7Ğ,h`�YA}]?
`0 򳴩~�"����
;Hx�y#sD��Ε�v��,'�N&�^������[>oj��U �ZP8%�a&:I�YW�,N��R}��I1���vGHᲫy��{#�7G��NZQ����R+(��a��#0��׵�<*���^��:��M�<<;kC"֯���!ܜ�"����T��w`^�2�¶�n��[���+��;��mX��x?��}=�}>��n���
c�AP\Z�$^� ��H�ݻ����Ta�H���}�"�����`��
���mno�N�Z����Ȭ�Q9F���^�ZLXbU����n^"Sϙ�yw;�X�tCX��rG)�0GaS��5�t�x=�Y#�oW�&�
��S61Sa�~���4��ދ�!�#������J�- ��"�zP�v/3P=�����)c�RN����F2��wP'%�+ �^]7�?+
�ʵK��R�]�ʝ�->e�=���&֤�0d�.���'��ao��'�8�f**�zD���z/;�G>r�f)�WW����-U*���N�j��t��)��(b9�����wZq�5����I�=N�i���^ ���%��9�~p����>uI&ݐY1�c犔L7-���S�^��\0B9����D;8Ll�T�uF��1ڼ��TF��Ϧ �ǜ�LyO[󨾦�5z�� c�~�}��5�B6��K����U��a�o���Kr���w�+F-6G��GFJc��G��D���9�
� )dv��0����ul�\YZ2i9-��^��6_?�\� ���8�����t Py�~�֕m�jG������y�Uj:����\f�Q��OU�|dh�Q�W�=&��?A.W��2t�����n�'�N�*�D��>N��5���!ɾo���\�$Y�ّ�ޱ�|1Fq��p�v���|������(�!�1�ź�UT�l_�V�hI�V0���
�ϔ�0��&��r#'���i��	��f�w�BX{� ����o��!���Z���g��A>Phy�� �"W�R<[��C�t����m�^&���F�۔�8<Z坢�]99K�ۗ�LUa�{�4.xH�7��B�Q:��я��'���
>K��do��Xy{�.m���]�O;�[��P>��D̞5H�A��\s��E�p�m[�3(�@�J�8���4��*��0:|9�2� ��U�"Vj���yN-f�挵 ��R�uz.dٗ�ph��^t��Dh�;�ýh�F�q�)�n"}S�f���v��-�M�g���~4�$��(�Ҽ�kz�L�M()U���wF�z�����u�]ɢ��������fl�aNuSP(���Խ��G��=�Y�l�n�(�kT}aօ�l�8^{�[p�v�ş�� �4�k�w�TU_!Tf�%�U�/x���� R3M ��Xbr�8Ǫ����h��W�eC,��ߞj��z$�a����OpQ��߆�}PܲI����q��X����#���7�s�������3J}C�ຆh���}"��t��ϣk7Z�f��Bp#�O	GX��ƿ��Gf�5��!�22#Q��7��cD���l�S9�\��HBm>OO��.AK������:�`�ݿ���)�U|-r̅�����dۅu1Fc��٬/b��v�>+���U�54���܎s�_ΚOl�t����v���f٘R�z�Ln��*W7M��(�	%���Rh�ȁ�h>FR��]���!3QV�d$5�+��eQ?�����J��h�0����,�Ż?�7lgk����RB���;�Y����묭!���&P�p�t}syk��:m:%Qg6Ф%��F��h@�ז��2ͺ5�a��w492�·�0b,P(E�,]�IC�+������b��K�8&�+�˧[�s����5?& ����_� ��>R,��aֳ�\f3/�W����;s�#�������ǽ�郱�!�ؘ����7�|��f��"X�Y�X\���(�E7�d᱑cz]iG?�����^-��+`��B���,[�}L�`&V`�g�]SvVW�G�[�6RM�ߏm��5��k�q(���&�˴6�`r�;�ٞ��T`�Gj�>t,���.G
��=��R���|��!�z��[+��%G��+d�Y0L'aL:#UTHO�~��嬥F5-Js:���#������9ȏ2��A�3���Ԁ�bŊ>�k�"贚ZVEa�.�.�/�]����7�G^��Sj��2�;�!�H�?'3��FA��B[긆���;X}=�qu�Ntt�o�W�r��t���xN�C!���4�F��U��ub��fv����}�]�u�~BP���qD�uF�V�}�'}��		g�2�N�A�<��t�y+
�i��ߖ�]'��MY�}���D�{��l���Et��6?�d�bi����}�KM^Y��]ՄGEF�C���HP/E�F֕�6�	H�,�Hϻk§M�o�y���C��l�~�z�~v��ڂ}����Q�8O�wk2�!�-n&x%YC��Mw��p�$���������ީ�v��"��*F+�f4���H�4������;�I堌:�j�( �y��~]�"�6�/4�@$��H�8��̂yM���D��N�/4 ����B H�šl��Lso��pb<���,A��,�kЫ����,]��{��]�a�V̚l
�j�fy�ڀX�rH�����a�W¢\������ngSY��'���`c�;�gU���Bz���{ma�ZݯR��gj�5c ��"q%*U�|p�4��W�y�Q�7�I`[H��c"��
���4�]��P9���]������4��ng'��wC`�/���)�L@����	À��؛��8�'�2���IuS�(C��KC���@�}��#���q��R� ��ɯV!���A%���;�X2��A.��\�����"4£Ȱ��r�?�/�<i��kQw�u��j͝[/t89�x�c�H?�D�Wi ��B�$���vǼ\���m����Oy�Uc�9��IsSǑP3�J�١9v��>�����[��� I�L�nO?t�� }��f�qـ'#�p7'�B~�A��hr���4eBIt?e�Rhh�b��{hm�>�ʜىZ�݃qg�����G�g)<�k�=�u<$���BsI��fߏ��/*b�����p����lv�VE<4a�o=��ü6b��W;��V�uQY'����.����V���<��6J��1@
�2/�V��`���ʓ<��3�#���q�@�>�����)-����F�TJx��-Ze�*9�.��樽�뇖�`��ަ�l�۰NUD�)�1�[�'�_��&�c�Qo�f���I��|-���f���j#����U�tsH}1�D;x$�~G4#~D3�@�"9��	��x��`��D@��ȁk,�Zca�d7�4S#�9��-��K`4�"uO���V�瓞~�\���L�bYA�q�7,g���E+b��n ��˶��ŪZ�S&�!��N{�!D�h�.�f>V���Z��D&�����k��r �~aĔa�]4���eϵ�<���Ao{w[�
f
�����z�ց��v�Z�^H�d�pg	t��ZˣՉx�+�:,I�Zz�f@�(�C��c�W�=`���Gh^��:��N�t1����n9g��B�i�d���`(�����BӿZ����{���gx���SQi4�ߕ��2�|C<�����11�Qv�V��>Bc���e�~e6���@�n�E�qp�/Mz-|�P�J��zh�_�5I|B�W�� W��Q��^���cˤy��׀�f�	�0)��nЅ�g6.^��?}�cU��k�<l�Ef.���Ri8�~�d�+��$j,r��rh�����T�ý�Ξ���h��$M�(X�;�N�eS*�ӕ��q�)�]�M�2�B��>/J��!�쫏h�%�7שN�R�[\'��1;,P��Ve�
�c��δ��[�y���.�Zu�d/z�΄��4�t�{*�Z�tbj�g�u���sXY�K�4eLM�I���Z�8@tr�2����o\���P+>���;�ۅ��N�лugD�q�~x��A[�,���C�!��M��J=��o������\�󚿿��3�mҖ-[,ޢG=��%$��:����m��ݍ�C������IK���tZ�QJp� ��L��ǊX�I�*��4�G�UѰ(5��&�i	
�SP��g�,�a�_�¢?O�o������@-H"ɐ�V��hmK:������V>�y�� ��IKBE�I�ٿ��J���8ퟚ��iR���������}*�Ů��+�M_J���ŏ��-�����S���w�F�eʛ�r�T�
����ˣ��_�)���mM���"����{�g�K"��3Ey]�_�\0�-���4�c|^~�N9����k) Q�*�'��MxA�ȱ=��KL�,JfbF���o\���g&'���L"�07��a�L2��P>*�h�7;�r���6A1i��h�F��� /���?KoU��4`H����~����7s*��ҝ+�rV���!h�G.�8��� �&,׉7+_�ұ�AG�]L��Z=h�ːȶ�Ɖ���$3]7�p�Lf���4� �����XA  |��k|���D��W+<$^�Dy*�Z����oꕮ���c?�Ol�������ʒ+�b�y�f�Fн�*`V̝�Zn�}�$O%Db���'�,B�YAA)�LBS��C@�H1Sִ��v4X�.})
�+�4r��X�����*,���B����*r���}�2����؜̫0��$�л���a�3���W1�5�u�d���Of�\h�𼽀ж���m��a��Ԙ�/ �.PA�^P��2�vO��"f^��P6Rt����S$��nr�G�.��GP���i:D�|�W�ھ��X|}�'&t�1�nϘ;I�9p�������2�l+%LQa�{A�X:�`L�/c�B@|K�c��D��'kV��]:u��
�%���i�֑D������&��9	�`�7@��'ɝrxO!�q���e��E׵��N+�78G{���Z3 ���sQM�!p�s�3g��(Bq��?ۂ[{�Kl�X؇�a>����6���e���U|[�S6�L��e��(N��q����Ϟsi�'����^E7�H�D�JX���Ϲ5��JNyg��j��!8ǀ�<��¡�H����C�a���ǛЛ�m։U��8wjc�t�9��=��Qu��Ȓޤ����Ŵ{�{jp�C�?p���>�y���	���n�`���Q]'�%��r��)d��K
��wM�T<���X�bC�ǁ���Ը���{.�5k�31b֓���z�٨�P�q�C;� ��sM8�Ȇ��|��M斠hI�]��ؑ�w5��.s�8���P��P*=8���pq�q�\KzB�C�JŪ��3���0`lzP4�	iO�v�Igx���g��-�����صY<D���%�|�&�EN�vv�J�1F��S�e̊���T,�ĻA=@�w�n��^N(��^ﬧ(~|�,������P�G�)��p$Wf:�e٤
�(~<0����#^�ޢQQ���� ����. ͳ3�HYZ80�>=�].+Ջv�hZ�˧$�֩�Ei���J�e�G`K��m�T�4j���N2 ����ؠe���6[,�N��#�Ӟ�:����UPxM����Y��"�VS�����)Zv[�ձG��Q���M{����엠cJ��4xS[U���_���c��W�������`)���pP���kT�QF��`H�AyT�J�pL�$��R��.�,���​�]
99��}���@���+�vN%t���I\;��a
	D�'P'���s35��l?j^9`�dĹ���W����V"�`�[I��j,hL4֤[k	�V��U\}?�I����QA���k�=��y��zM�u�Q�J�W=4n�CD_u�ϛ+ d�*=�;P�lMMn�m�� @�75���V�O!B
�z�� �%�\~�YÖ���f"�Ӷ��WZ���XgBp�A-���Q�2C���‎H֡��K�Y���|.�������\ �P�aK �C��e�3P�Y���i^�I�q��;�Ŧ��A��v���|9�([m>��y�%��)u���������J'��;�O�X/�7E"�$0��9svE��S��糓�w2W��h�m�1;�� <�L1�8� �ʱg�8��Tw�͖�w<��Ad�پ���
���u�2�4�����v�f�l�,Q�P�k�d��~���� o��s�p\3C��6mB�k(�8�j�@j0p���T���k��ވ9����,C��:��6�]diHe�Z�*ܱ�.���aO������pP�~��v�X���u�8,pJ��b����ԏ�E��S���ҸF��,����:.�xdt���jl�5��yg��=�
y�ST�x��j��(ڞ��
��y�%��H$�}#�e6�EHb�%�DQ�"1[��th@|,��Bon���H��ۿ>�	�i %�X�o��U�iy�C{>ғ{�D~*�c^����/��r�:i��}��$V�����B��v�.J��3ڧ~�!��0�c�zˉ`M�P���r�|�P�n����M5J=��%s�v�h��-����A�72%��i�4��v�D@��qx���wg��������7&gf�dtMQ��'+v����Ʉd�lơT��U�����ǽ�����DΦ	�?%�/w��n?���k��L�pÉ�뛆�B}凘09��v�����=Nsm�H^��굗W�����g����P` ����CR��w�W���Ʋ��h6�߸��R6zצ>�6=�e /��8�m�4҅��9:�T2�y�R,Kc{�K`��k��r����/�� t�W��h�vA*�V�jGc����%��?�j�l���M��@�Lҡ��G䡹}~�o ��r��VQC��$}2e�d���|�^u�f냶d�3�uB�P����:;=&C�V K�� k)N	�;{�u�Iqb`~��~ZE��i�gR˫4����,įJc����3Nȓ<�vƿ,����N�E�O{;5t��3z��#Ue ���������mTD�l5P�X37�uA�3�&�|
(��l��X���g;�K�Ñx��"�@<p�\����;&z�Uߐݮ���ob?�]*<L%�4�Py����V�y CC׋��J{q �4p譴�V����p��0�b*(%��#�Kڻ�X5n0T�-��
�V{������t(�9��X�`��-2�+����'��2�N�}}�]�)����+��}
�{w�ޭ�������K���E�FJ��5�d�3��zu�Sq~����3�	uZ���� Dc� �S��.G6	T`ڴk��p4�۝=���_W�hn`��k�o��"0����9����K���_�ՀZ9��=x6���`3<ܟei�^�.�:��֞��:.���˃k��'`?�r{~Jn��9��.G<KѢ0��_?EZ�l'zTGX9xi��SG��y���;.)�0�  ��gf�|tAM��R���>-g䉹e��n�f�% L�;Q	 �� �T[ �yXb�6���m��~�JM*�DtY���e�9܏쟠���~�_Ho�N�9)u��N
c�P���
CE�*�n�G�[l��/�ZtȊ�e�-���8�ߋv8��/="�>><I^�"���[~�h4��	X�6������6�?�`��}�]0B�|;9���,�Ѷ�_�����F�=�<�����2{�E�x��J���n�g�lT=�<u_pG,3�V�]��5*����&83}����-�q�(�&G��D$-��$���ߕp�Pi�͗TY�鰔%�f��< کe��L ��ˁdw���~��e�2L����c}Y�T�3�5*�ɘ�\o�Ǐ��{v �!��o��W�B;l��Ҷ�iL�����)ؠ�+�&���C%���Q�<$3fJ=|ɇ�No���D߽Ǜ�n�\o6ci\k�؆��}h��d?��� q9��� L�:��i�ȹ%�I�Rg�#6^�_���d8(#�կ�g�?�z��_w����ck��{"�0pP�*������s7p�^���k�Ա��#��!�[u�	mL�ϧ��r��N��9D�+73���g�21�h�z�PyL��D'cE�8h]�*�݂t3��T��VN��/�jL�j�s�IĽ�<���];�W�L���c����h�	����
�\[9�Kz�@�t�wV�#;�KL��l&�:j	�Z�b��C�mց~=w�9�]D�U7���4�B@���p�����%�D����Ƣzl|�N���6^��9�+�B@w���a�7�J�*VO�Tճ\�š���­VE!�F��<[��CHi�0l��=�
���MzȎ���c;���S员��
��H���a7���{^UF�����c&E����p�������E�8"�-|�a�t��T���H2�V�]8�U�"�)'S�v�;3+���֔��h���I�q{�̘��ȶIP��,身*���+�pv�J*e�"l�^�����&�f�kZ��7�(WV�P�R��'-�4�|&����)��^
,�L3uˈG=AX�9��g�	~o�ɐ�:e���k�	 ����54�(��-w�	L�t ɂ�Z�0���%�>�����YВ�1���@�h�aX��1M#d�q,����zTp�^{�o"<��u��R�u�^���]�Wf7����k�#�0�'��??>}r��<ij�}W�+x]9�ЖԞ���:�S�{�oP^v�y<e�}*T��gj��0���i/��lߴl*"�A�N_�^*ծ�#8��S�_R�9�,.�9"$�z�|��2g_�k,��EP"
c��s�ʆ�d��Ou���L���	��b
l�)G��Yfc���-T[�Y�r�s�e�*�VE�,>��I��#Q���@��;�~���2*��}���@�8!\߃���E��ݦPX&�j����XH����Б�좘c�>�p�"[���z,ʙ�H��h�|jx�����8����ۅÿK|����~�QTZ�MgÛ���Ǎ��*<]�E,*nIM�;�4��zm.�h���d�Z̶�܊s�.�~�n��v�T� PZ�gt�7x�Y�s�`̠za$~gM��/��f��Fĩ�.W�idRJ�9y�0}-"<�D��h��[^z�<S6qw�{��"�h��}�9HXTLwh0��k���	��ө�������]�R�� /��_P**C��_�m����!.�ꝱ� �:�d�D������O���p�1u>��5
~k ωF���R�Y~Vh�?�r"9���x����b����aHr�_�eG��U�@a� ��J8�Y;ESl����ID+Ȍ������_^�W�0J9z�,������]�)�s~ �Y�x6��w���m��smJ�z�#���p�x�w� 5�g�-��������y�(M-�X,��1v9ѐ1 7�[�X��5���i��:�Nۏ�	e�ۜ����,$0�1�:�4�_���<��� h�e&��o��{j���O΅œ� � �� �}k3����z�g�w��̩�#Ç�\����,��Q����Z�'s����Q��~x��A����j�q�qnt`\M q~�Nړ��� ��Q���D���XG����>*7��Ӛ�v��f�8[_Y������e�IF�PI�,M��0|�wS�#���Y��J8��".g�����L(��F�f�!Pe��f�u5Xy��=�����f@�x+YB���̀o̴^h3�XU艽WXF���(���$�K�ݨā���:�G4K�6��C���ѰuTf�k�y�;�
�\��~y�U ^�?�$�cP�w��ٰ�6�)l,��A2K���]H�Z�Y�Ovr�3t� �:(V/��ĉ$H�-J����X�� M_Irwʻzw�셠>8�V8�®�$�c��Ŝ��~?�P{��/�ws?�Ð;:ð���M=�9��?|粵$�B�[���i�Q���&�iB��(��Q���÷m�c��Q���=<#�ub�;5r�Xձ�ĭiִy�n��hzd�m��/��>�9��lCņ畼�S���}�Vz��m	hM���f��ڹYOD��>V?��N]�<Aۉ�.��mFf"��!d���N8��CӠeF�8Ł��y�\ڞe���Ԫ&�^C����� �tض�H�& Ǆ'BZ��@g�i��|��a�3{��!�A�c�nʸ}�Q1R��kQcW7c�x�#s
����.!c�����a<�%�d;�Dwj�1V6+�St���X6�_>B� FBDᾀ�WhËM8�^������?�v�����[�w��(R�E�W�H�C�Ak;�[�X�"�<2s4dQI�����&���#�޹⿔8�����r:���QF�:<��?,�8�q�5���ͼ�ժ��X�.]���V�M4n�q���%�0��2�M�F�x��X�����H�QEl2�9�����A�����Ps��B���X}V&�������=�m��$���y������R6L"iEc��>�����ֲ}���h�__������
�<J�,���5Db@��y�@��|��?�&)����(]�ݼ��k�T��N���(V
O�g��o����Q(�����=����@��Y3e�p>"�]D�Ty��2�9�Nb��N�'��]�v��&���S��!���Q�������\.�#�r>�L�� ��w�
�V�xºY���Uy��� 6D�P����32���1���!'7�]�7At��V�Q7 ���b�������K����2��c�ط�k�?Y}F�%9j���d��`m���}	HTb�x���x1�_C�)��3&�Mb�g�^.%;�Ĕ�?�_�W�~Ӝ��&�1��\�[ȩ�x��t��3��Gi)��u)�A2{�9�D�N6�ӄ0s�I�~�V0W�l3X����=$���y���Vb #����Þt2�-�:U�j���W_g[�E����k�&Ʃ3��љƋz���������oVv#�ΎG ӗf��$��*HA���E���%y/�̧�zX{6 s0����L��j��?
I�?�)H��2:����՘����?f�q���5:���Nk�j�6�1*�S�	V�2�L:>�<�$.Lvi�X)�pc�E	��r7�=ك�e�Yg��#�yQUXS�Np���?�Y���������8M������;��o���p�>���瀂[��[ʰ[i�q�.�6��6��x�u��d�#5�g�0h�^�����_���;4[x�n�&���\�5�^��7��b�D�A����ڽ?�� ��9D|�lz ��%9��^MF���pH����D�(�	��A�Y�HJr)��+�!t�9*�����P�⑭��g�mc�D�N����)��E�dɚ�>��^�]����ry�&�Y*�S����j�y���+��{h�~�n;�2��*�W<0~Ą�e�> R豾vV�L��.���o�y�
��n#1(c�����+}����s��I�C����;������iYx�D�z׽�C���#����6z]GMO(!a�٨�-�Ȣ7oB5F�έ�������Ȱ0�2������z��G���
��D�¶\u.���ꭟ��G��Q;�S��#�6Fu@|�U��& ��-C�c%*�wd���Og<�[���.z��m�E��\�@q*��Q�2�����s�}�#�K�w�ze�[��\��q���[�	.��*�.Fe}m����.�'a«�*������pvdeA'���AB-�&���R���a�c,g+�KBL��p1/�g&rK�b-�ZP�:sR��+�+܋p��`��}ށ�qn�]!_my�6�Zi�C��TE��ͺx��u�5��,���䶣�,�^+lvz������$-}QMj6j@ƫ�� >���<�>y������&�"��=���^=fO!���<����v�R���v�'>�_��í�Pt-Pt���Q�^���?U�vӽ��~�@�M-?n8� ��E8��zxGc�g���٫1p���ƺ����vH\A����Y�tED^իyVf�:��CM�MP N�V�.`�M���}����6�0���G�b���̠�R������),�T�Ŗ�>�{���M��bla3��ǡ�=4NW�7:t��}b�r��sc�;�1��̴5�_�Ҙ�����#C��,(�`�C^��Q,��b� /A&!1g@Q���cyV�U�
:3���5��1ͅ����q��WORr>{��i���خۓ�����9�.���A�C��"rq|U�߃�r��-�28f��1�D�m��_��hQS7�Z���hh���[ �o�S��0C�-������������B��`�e�=AYE�+*�~�x�6�%A����&Xl��"]��M{-��nko��lǵH@�0�'<O ��ęPMiG��C���R8) "~�b�Ҧ�:��� v�*(��:�$C+zF˨��%�ə~��dP��9�p���������ڌ�1�`����maR/��iFf��'|���Bm,t2Jq�`��0a|h�n�Zg&���5�H���ۦ�� ljV��Y���l�|���)� '��B�l��[Q��v,m����0����zG� �f�ho��4Ԅ��Q���h���p�x��̱�"('y=����χp	^�%~��3K���֚����>:�qCUW��|n%	�ɸ⡭�G�,�sn{�zj��	�5К,7%5�+g!�R�����m���t�]��e�w l�.���^rqU�JX�@���iw�����ܖ-Ì�*2�lX r��,�o^U8�AQ��63���Dt�k�.(b�2�YW��`h�&02��\�Ѵ}�pC&�D�/k��������Ԋ�U��T� g�HZGT>C@�7)�W������>�2�|�����(1r��w�������u���Ŷ$���X���v��D��P�� S�=��w �J�yyʤ0	���[�^U�+;���o=a^1�@�I����?�4�� ��ć��g�����z�ʶf��̠����Ֆd��q�'��H%��t}�K"���(��N�0��#��H	R�h��L��C1<��&�=�m�8AB�ތ��3��Ԣ�8$LZ�q�ͱE�a9��4�4J���s-���YѨ�c�?{���+�vƗA�3�G7��*1.�+@�S����_���;d!^�W���s�<�6��,S�8q $V���lr�;���q��WZ߄�\�
��^���U7�0X�#\�+���|E+�</��@��2K�#pS#^"�:{Хd,�n��D,��V�U�+���h��1�sR��#/MwI�2��e"ߺ?��w�|x����r>@�L`(��o�-����F��^\��7SF�gnS	$�wa�IQ��8뾟�B���1]�ܙ���,� ���^�w�լUb�+wu3"�p�fw�ǋ���? �a�j����(�NY���yP��Q!���R�?Y%��6�ٮ�U+�aL����Y$i_����EA��̌��k�T6�%���1���5�\k��	�咄
��m��*�[���&���Xv��n���;�z��'�l��!��A�X�!�Zߎ��ͬx|����\qf3��%�Z�8�In���;X�4
@ �&�幵�,t�M<A+7��:����Z�����:��������c��O �X���#b��S���h \��O'��`�q��Z�b��5�X�;FN�'�&�b���1p�;��K6C1�A���Hм7aW)�!�1@u��_5%	'�$SvN�[7z�ȅ)�%䌩��_����c��
������(ۜ��V q
��5��n�S�*��J&	�����ZoJyX�I�z�I��ys9�&}��"^� m��WS����(�N\�k����6��P�9�p-�C�^��S.ɻ����s���������k��I�4��d�	6�跼�@p�����K6P����5�A>e���|p̖I�_�7Kt���K{���$�*�� #,�RX��y��h�
-���A���T�3�\(���m�[X�K`@�5&>ۇ>1�z���<��ǝS�v���)>�t�T������e��Ɲ���x�[�b�j���̂��"8%�����35{*7��9���d�H����Z���$�T�Ւ��`��[M;l,�c�c�� s�)y������u�	|+�.y��ַ2�'韍	F�U���E��@�O<��nnHi��K�3e����I��b�!� R�:x��� s)�_����2�X��e��K�#�-H���]��r�?1�J��6v���M�U~���e�����=1�։W�;�g�~�R�}�Bi��Xo�F� �I���R��5T�g���Z���ua+��Tѽ�֍�r�"���rn)`��O����B���>� � �Qo��[�+\f�b0>���}evQ~QZ�)�B��E�?Zn����ˍ�$זT���O�N�O6gԠ�C-��F��4�\9󰽍��l|�'�$��j}��a�"�y�iP�n[�M���F�q���L�U���B���1��E���BEJ�z�Լ�a3ioq/i�RۿQ`��KD�+�}�_�SX�#|5ޱ14:�w�a3���b�|lk	F,/%�06bҫ�tU��j!�tu�2�j�Z`[ӗKfj���.,j#�6��;w ��x�c��O��߅ߔbO5�4���D	6+�o��yu������]�=�,i!�%&��������h�+g�H
C�T[&OQN54Y��9î~|��Py���t뀗�"�_�=��=4���ap}hd�Dy�c�	�3�	�8H���������rB7G�ٻnѡ1J�J�����!�������TU����}s��j梅�oT��h�2)�p���qy���	��R�z%�g�d�������{����Yz��2ݻ�d3��̋�x��A��k��Pa�,3x]Z�7���,+�H;�+%�a��-�<p���}��Eɸ���^]!�#�]�@�1�_���	x+H����^���b�eqI�o°�p�Ө�S'���F�w�����l1x�$�b25�j��^9��N-k:��ncۤ/�H]	}����t�F�)�C�{�g��Z�u�]06��Fi}� ��5w�E��V��?�Q�� �Q��a�]���|��fj��"�]�i������g-��*m�Q�x}<��}�<bD��Xc~��)Ht�Hz7J-?�ځ��xM���y���%��tEWB&�X��*|�a�Oo���U��U�F�B%k�p3�-�~���Yxs�=+��f��bn=�v�IФӀ&��|�r���?����]�N���=��t�}����ߨe���D�,}#jڝk�����H�@ ���#IG"[:?���P�x�? 9R⣽镬��1P���iz��uQMv�n(',�İ]��%�N��UO����"��uU�b����kW<@��Ӵ�{˓���_)�D%JMJK?��`K2ȨU?���Ӱ8��X@�E݁���a҄��6R��Tc"���؉��dz0jQU�u�BmA�ol��hX��]w��n�����[��UInj?-�Ow{�[S7�	�0wji��� 
�L�h��?
�f���i_0��4�ʞ1�,ꬸS`$� ev�i�tU�>HΦ.��V[�k����W�{��@5%b8]U����.'��Y�_ɧ�-5�nФѾu��H^މ�&���������ݦ4�h�G�ݍ/�8��E?j��wU�Z���+̗ Dەx9ǧ=���Kx�����*#r�cvٿUj�'��[5���;M�ZI�S8� �G!��[T�3�W3���F��O���O�.+E�罞���B��D��/濎��kU�F�n�o��.�F���������ِ�AҀ��ǃQ$���̷Z7��$̠�T�x�I6�۶G����8�OZg����X3(�] 
����T�� 1&s��k���h�O��V��T�k(�%| _�c8�9�6�6�=m��X4�a�ޖO��Cܷ��W�+n
�@T|/M���?�:��������Y���uT$��j+�~ɣ+~�2BVj�
���m��v}����y�nz�<�?���x��{'8������?�i�b�4�4���:МE?c�u^���k��rC�|q�@E��a�R��B4+4Ȗ7 7��Y�0
p=~WK`%�Ę�_Əfd��5�����e���_�.d������i��8{U��+u����2PɆ����XL8�u�ކ<����X��R=��5��~A��7݃��5�Ե�c{�:��"�֒�YS."e�}��T>"�h|�[1\��~N���?�R�S��'�乶����1�%Ҁ����/�G	�������0=YR^�d�{��y��j}�]��B�$P@N=l)	P��_���o2�,t�5�C>W?�� �Im٣�/�n?��T�!ԙG�2ކ�v�G���>�æ1�Gxc��9�a#�'V"O�Eݡ�.����D���{B�i3�5{���'���܉�xl7�H4a �=��L�"��L�pX�=z)�>�T ����`��� ����?dF��;�c����E��FK�{D�Ug�H�D�+
����z�s�d*-$��j�W���|"�vFBG&���3�Z�H����{��+�"Zoφ򻈐�K����:�o���-|GYD�w�DCX�)L���4!:W�5�{���������
�",)�4T1�T���d#�|5N���ЃЭ0�Q	/Y�l��_��n�C��Kl0��0Q�[�k?]x�A��j?M�@и��pznGeb���6��p,�"�Nra[�����V��$ui�}�?���wK���;��\�o�"��~���C�j쬤B0�T1�m����C_��G{��S_��asաᔺy���b�}����w"YF'���H]�,N�Ę4]�9��<�1�,����Ҳ�r�ػJ'���{3�|F�7>�B���98>�zi˯��� �u�`���䝜���DW;}��8����p+��MAޒ�܊<�oW�җ.�����0�|K��
χ=H(�h��:��/y�F�h���H��)`5��(1��������/*t�.�x&>[D5w�$�n:��6��Sf[(wx��D�hN��b�:T	���W��+��l�w���������u-SM����� w�˥��֪�T��zc���YG�X�܌��f���ҥ��p�0�Q�Q-���0J�m�q������Rw�hX(����d������4�?[���
0��@�)�l9"W�̔�Q�T�7�#,���sb��@o�1�_��1N��#�"m��*����e��
�FH|M����	�Ф��OՑ��0�d�g�����[B���{��B��.y]�9�'H�M����ۅ���pc#��՗x��?�e�Uf�'{|��H/���пMK3��^y%�{8��0�ASi����?�ś(�y_sH�(�ש[[����,�@��|�g��Ed�S��D���ݣ����,G�Q�n�Z��!þ%��7��!(�z���D����b��#��Y��$��?t!'<�n��k��( ܓ����	E.ZV7�e8�$�
�CPM���#�+J)���*�0ǵƜ@��	YyP%�nU�?�p��yw�c9�sQ\/K�ٍ�H��
/�����o��Z?����	��~ۈK�I�FO�
>
�wp�S�T��ͻ�1>���R�����h*%��]����ul���#����%E����d+Y8�!c}�	?������Ԋ�k�cǟ�rR�u�1^��"`�H�����A�3o�Æq텴��3Qs��d���혙��T��T�V�M��$\����딵0Pa����0�s3�
�����J�A��� \�\�G&"��_^�C�Y��\�,�h��ywFˆ��{�����/������<��"�jr�	����գ����a��Q�jcN���~�%�/���<��R�ia;�<�._q�����$>��P���SHx���N�����UVē�Y��W�6%�S� 	0�Gq�z�>f*�_\�Vfl���(�6�t(ǁVݠ{�Y��!\�=#��&��H���o*��������~�������\:I�̝�΢_��akD�]0������ݘ�J.�4AY�)MP����h�%C�ޫ��pȚ����������+�^���/{�Z���>.�6~sQg}L�W*Wp���f,��?;��1c�K�;�b$�7����]1[���R1�g�������{�Q�C��f����tC2Ƹ,�e܆�I�����ޗe�R��`'9t��
h��U�Z
�(��(��k���GA�v� 6���t�{�$^�Q\p q��o|o P3^�xN�6�1"6X�D��l��6�[�~�6gH�M��ϫآ�Guª�/��,��7֙R�̍:rB���Ye0�z��J8�5ל+բL�9i���c��GZ�Ē�����Y��]��@���~�Q���i1���ˁ-���-�+���KH���M��S�E��GwD3�!Vr����Zku k�c֋��D�_�>=\n��p7JGٮW����vcL��6�'Q*~�}����\q�83J�G-y�����>�E��e���u,��uJ�6X���������|���г�Y+B`���� Jj�=Yn�L�l`nqFz�,�A��{�Mٮ�&�gV�*�4F*����cM�lnn5k,�:�}�_��#F�y�`�T��'�S�tgs������;��߀j��m��w2�q�wuB���[M���K�}���TI6����I��@�g'Q��jOx�Ѳ%��q}��Y��/)�Pɀ}л���k"o�l37mh���eW��nœ���&����M+�k�l��I��������v�9��?��7�G�I�/�3����]�No#�(��!Ȼ���1Z����.i�����86�x3�V#&
���R�60Av����4S�Y$���b��"���i	q	µ�f�KK>2o�m���#OخW��EĜ�Ц��ŏm�cg������R��f����5kS32�?J��2�e� ��I+ڑ�����%�_�bГP�O-�}%0�v0�y;��'Gί�=��[��j��9�gOW��F[dWɯ���{ba�i�u���������ԑ�HE%�<��S���Pz�b�! h� �~�1��7T_�oz0h��i&%�UD��t��8TD�	�P����z����2�8Y<�"8����i��k�厐R�~c�<��}�SZ8r]�BWg#aʻ�������5^�h�t;�c���P��zғ�0
�߇��M
�^�FΙ���tWdώ�s	���nue������(�x{��nk�ʤ�ޗm?�-�8<�*]�3!^���bh�GX�*!�t׶7Ns�d�a"{|m5�}@��,��:�\�N|�1=���q�
�Y��V�L	pW���ͻ��ד+�Bb �6�bkЄ���7i�K�� �ˎ��.�+۽Ư����G� �բdm�k�d5���:�=�	� �Rg緼O	���
�|<,���̮)c�{ 4s���qt�*�0ƪ�~-�������;4�;T.��ew:�x64o�B��6��{�+�z��N3�o�M��0E���?*��n�ia�]��
$8�x��V�ߺs$gg��L���Jg4)�ѷ烆[� TE-�����3\��%.���Q^�I-ɩK�9�`%��+��O
y����ބ�P>�|�w��}c:��u�;#V�{��)��Ɇ�z��7P����|��M��U�~-f�o����NVAG��ϻ�ot�m���K���,����j HpxQ�W�0���^خ�k�E���yj���=���h�F�ij���x�EË��Z]�H�L�Y
,7u%Mё|��P�V�u���I��^ug�cu��d���6��x���i��Jt�*�}��<���q%���:qnb��(Ο���w��c_2��Id�� �u,Ί�'��T��P(b����R�gq,�/ݥ~���`c �Q��9KgNRJv��ų�=�
xZ���I�]
}C�I2�C
��{��Oq]�l��>縷�iC\அ=׋����p�e����������PQ�ܫ�4�'��&f /_��O�ф�`�_?����\1 �y�N��NǮ����,n���gr, U\i6w>�V$r��	�@ �@�H��~���*z=�c��)4c	����3������$?빧c<|���7���8��OoY�H`�$[� ���W���0}���xf�4�;�h�B�!2%��g)m�������j8�P�����Cpds���0�{b��Z���e��YP����Y����C��?��HL��� �PL��9���)cWk�eu7�NC8�箄܉� �W�u;h4o7ׯ$���U�{ � `t-��++���	����I1�5�\v焈��r�п.�ͨ\#�]�F�rǤM'�r�,���m�b�2�<�<�xYy�[c���e�l��:�ڑm0��ܰ��!R��MQ>�CQq�J�����$�(�����ِK�3f��Ɍ����B��`\����	�*�k��2���b����+��r�}�H�p���w��F�w½׸hh�(��sa��#N����f�}O�_����W3��SG�]���v��4��k1�;z�R��zQ�R�<B>��Ki,5��O�$���QR�Q,�Z�qy}|C�!>	n0��Y��P��0��1:�p�0A�6�AF��w���#A� xċh�[�k�X)P�ߨ6����T^�$a
� �S��}�� �a�e��vΔ��/�2)�q`��a�Mh� th��M]dU�zSE��"<q�0>پ8��d���}>w9�m>_���^Rn�	n��k���Z���[�^���@�q�Q<T��!"�H̞>U����Q�
��h�3�7����,�ʮɓ���!3Z� �u��6b���lyP�җimĢ�2��^M3#�^�Qs���)�?�f�� ��{S���VKn
:և4�,:�!�F"#����Fe��R����l�d�a��8�dTw8��f����XRf�A�lUC��-��s��V�/~γ�4yIv�5@ۘ$nKi|F�mfg;�rX���]�tl��/�۞��x@e|�o����q��uޗ&~�^ib絆��5�ώ-�����@^��.��'�:G�(fR�Srw����r�Q`����Hs7�>ksV���н��E�����̜Zi{"��a�[�,�x�Y�`���%H{(_f��9�Un1�[��5 ��ۍ���nmn��J ��R�� i���ڎ�jj����R@o܃�~KS�hs����������f�'�k["�_*��ךٙ�-G��L{x�sHGOr�� rX�N:]�-C�rxb�qd�w�M�"�"�_dg�w������Iȴx~�C&�sS��b���+�z�{�tD���XK;�-�}{�'u=�,ݵ�P ۿ)�4��r�cix$x��nl�����v�V��~M$�W�L�����ꟑ���B�OV�H��ܺ+'�1�0�5��)	�E桬\�%�n><����N>+�˭�aTy�Ǎ�E"B�#�a<��%Oӄ}��v%�Ʉ�5�ɢ�@/�y|���V�3+�a@m�ke,C��DoT��y.g�O��(wu�EF��BY���5`r���L�K�Ҍc�+����!^�*��'\.B�����F�/
)L(�	ŚChj��������qv"�����à��Ǎ��a
!��x�0��vvO�Z��{�|����e�-��:�g��R��tE((��;M,��༦�X˶$���WU"{�������|����i���ii��(/M��� ���p�UM��3�/"��d��l����˅���̸`�qCŇ7���,h����%���1�����/j-u8Anx8���؟���?Ñ�R��GZ'<���%#GG"�ؑtu�]���Q�B�"��^�L���Rpu��5���g����wܲ�!�a��� 5��E��]1ÿ}L<��5����MM�~�a?�x����C�ƿ��l���u�m��:e�l�� ��W�aߝ!N�A���q$�÷��"��\*C�̧�4o�E��.SŤ�����8��.���=�~�H����(T��W
��Vk�j�W�FƤ&D��r��5NjG�� �mZ�F⶜��2���Xj�e��H���.]ǟ,�XV��}���oU��q�/F �ӷxz�=�0Xf�D���>oJ��fe����[5C�5�9���ૣC]҃��A�/�#<I|�_�5�%))��ϴ�����Pd�W�Ͻm����:�� X!����I��L�����3�2��f���G�v�C�+TYH>_5�����8�s��l�:�C�U��|{3�%��+q��7�o�N��~;ɠ��M[��<�)f��pb��`W�=��Fv�T���������.*���c�Bb�������&��)��<�%�����ժ3P���W�0'�)�^LH�N�_����
 f�����Q�$�68j}-��!x�\BSl|N���Ǎ��c�ø��������/���y_H�O��{�6?~˪�w��o�~�ў�h>7l�;��;0��c��'�{h�w_uV�� }�w�����+咤�Z1,D���&���:Z,��� �(�}a��w'm@���K�0�#6�5�N�����O$/�@� Zxl�+1�놓�Rw_�h�G�Z��
����ʩRqri�u#�gՃ	���}pV_�r�*�$�Ae��O�a-
�s�5�{��3��<3��z������]�%���:��t����)+���02�rήmZH�ؙ7��4Z��$
�!R��oP�oO�
w�����i-�����MC-/�ݼM����Q	�N>��Ǳ����S�ަ�p�Ì;�����Tb���� V������ϧ��`���f�A��;�>���U� n����|Hm�=i�4BU��Q0[ϝE��Lz������k$�js�W���W��U�Z����"pHV9�A͔�f�$Bw;)�G�"�<L�S2��7��.'������l�8��t��.��v�����S��=u�@�cyg��V�?��T;�}���� ���wv.�ilhl^ӉL����[kӬ �J�eA0'n�T�/Z���\����GF},'g�咍�ک��4���jV&�8�%Yh+�1ho�3���n�썉��8�8o����Ze~������k%�8u=лJ�D��+�Ek��)���霶����i����ƚoH�����DD�˂+�%ݎf )�⩩_��JJ��y�����y��ȕ���'�Z�{ؿ;)��a�y�C3d��3J�'���\�RT��?�>��2}�Vg"UJ�3)
�3=�=1�K�5XD�E�f�{�'�Z��_��Y�b`�,8Pek����a�c�r�)��=q�
�$a=�!8���k�5�M�>�0Z�*^�ޢ
����۽���qC��+� ����Dڍ�f��/�)m�}�����/��۹*�z��i��Ҭ��2���%�V3u��!�s��#�<݌�k��8M��_��k�?����	�,��&�|�M�ϔ?�5Y�#W6�;��|9��8�_
�n�(�rF6�˱�Er��q\A�K��w7c�]�`��u��8\��uG1��d�����1��i��3Q.yk�T
�]o��G��트�����@�o,�H�����T_V���0P���ӧ쯙^
�7EzO��Y�s5g�Ե����Fߗ 2�1�I�L��_��✕k��GЉ�=B[!�H~����ޭ��h��@����7�Hkr���L� ����OUž�.@5'�G��	�����O
��m��6�r�^�MX�����_�խ��a��9��@��uyIn+D�g
w(78=�L2�`�ߛ';��>�ws}�t�&o�2P���/��D-*Pjk���~=O25�l� �dn9�3����gHB���ԺY<l����4z�'��bG�hGj�˷��7�	t7��\	�]!��} -�B?�7��+�Ԃ����7��dߍk��B���/�8L�)���� 6��O��ȢW^�+����(���s���e���y|X�F 0����6s㖽�Վ���	��$�1M��[�A�L����g�C�q�(y8S������bUt��q0%h��@7��pm����|�ؘ9�p:�����3���2�?��z��~�M�塦mۓ �<!����M�ÀI{�BI\q7���u$K��\a�~�(B$�(~F�Q����;ˣ��\�so/��˨�j�[YЏ�o�5�r�l�"���GO���֓�$/��bBץ��.l��Hi�+�# ��Y��#G
9Y������sb�D-ՠ��/;�{.�[J�:� i2s'hղ�%���[Hu�l�"�mމ�I#7O�5����4$ڎJ���iRV]�n���H���B-�WH�m� �

���j��6$�Ȫ`E��̼���ƚ�R0��`����ȕ� j{Lx�#[H�[ԥ��ZaZ�jF��� C�{Ⱟ�m��~ ?b�����C�s�M�b�����`�Ah��8��= %�Z��Q���w��'v�[�-�p�5}�a���#��K4�q!U���MK�0K0�ޗL��I�'?�̩G3ͽ�G:���A�{:��#�,����e/�ŢU��_m*
G���G*� �}r��2
�SHI��D���G��)���� S=4��-c�j�� F7��!�=R�a��:F��O�G+���4A;;%�n*%��~�K�nT`B)���E� �,��t	m�O�t��9�ǈ����p����~Ņ:����;�`S�Q��'�cq�Q��z��� �ЩJe��\�w�U�gtꆍ6�4p��w����?Ѿ�SN�(v�[�AL�ɳ>�����[4)�>]T#���m��JK4Α��P8҈�K��n~�u�g,�ۏ7��0�]}�ļ7p��I!�%��cL���<��z�d�}��-`��f��7����|��p��~y�n\��
��G 1�nQ�ǚ=�ڴ�5��(�� �.3�]��%%:<!F�J�N��s�m��:\�6&��S�R6�nKpɡ@%���(��C������kO�nh�����ߌΏ�a������0�ݍ�m�f��6j��a����^?�ɛ3+�/ؐu�oW���xN����BM���ei+J4$v?Ӡ�Z�c��O����1������G-���"������ޟ��jG�C����s��+�����W�3oe�A��"����ծ춹����u��pB(^��©�o��lz�S��|�%c��k��M�k�2>k�K�#��f�/��;.��sxGy�󤺌��/z�1>T�<�%�[q.	^�_����A' 05*��j�h*=L�#��8���h��|>������_��q��Fq��Bh���S!R8p�1�dWa ��"��P��͛��*^?��>-��(�'�5��x�#�u�C���K�n�J���Y��T���CvXKW��f�J\k6��wt��o̘���vJ�874">ط�'�O�
Mv����=�8�
a�a���n�b�35A�tҀ��$����ǌz��_� �T��$�'+f��JŠ��0����TE�E�XWC��ɖ��nbQ���~ӡb nYE4�r��λe	`f�fo^$П��<-k�d ��>>i,:����#fY�L�m��X��������Dn���1��%CfN��;H귚2)��;����AD
a=I�|��X��
���3h�@�w�;Fn�j����!0� �(f����)6M5 0��z�=��0�
�6�Ŭ뾦�p`��n8��7��	oj@��[���b�> �|G[�����!�!���=����a�G5�c��g���5c�Y�DG�O��!D�?B)�X9%uﳲ�1YrUL{�����	��
[)���2v���*o��?@G���C��Hm�$vs�h�,NFsI����i��s4���5��R��g��W�AX<��0��{ך�NцP�%�.�}X�sL]�"|l�DT?��RfAvKW��`Tj�>e�W��I�H��Ҡ�й���}/�%ЊUHK����R�Z�ދ-܈��&��C����ё���|#��T~3�#�l�:�L]<�гl�0����)��.Q�P�;��x%^�T@kC�j/�j�?�a�E���}�FXC,�(�{qH'�'�=��mϐ}�ONu�7u��w�:��l�]ͼ5l;8��%�'l���h�jy> Y�7������*��h�����DN�#`"!5��;��単Z�d$�7ud�k��N&P�Rr	�d�������`��0�rT�43᝜����	"2�~�-��C���a���x@1��|�/7����Ds=}:X�7��H}}f�K�D8��y���[�|��#�����?Iny[{�죖�p��vi��C�$s���� d�qq���^@t+�����⦙�VA�e.Qg��o�ݮ�kg^$C�f�3��FQk��j70V8�jA���*�@��fo_S9�+�L G���G���L5%�@��	��Ԙ����1�fn������|�82�1:�-Mg�\W�dRm�I�`�Fn������������5�C�c�W����g���<���ik��n�l3���Y��1-�~�T}/^Adqñ󖥜�04���-z|�+���1�e6�H}iT_h�.v��>t�x�k��Pִ�b�d75ɻ/9��Q��
ΒZR3���CǮ^�zw��S�1��zP�.�R�-q�[��h�M���S":���V�q�D�-�����M�7�� L�З�>��p�:�%
����H��z���e�hY|@����=tl�hx�$��PS/Ek����O�q�3�?7d�)�"9X�_a�����9���%����U�?OMJܿ�*�Cg7�YW.V�D7١>4{)��v��on�!�,{n� $%b��l����*[v���OYV�_z&�k���su=[�G�a�;�o�ӆ ����� M��36.�tD�7Գt��V�-�%	s�+�҈����X�%i@���4�׭����m�W�S�)LL?���㶮bCiO�{��@�)-D���nQ䱏J�w!%�%^�4��gQ��Q��?�Cg�3/"HN\{�R-�몥�yX�a��'��*{P�n��-�Dpl������%��rZ�ج�����c2�/��/�9w9K��@5C\S�����Q�d
vB��c/���Ç�c������������D�����d(��Kn�g��������J3~��!��u���:=���e��H�#��,/��M�b�[D�R�Ύq�i~*F��U��Io���F�E�(*����@X^||f�_�o�x5���=�d���m�N6���9�Z�4�j���ﭕ ,���ZV�͉��K�Z�m����U$!���z�9����ب��u��(���8�Q�����@��'n�轴�k�Xr��Ga�p:���昈a��~>1>>��AF��PE�8�X�q �/S�X��a*Iq���D�kU�l������RQG+��|����}QȞW:����.l��2�9���B�f)U�墤��8�m.G�������j�4�ӞB~��B�}���qѨV�D�k�`�>W��l�4CcΞ*�f����� �YD�#��Pf��Y���;��B�M���>��?ZW��u�!1+JO��`Z%S��l�0BE������}�߮�~_�)uk;]���Xx����+b�F�7��,�=�w��cxz����y~��`��EG�3�d?��X]?�Xp�T�{k�o`��9ɒ��	�@�_Lr�yŶ?ů�׌HU(���|���%���ã�A�I�G�����?�Ձ0�䧹-9 �@��~�u�??�%J\���B�.7e�rH�k�y�8hD�9琁���;:��B���!�c�7��<��T�rLJ���Q2��K�In��I3ש���kzz���G�-���_��&���WJ'���
�!�i�O�y�(Y*v�j�NQm�ܶ�����9���DmHc�e��U�����'\����Ckq@�a��-�#��HK�o%�~9 ���dD��Lbp���E�6��a8����Ͷgb	��ږ灡�yJ漀ё}6d�O`���I-�%:��oCh.ksE��SXN?M�@�1�0�O�q� 	���&�!������l�8��`��.q7Gm·/��g?D �!���O��{xk����6т�|�Z��߫:�;�9���ԩ�Z�8��m�t��٘�ciJ1k૦k��Ȃ򑰟�y��E��
҈�XY}-�r�8N�J3`<Jlԡ[�_���iCnj6H�"f[I�mȓpb'�����J��4D/����`�h����$���O������`W3�������U�c���;��Ì�D+q�8Dq`Әzr�.F?�g���4����V{[���!vz%�0���3����c���g~LB��|@Md��~�+歑z?)0���l!�M��m� ��~�ɔ;gH_�$�9�k���Z-h�0�Dc�r'�!@/}�˼^�4(lz'�kN٥��=voۨ����
k!R�����t���P�I^k*D�`��2N�L�������_��M���wۤ	s�ӏWh���F�O�����5RX]�A�	���R��S��+�$����4�D:*d���u�̃ �#��`���<ӂ���Q(a���/�7s(a�1��Y�|s��v��a�|*���t�WueL��K�G���z����X�1�tI�s��}^j��jY�;Ra���z�J)3��ޥ����-B~�D�7��	~ ;���!��3,A��3kt`��T�tM����%��&���G[����x��Eȗ��GpT��}��@���R��vka��V��%�ص��z����LpC4�9�ʆJi�guH�M�/Vh�<��ϣ������M>��2,��?�'�p't3 s,�C5V�,�12.�9Dr:z������}\iv^'BL}��39��V)nvÅ�! M�SÊ�H����Gq�s�_McGF�vXiW�8�T_p��\�@m��)�<�{��Xz�312ˀN�✜Ev�i�週��E?���כ-%��d|z��*j��$a�զp�
sa�Jb������٘Y,����Y�[q2O�1L&�q���"Fa֮$�m���#`'Fv�@$�)4;�`%J�%��	P�a�"�qn�&��'h|pM5�l����7�iְj�ZT�o�{^����e�厂[�g����/'�f�~����C7��l��ܓ����gU�\Ͱ�*���G=��ZǴ�H�g�w�@~St�_�c��1�q/���>c��'*�����]QB��KM����	�g�jQ�i}��r��UҔn$�BiWz����6�eg�+`QP��|�2�Oa���b�DQ9�. b=<�i*�[��C��8��e~�PzNq�K���P�,����~~�˺C5Bg9����N���]R��
��%��Z�x?(�E�|�NЂ��Ф<�wO���1`Ӟ��@/��Qι7��@#��b�[b
V1@��l!~�-s�����a��|kuP�_\��o�������.����EZ�Iz{����'��o�Q�/�.g�'ל&��8����"d�T�]PA7MI�k�U�L�P~��-dm�eS�5{������$}i��7ŗ�O9���e�*t��ye�׬��op�g�Q�LO�?#�����;�<TO�!_F��=���9�#L�V6ۯ.��p =i;Ԃ��*:š��} E�����x�~����vہ���&inP�X�rr�G:|�cg8���ߞ��>潮�e5XW�~|1�)�|pr���G?�Yo艩/`e(���[�u�
�h��㡇�o"[�Z��-F.��+�⊞��1&{�1YʊR9r��/�aB�Ԋ[�	Ԫ��-�o[�1��NK���,��Ev&��Wa�i�����]1톦�ݕ����X�a3�5@�C�ٲ�G^��!6s�vC