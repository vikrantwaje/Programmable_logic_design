LIBRARY IEEE; 								--Importing library IEEE
USE IEEE.STD_LOGIC_1164.ALL;			-- USE STDLOGIC_1164
use IEEE.numeric_std.all;				-- using numeric library of IEEE

ENTITY hwseteq1 IS
GENERIC(SIZE: INTEGER:=9;		--WIDTH OF EACH BLOCK WITHIN FIFO(9 BITS IN THIS CASE)
			NUMBER:INTEGER:=8);				--DEPTH OF FIFO=8
PORT( clk: in STD_LOGIC; 		--CLOCK SIGNAL
Rdptrclr: IN STD_LOGIC;			--READ POINTER CLEAR
Wrptrclr: IN STD_LOGIC;			--WRITE POINTER CLEAR
rdinc: INOUT INTEGER RANGE 0 to NUMBER;		--TAIL POINTER OF FIFO QUEUE
wrinc: INOUT INTEGER RANGE 0 to NUMBER;		-- HEAD POINTER OF FIFO QUEUE
DataIn: IN STD_LOGIC_VECTOR(SIZE-1 downto 0);	  -- DATAIN BUS OF FIFO QUEUE
Dataout: OUT STD_LOGIC_VECTOR(SIZE-1 downto 0);		-- DATAOUT BUS OF FIFO QUEUE
rden:IN STD_LOGIC;									--READ ENABLE SIGNAL OF FIFO QUEUE
wden:IN STD_LOGIC										--WRITE ENABLE SIGNAL OF FIFO QUEUE
 );
END hwseteq1;

ARCHITECTURE behavior OF hwseteq1 IS
TYPE MEMORY IS ARRAY(NUMBER-1 DOWNTO 0) OF STD_LOGIC_VECTOR(SIZE-1 DOWNTO 0);	--DEFINING FIFO QUEUE
SIGNAL FIFO_MEMORY:MEMORY;			

BEGIN
PROCESS(CLK)										--TRIGGERRED ON CHANGES IN CLOCK
VARIABLE LIMIT:INTEGER:=NUMBER;				--MAXIMUM LIMIT OF FIFO QUEUE=8 IN THIS CASE
BEGIN
IF(RISING_EDGE(CLK)) THEN						--ON RISING EDGE OF CLOCK
IF(RDEN='1') THEN									--IF READ ENABLE SIGNAL IS HIGH, READ DATA FROM FIFO QUEUE
IF(RDINC/= LIMIT) THEN							--IF TAIL POINTER IS NOT EQUAL TO MAXIMUM 
DATAOUT<=FIFO_MEMORY(RDINC);					--READ DATA OUT OF FIFO MEMORY ON DATA BUS
RDINC<=RDINC+1;									--INCREMENT TAIL POINTER

END IF;

ELSE
DATAOUT<=(OTHERS=>'Z');							-- IF READ ENABLE SIGNAL IS LOW, TRISTATE THE BUS
END IF;

IF(WDEN='1') THEN 								-- IF WRITE ENABLE SIGNAL IS HIGH, CAN WRITE INTO FIFO MEMORY
IF(WRINC/=(LIMIT)) THEN							--IF HEAD POINTER IS NOT EQUAL TO MAXIMUM DEPTH OF FIFO QUEUE
FIFO_MEMORY(WRINC)<=DATAIN;					-- WRITE THE DATA FROM DATA IN BUS ONTO THE FIFO QUEUE
WRINC<=WRINC+1;									-- INCREMENT THE HEAD POINTER

END IF;
END IF;

IF(RDPTRCLR='1') THEN							-- IF HEAD POINTER CLEAR SIGNAL IS HIGH, RESET THE TAIL POINTER TO POINT TO FIRST ELEMENT
RDINC<=0;											
ELSIF(WRPTRCLR='1') THEN						--ELSIF WRITEPOINTER CLEAR SIGNAL IS HIGH RESET THE HEAD POINTER TO POINT THE FIRST ELEMENT
WRINC<=0;
END IF;
END IF;
END PROCESS;
END BEHAVIOR;			