library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY LAB1PART2 is
GENERIC(N:INTEGER :=4);
PORT(
X:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
Y:IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
S: IN STD_LOGIC;
S_STATUS: OUT STD_LOGIC;
M:OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0)
);
END ENTITY LAB1PART2;

ARCHITECTURE BEHAVIOURAL OF LAB1PART2 IS

BEGIN
PROCESS(X,Y,S)
BEGIN
S_STATUS<=S;
CASE S IS
WHEN '0'=> M<=X;
WHEN '1'=> M<=Y;
WHEN OTHERS=>M<=(OTHERS=>'0');
END CASE;
END PROCESS;
END BEHAVIOURAL;