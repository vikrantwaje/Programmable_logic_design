��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#��:fN�5{�bA1���6B��f�::� �ߒ���1�U�	Fl��T�,�@�퐺FX�&RqJAL�Y�����h2�L��h+;���*O)-�uY���r�ax�݅{r#IX�XMq��e�����~,�+��~�*�D���N��s�"^���Cۅ�0H&�� �8z�7%%����n8ҙ6�.������#��2չ����㡷���<c�&�%��WB�"S�%oa����Px���7�tw���:�7p�3����A��3�l����qt��3	\u�,)̲70��b�-ҸE+bK����}[��!�?�BD����H��(��q��]ŽOtc3Ϛ�<�Ǝ��K{�Y�ẝ�P���?�4�JfC�nUx��=��x�1_��2�S�x�+CǑ����U�X,�λ�I�% ���.��ĭ��id,}؄gqk���i� _c�FYߝH��.�r|��P�qR}9 �,:�M��v�}-X�I,K�D�ڎ��@�d�bþq�8�;y�A��)����I���������2�_��9�+�U���[�����3|�pY���o�/�r�5iB����Ɲ+�,r��΄�v�$|3�N2�.��Lt�K2z�'Б�6:ytA�5c�fA�{F�&��Լ��s8�*]��QI��}�/~��R�K�o�ta1��58�}F7kQ1�熢���c)A��Fb��׬��1>���9W"P���������0/�. ����M��~��n��	�wnv�f�C����n�2d���M/�f�0ȉ��#\�l|P{�ؒ�$�",M��Vl��M�?�����mY�Go���W��68���b���F�,�~0U';��`/4�ߠ�~���VX}�Ŝ_>㺏V��:�����~�N��B��P3�5ᗰt� ������a��3^^V>M��s�)�/�i�yO&e�}�1��>&(>��> [z�S�T�oK&Q�9E��|ʁ��R�IJoP3�0W�.|3ᘛ ���nȤ�8�NKT!��X0�������g� ��%Y�$�,�z��F�@*�.��#�ڍR8H��n��9�Ojow"p8!Y�LB�ooTKa>/�cH���3ʦO�d�y�hc���J۶+���ބ��
������B���YZY���K���z�Ø�vG�V�70�X�|.cx��	��+��,���	-H��5d$��98]�&��b͖�3�<l@��T�����׳�P�p3���̡E�s�(r�&g�V��E�$�����0T݇���	Вǟҷ���D��,���l:���\*AY��J�"�vU>q6Cn^�i()ĭ1!@"�e��I�/���pR�-<��|��W��i9�C��<_ׄu{I����9t��M��I0Gm�������w��Er���R��ֱ�Gf�Ri��+f��)u��NY&�'2��뉀\�7 ���R��3�U2>�n�[�3�{�/XJ'�q�!��/����KjZDy����x�nu!�#�g��#  ��H��m%�v4��	�~���a���{����3�6���@'�+�4t���6핃_W�x@���pkBE[�1+�K�}(���8�7s!�5��=*��lJF7I�L��|��Y
2�BşKVc�k$!�Ï3{�CG�pƳ���ڋ�����c�d�s����/E���KH����`�|�U�,�1�,jVX�]�u�Yl+�*K������V��y���[�,B{�ᛅ�q+K<FIC���J
�0�9�}���u�����/{�����?�����M�nW�-����艸�R�P_C��۝2$�P7��bT�R�D�����EK�Q�C�z�B�S�f���_k'�!E��i��F�1Q�kz�a�#X��g�l�TKÞ�md� ԆM�{��S~�v��j-G� ;b,�̃Y[hK����5&�ß���.��t�Y�������U���f� �+~w����C1'Eܲ����L����*���R��PfZ���0	8ҊF���YETV
:c��$_i�G���8�q��NT9��S9�,R��=�K�n/�������a�1nԃ���&Y��a�hV/ w��sMJ֜��j��3
 Z�J�u��s�$�q�B�õS�&�FSg����٠�O��Ih��O�T�+}z
�|
O2��P#�
�s��`c�=���Z݋���p���m�9�ND;J^*�m��=$� ����C�d#f�ũ���6m�ǣ�@�?P�+�=뵍t�),.��0�