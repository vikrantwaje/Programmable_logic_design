��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2�ǣ_4�^���� -�������u�o�?�P9��!lN��6�]��B��LS����
��^]C�O�����>!��4>�6�PX���g�B	ײ�kb��OB%�Z(�1�e��s�z]F�˾�U@.i˩��4U1���.���|��B�V�����`?���^i�&���)���ya��j� UH QU�F��>([��n��B���ѣ0�om�Jv`����%F�F@J�Pqn���J$�	a�5��ڟ�Ҏ�KN����Y�x���!N�G���I�Jy�a'7IIp��{���Zb���Xd�1��MQ����E�,Z�!{r�fSe�~\a^2(��}�X7�j�xfk<�2tŗ�gCG�lk@��s]�ɼ�Z�:��8����2^���CK�� �2[Z��5v9��a�M�ĉ�:ԡ]��A"" :��N��ԫ
�+/�]�iڔ˞��|�EZ<����r3�)�v��>��=�LS���ة4�3Ɠ�Q�"a�'���6�Q�S��>B��$�}��b=Z��$g{��ԧ��0�S��ْ�)����?u��c���A�·�%\��&�޷��l���	{~x���Q�E6���,�>��o5�q�_y���p�ӫ�^<�:��]_���a
Yk%���]��Q�k
�9�zK�2p�8g;K͜~t/=���lӶ(���!�z>��r,�!l��S���{E0�ϖ���eo�u�-&b���v��IIW� ?���� 6斯B)��u>xDƆ�5H��j�Zf�yH8h7.�m���h�RN�*�Oz�
\܁�� �?䃗������E�9��t�G����k}g��˱L�7+�*2���W��6.�A�y�S3���	f�ϫs�Ws�7��Z��e�7MzL&��7(��l��w�\�E��y<����s�W7BA��9�r��O���}���H�y�w�c���/�����G�腙p`�ۚ٘�v߷G�&�����~��I��W]��r��Ρ�#�IB�*6C��Gl�!������̍������[�����+�j��q.V�kVg�H�2(�,A
�m�,��C��k&��Nj�T�5�ߍ�/�~ENߦ���,�x0�%[���G����X���� L�V).x�,��:��v3�WY�;�B`4*l����6��6K��|Bd`�T1����b�I�_�գ�5�.R�ȅ$�y�v�j@Q�-0����&�vV�@����Vk���\�xe�+����h�*����8{��i�:��c���0e�����W���P�
oE�d�]?t�0RZ6��8�_JM���8e��?,U��;O�,8�xQ�2�S� �i��b�����j���rh����z!�$�+����b���⠫=�r�o����V��T��uӻ0�� �O���X,����hJ�G�8s�Ο���힕Y����]�
>U}ry*1����.@�bm�}�����6ĩs{�d���U7�qx�a]�+:��e�w^�/4��5����ǅ�a�&K��@�	�QQp�5u�3'7v�g��T�#��Y,��Ău.4`�`o���Dw���E�Wk�p�����u�0��$�U��zx�2������X5�T4���z~�ij��5���5)&�j���qW�sS��v!<�g��֖`[٧������.hh����k7>}����ȴ !���0���i'���B�GA�SJc� �~�ީU��b�	���r΂w�ͩQ㢤�9,ye� J�)|��)�ÿˑ�Ęi1�����a�d�S�����s�'�wr��?�������Ԇ�C��C|^D%#
MSB� &�$S�wjg�zNVz:WesX��]mcVW�y������x:�ُ7��l%M4�_�A��/H��د%'`��0w��Z&���y�������;aк��Z���HK�wV��T{�o�1�����9�#w�H�mY�:0L4(GDc�4