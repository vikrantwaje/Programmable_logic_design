��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�����uK~YSokj�&�9ȼ�P������şd�rU�gb�nEg��e��`�"9H�bLr?\��~No��6�[�9z�=�'�곙���K���Ӿ4��:y�ۖ��nż��k}q-��&���z1HE+�j�<���J?���&Ą�p���s�	��+"紒�Hb	 ���5��G��r>��T�CF�/�ݸ#Ɍ�td�M�\FxT$��٘��ߔ�M�"�䮤�Mt����  ��{�������]������
�P8��z��c���b�S?�*K��O�~b�*����}��f^鎸ݯ�1ꆃJ��LG7��;t��G:��r���b�c�W✡p��4�����d���8Րq�������������}W�&��tsY=�$�в�L:(��g	��Yi����=1�-�u�Cmb,r�r����S����F_��KowR����tC%�緂�Þ�x��n�g6��~��N��h^_�1m�^�`��$$8��t����s�r�9>E�a�++�pbr�^��	��V�4{+`a����?8��Zf��Mp
k4|�_D
�V�9�p�]R������Ê�q�P�J)�ڥ��0��#p�Cc�mtbY�K���-8�m�e���(RRk�\�����kY��c̈́
ap3l��t�⣹�awo�T�xYt����w/�US����{��?����à�����$ڿ!Y���e�)�ЗGC�A~}�$�x�F�۞B=?�0�yd ��H�{�U�V�S���0=��r�rt
b>t m��[�Ѯ[Ap3�I���{��?
T�Հ)j�����4�9��?�5�n�ɝ�~j��J�`�I]���Ծ1om�KY/Yq!v��Z��[k��2��������Z�d�L�F��C��1��õ�6%P�A�4�[P��F���B;m��?>vnF1���L��{I!�(�, ��%Z��4���/~�����ư0Z�9�����#܌���uw�3���r�钢����T4B��������&{0�	�� ����hk�<u��۪TTd*D6�MH�9��P�%t��U��M��j�ԅߔ7�/T��_��c��?����uq��(&a��ǈQv�.v��CyCn�����*��c�'f��P\�,/bZ�k��A�n�'��ʊ[{��v�R@�K�)r
��I_z���j v���y�������M��4*b��f����uG~^x��,
Þ�)�Ȟ�Y����f^������$~�2�&����%�¥)H��cp��7ѧ�43*Z*���,��5���I:�;�/xlF40��]VD6zQKDWl�$��"�s/��0����#�zcu�-S�1tB�9Mѵ�%�>�T�0��,��峨�}�����9sB8���J��c7x���<�Z���\S�������.xD�#�zʠbƮFEv�8P�T9fo��hQ��Ru�o�;�÷��ظn'{i����`L����
Gi�j|�1��F�M��F�D�ۈ�'L����~n��l���켹"u��E�:�Q+$����t]M�M���<�(�r���h�cH�#���AXaۆ�o��xت��v_�I
?���M�_g>��"?Oǌ�A�n�Ó�����=����l�:��-���<�J'����=��2�V �ʷ�d{	��Z�G�."�{��yx:�4X'R@�6�<�����6_��H[H��l	̸e�&�K�w<�P�Љߙd�r(�/YX��W�&��^>zG��N�~��Z>��L�zb91{${c8�p��\| ��=�#U��A#���P���r���\/�p蓚XǮ|�ٗ2�h���k�|[0⣻[zE�ʆ���:���is��'�%����e�-�]9C�Nܹ�є���˸ϟ�7�0�/�6�3�I��]rP\Ե�����L��9��$������n��͔� �ڦ�"N����M��[��0@���7;�Ի��Δ���iLA��~]��5��L��פ��G��.�T7Tn������;J�ƺ���1����|`|�m��I�i�Q�ح+?����?z�3��w����"w�<���{l �<�3�0I���vY��$m	�nQW�!I?���c���"�a��/˴�]�r6�̈ۮzk�4��^�2ZLWO�Q��XAM��ڦ�i3��W1��}� 9f����1�Q���Y?���d��E�u�G$�4��Z�;pjR��Tt]�p�����p1�����t�jn��N�b����X�<*��9���%]��¦��� ��n�Tc/S��ҿ�EW�@� &���}`T��3��)�w�Q2<Y�����J���U�%�ڻ#�D��	�P0S���ť0{AU���C*]qH�2�\U��3��|�֊rzW"�����(��p�s���P��ʸC�0�Yu�����j� g��Lo�q}���8��Ա�I.l5�&i�*�{��,��W	sS9�zr���'�J��dƽ��!����)ZN��:�u��ُ:��]s1g�B1��Z�d��,��
Zz(+�%�sj~x��L|^(��6*Q(a���2�\ę<3pF<W�N��R�x��
gT�Q79�]+v~ tu�P�q#c!�dw�'�%�ԛ�0�ԧ�s��e���`�ڮ��x6c�������������	q��6w�H'=���_��#i3��Y2<��W��Eh�����HDdp��%���.jx�O�$I���s)��qe�䪑d��c����,��?�~�2q����jH�������u��NF���;���#����ϓMD��g��=|�s����:���%G`N�'y���^��	�4���Ny�w
��{�B8E(2�qUz^Ӥa��fc��rdu��/S�E���W}�?w=��"
~��}�����0��l ��%9֧G�=ʢo!��xOM�X��?ݫ3��%�E�eZV������C��j�����LLɪ�B����s6�iO���~����+�<�/&���Y��fN�qo�� ����Z�p�~� ��H�[��G��RI�!�v�����L#���5X2Q�@L����p��r@o�v>p?�|$um��yL�]%5�I��hI�hw����%f=6��5K�S�V'B`ǽ����F��A�����s�^ �����`=�f�#�V�QU�0�}E�]8�3�d�N�:{L�u����e�=-�^2�������I��sب����c3�8���t�H�W:��\��-0>CQ�`�(������s�|����lq�%bpU�J��f+'I3Յ��K�~(.�B����<e�
������,m�" ��B��H�z0�l����dX m�fd�O�/2�M���)�"N��,w파�=/�
�1SqW1�%�����S�<eU�%�[�}V5~--ϊ��ls4�&�BF�RM�u�b��t�!�c&�u\t��"1_Xx+̈�A��׷$�i� !�ClA�6���y��B�K��۔9��;I���K^�کv��w��	ZE�$ �;V�����H���v���z��ګ��Wȓ��H��UȄ�bL(�%��"�̈́f��̪��~�q*���JNa�leV�WtER����^�mV��������e�~ɯ��ib�
%�,+�����= �X;��$�VK{֘��&�������9�:��a�(ӣ�����$]�<U!�>�S��;�ƅ��T���dw�5 Y��ߤ��{n0�'�F[��n�r�I7�?�K>�8��wO���	����κE��E�ƶg�ƌl��;1UJI�\�A{g�J�(%��w�ʀbNL�?{]��5W ]w��q4��F��^q�������櫚}2��X+�K��E�����74 ^]ޏB��	���@V'6vP" �8���� �~9�#Í��y1
^�h G�u*ox�Nߙ��"����4f�X�\Dj�]�K��$�zr��[J5�폼O��0s�ѿ%u��r���
ړ�F��G��r��'�/3���f��U�7f:~�M�U=��u

Ѥ�Y9��Q�11.�O3gۘ��@Id�H7Է��@�C����S����nY�B�K��V*�b ����	�h9$=��g�6���i�&3��w�a?B��]�6��aH�G�K�ˤP���]<d\ȉ�����C��2m's���!^q�f�4�� �� �+1I�^�t����Yv�(3��-dv��\V����YS��iQ*���ɲ�n�հ3�I�#�7�`X}$^�S��n�<���p���e�R���>x�����;(�G���;8P�}$�{Lk�3�Y�\=W��f����L�_�T辬ЪW $���^0DH��[m�#fuʾ��:[Oc=����-\���f�� c��8CJU�t�	܍fQ��x[�O�������X�n�#�[p�(��[o}�< ������Mh+����O 0;�i���14Sڰ����b�>6�ܙ�����%��J��-����@�Ǥ�yY��N��d�:�ү�C�M~��Ǣh�ک�\��᫮")�I���xW�,�Z�i��4���'��.|h���KD8�Һ����n�':������	�nJ���*�Ҧ�2���p�*�v8Ԝ�G^R%W�r+��F�Q�넄����Wb7&��V�l.�3{jM���[7.WJG^'b�)�r��;@���`�<�b�C쟜����8��F޼q������a��4qԌ�a��?Ι*�6�l��w��s�m���fy��?Yx�f��4Q�b��܂�3&���ԇ�:G+ܩoY [�U)���m�3��~\��Ql` �ۥ���=�G׼��2�{W	��>�l����?n�LEg7��E����+�T��5�()Z{��q-Xb���C�fM�e h��M\�^5��'��1[��N*�gp�ߟp�/����u�%W��z�{&�2����!R�b�T:�DV,��╯c�On<J2C��s-���jϦ�jz-inK4��$�)�,�1R���Q��0�
���W�3�1׷�/�@+C�f޲(�*�e��m��h��֗�Ʀ��c�W���֓��L%�?<�`նq�ܺnE�X�bBw����h8]gwnN��M��k��c��C~!�B�H��&��Hؚ�<Xr�m`�k����#�fi�7%�����cH���PL鱈����/�ǘ]��G��0��q@���P�4P_���A]�m�>vЙD6����7��Gƶ=�j�m�fɺ���t�ܮkT!������VeI���é��zy~Y���[�ӽ4�b�H�B��mH鯌��!�����ה9�>�y������ѽ~c���"�S.�=
}���Q��WD��$:SGp��q��q9��Φ�ۡ~ʪ^�5cIk�f�9	�� TN��Kw%[��5r��F����q���l����7��|�]�B�V�';TN|�C��t[j�D��ܸL����?7�um�f���f0�S��a�}�v��#
�3�>�V�z�YH���)�s³�p�M�$�c�i�B� [����zI�&��g9[e¸�@Y�z��1}�zy�J=����L��!��e��r��&o��I��A�Mt�5�	������U�߇�
�^f��r��}�E��1ܭ�p�b ���;��v�ӯ�<��(�Zb �u|W13 w���M�����9�_EIMԈ�P�_��T�(/x�=�}oKc� \� ���9lY�D�]��^���#�ƣ�J�>�p�m��-B�ϊ
p�Ǫ59�#�V�B�f�-��2�Y����Qp����a�u��ڒ��L-\��<�u� ��uag�@	�!�,�>��h�S3K����p�qЖ9��s��@/-�o�'j�ř��z._ш.�={L��'�I�{�z�� ��}+�CS��L�o\��r	�6c-�Fq��3a��PQFE��䫪�hP$K�Q�óOE;�QO�#jwɓ��6r$|���'��D��W3��\��\���m�lcp��֟��=��M=B0&Y����l��G��ʑ���%C�Y5����0�PP=�Y"�u�z(��C�.������s/�Z�a���euey��S��F[-��{*{�y
��N��Ikf��k
fC#�P�)�E���'rT����<�,�Ϝu�tg���+�7���NEeû+�4�����5�)y��H��9�U�����J�Q��?l���=ʻ���u�ܯ�	Br�Ăo�O�.�R���g���i���@.M����P=�����<��d��3�ȵ�2aR���܆-5^O�3�
lѩ���`�].�u�l����)s�t�d�Zx�a�7��ve(�~<���N�8�ĉ�E�f�8|���$�h����b���k�k.֔� 'x(��0���<�]��(�.~g�ˡǆC%
Z��1;"���].�,�S
Z����eI��7�
`�JI��J�@��ӂ:�[c���(���3�/ks�fI���������҇�
�ho�=8�������yG��n�)�%5b�9�N#���9^�e��d��y� �D:=��b25�6�G	/ZT��G�CH�Nh�f�-��|�[�4�8emF�  ���k.����)A%Q�c��jKA���\Y������frxS���2K
r��߻��8!��*�FI��m�D���%��`t@�䥵��w�A�Wc�5A�#6=Bī��SO'C*�)��|.�f$��E���_s��9�Oǚ��.c�"�u���Jo��x3R�h]ū�P���xvh�eWFТ�"��	
%ToR�ijhR�����+�P��ϗ���)�������k;x�x�fM���!��n��"�(ז�$l'���_�i��]�T� ��]$"�Γ�E�������YF0	�U"��,��
��6��(�^�o��Җ0��,W�ќ������ȟ�_�'	��c�g�7��6��!��ː�`[]�	pCLߤɪ^ h\���ᷫ�r�{��u�@ΐ�~��Lo����P�r����T�/�LaI��a�W�0�Ô[���R����OOI�	�kAYW��)�yM�4=��hQ"��B��Ae�E��t� H�8¬�S�K.L��;;��2z�5o��ro�{ g��j|$�i�.dnWe-��̤ԭ:mN��|�>���o��������0��@��e	Y�ΎG�7�����?��#��w��_��MkS��,����p��%9��P�Z��;P�{������!�ٯ����iu��>y��H�� R�l��ލ�X)�7�ʸ�2,��B�'��x4�w���q�gf�%���qL���3�[�d&ބ���<d�q�+ �F>�?
�ԇ=֝�{V��H\�����5;��+��h|�Q��"�wb�g_��'tb�P2>T_�|�����m�"b(�Q+���؀��g?�PmJ;/L�Z��D�4�;M��x�Q�I&�R�ZM��Ś�
��6�hL��3��4,���w8�\Ie"����iinI�)�n���Ou���8�if^�ģ�3�yj�`TjA�oR�(`,�#M*�@t��t[���1���p�Y��,kN|h0���7�M����� ڙO�j�0#�}H���y����ф^�K �/Wk��2M��s��ը	>����K��(��}�Ok�)虛��jvӹC!6�����a���V�5����.t#��5~��@а�G&@n��c� ����#[Z֣8sԮ��*�$��^���L#�uk���l���r��N�C+ˣ�T\e,�\>-�`��_����6��ך}��.�C��xÀp��4I.ia��eM�0'��Q$(u{�2&�����@*�'�l�ܠᝢ��
NX�ﳬ���̷��gG_
�jOY��1+Hw����ss/SO'��v�������YF%J���L�_����㸨�x�#�/�^�<����E��~���_%,�nւ�TB�ǉ7Ɍ;CS���=Ҕp���S�9W�Ǧ�Ȥ9��<�Lz!}��v"����:b(\2YN��R4̟�@��^��%8C��ҤL.�0_��,Az�9��u
����V�W�������[
ϳ(�8bYf�U��2��w�xJ��5Ԡ)]�Qw�'YJs�(��\;��)�<�-7�@�?å8�T�p!8�&ud��W3)Ld�㈤eP�>L�ǅ�wGM��+}`5���%	C�,�˛�3�e�y�~Je���-�W��%!��5����B�T�O�;S'̢��p�2����'׊��C�3O[�AB2B�7�V� 4���ŉk�����:�I��xW�l2li�1�v�q�'���r��w(0I\fTi֘]K�_��tI~X�Dߟ����,�r��6(A���O@��һ���)�~�T��
��]�c�I���K�lڑ��@�Qf�0�W)�c��a�J�@8��q�J�R�ݦN��[�(GI� ��蹙Ve�/��zJ!6'���o��!o��*h4wA����d'�h�t�U��R���J/И�+���q��}�E������q��O���eyU�%K���p�L>�M�����m���5�/U/���!����5��%K�{a5�*w��y�J���di����)E�'�-�>�L�|(Qq����6 �?���D�-�'��B�1v��`M��3���F~�BЌ��W����5���x�:����A��r��D�G��e��~u㬹���
+�����u��kb� ����W$�Ć	������ųv��lC`�����ozɢ�c��M������#�)��zp&(;�(�����*$�i�wҴr�ߵ$̣�{�|��B�nr���6��3�<�V\N�fq4Z�|���}N3LS}"�G��f�*����Ա}�vlFD �%V�ǯ�	D]p��=���*�Je$i�ނ�GQ���A���Ä�_=��Έ��>�eTo����T�,Bi�?�}3��bX��	�6�D���k��"���kY`�2t��q��Փ��Zh@ͼ���4��#ck�K�r��O�o+�����5E�����ZO?���96��7x'y��:��H����$��CY��Z����Ӗ�fɩ��t�sX���?�N^��;��iOy
o+-M�Ӝ��PY�;e�i��r'����g��J�K?!��[Z��=��w����Jz��k��w�^�ԌkNʼ+y�N�Dձ��1_@��)�
����Ș��<@��޶d���;��r q���bojeP��;,�?��Zs"���h,.��4P(ܵ��;�Ɖ.9 U�A�񰋵C,s-�i
��^.{s�(�q���&���)H�}d��i'Z�|0>�:�o�	��`[.e�f�Y�2�"����ff?5�b$����!$�z,7�ys���e�px�Lfk����"6+T�N��oh��*�:�v���yI���5N��cBS���֕w /�-�8�@E�E����$��}�������:��(�;�Rځ�\�%ʹo�ïl�B�!�Kc��ރ��su3�����L��Ԉ=����S�I�^ʹc|։!�QQZ��0��*B��H��|5 �Z�o\
H���ek}|i	7���%G��p��M7%Dg���Mѱ=���vYw�� ܯV�^�n�����c���xkZ%�k��Kg5����ҽ�\%$�@o���(��9MK��ȯW�i$&���dN���� ��~��풳���ܬM8ơW�!q�����'A4#�qT�[d�>n����`�S'P+�wȦ�!T�*$f���Af֙=���2��΁hb렬�*�
.�<�T��|C�\�¯*�W�]�y�2����?�aى�T��xG���W$cѕ�ܬ�ג�3Q�[�.�'�_jĠ��e��gp��g�E �[ZT����˟�ګ>g�t��Dv��H�d<�f�����q�z����a��vVj�T���h�����g����ƐV�&'#Y�v��u���Le�ɫ$>�N��L��o�I�;���P&\/������ZKJ��i�IT��ڦ�)h�@L��D}����e͙�e����Cz�lY�iRv���~�5,Ｙפ�z�n�w5~��+���͒|\ȩZn��`gm]1>����V�v���#7؍����Ϧ�(�_c��y�)�Co!�qoۮӍVM��m��ǭ�m}�w�6�s��R��·vO�ᩯD�;�o�0�<���
s`�����NQ���x/����b9�c-04a3����]��O�{��%|��&%�</.j�UH~q&�y��RX��$i���$|4j�uv��5&��n�>�ӳ��~+�q s��9̔]�3�n'"zѬg��i��CJ����g@� ��g|��z�� ����'y���9�ip�Ӕ�}��J���'�6	]����?Wŕ�U}�G���Վ7'X�#m����e�s�.%�^�snK����9�m��?��2M��>���X����	.cn�EL�U�$�v�UC`?���Ty��|���S��U�KR��1D/q�%�@I��'��#+���_dc�|(F�~�aԺD���M+�i2��Cia]�ˈ��N}��W��+���E���j��P�\)�"��З�s��=!�eI)��v#ؕx=�SA����đ'�P\��$��y�� l��g��ǉ�wܨS��O��=��l$_�Q���!\�WF��d��ec7^���p�]~á���TN�e�l�H3o!	:�G��2f�4�:�x9�7K�;��A�ZX�@�0�;��k�ei��0�����IyE��M���XH�yF��l-�I_?�?Xz����p�8�*��W��M�n�1��{È �d�A���	���vw2~�+��4��O���P�x�~�pݚ����0g5B���'� �����~�ʩH{̱� 8֬�����$r������*n�^7'�P/NVbMx�&��j���ԃy�o\b/C%ִ�bgd����I͕ �ȵ?N |W~)����cKa���tRZ��f����<��]����*�r�p��.B�+�@���飯.=��t�aW��=S'1o�i-A���� �Mi��f�⬾�Y�3Px`б�(�0����w�y���T�9���*�i�L�rZqq��G3��p�z�����:m��?V���z;��m�pޯ2����JV�����IP^�?�[�*,�� /"���V|��2�~sm6��R)�mv�te]�j ���\8���Q롗�#�����{�y�q��a�b���K���T� g����}�|���M(*]�)5^I�� -�F��r���Q�8T���o��D(�}���EkK��+ż������ŷ��w�p ^^d
@~"�-J��Jevn2�8K���_%Yo�V�x���:ΛԽ�B�j꽎�);bGE��u���\��v��}���T��{Gݷ������<R���Z)�%δ�b�C��@/c�H����me�[�o;l�I�@�,���/���J�Y	f�C��:w�����uj����]>8���8�ޘv	 �U�ۻ �cL��������{i�|'9�^���j/g΅l��	��#����{P�ڵ�Aʰ�~�?��,Q�ᾲ"�tԢ;0���tca��?�kv�}���.�y�'>��G�D�P��-P��0롄;�i
�,Ӝ��S�9���G0p�h�w�<e���ep'�r~����Q��Ek~
al2��.^�Gv�8�U�
8B��^|H��T*�-�®b�)����ed=Цƶ�?#��Й�$�,�߬�Ά6�I�3��3��5�"��eͦXf�m$O�"����n�|�������0z���_�.T��b2�^B�	wB�aVR��Ќ�j}W8χ���#�{��D�ٹ�q�Av�}�O�BJ�\�pX��0?��,e�꟩Y)���u���#�EBH^0d��5�?�4�C#���T҉�	�~�*1=��Z(�aO�~�\�ݭ	=�Up`���k	�� �Py1��-t�����c,e�3��;f�b� t6��E,-i���)�_:�%M�S<���t��3�N����U�˰�e�*�|�����G��$��Z�����R��T$O�" :e���l�DT����H�53�LhXc d��p�i�����8�#U�1�BHVp�B���ĕ\mؾY< ��m!P��)�D�u!߉Erx�AoDrW:w���qk7k�;�Aa�T����ڬ%�e��E55P9�jRu ���CǞ�����=I�Z��A~zZe��g���ph8���dR
���?��Y��:�U���N�;� �>�'{��%��^�V�<�h�yp�L��8��b6x
V�X���ժ.�����^mC��h��5��=^��x���g�-|��ۊ�P��"3�s�hq��ܔC�2����gք�@�紡�<��ԋu�I�� ���E��y:�7�D�Ι:�� ��.������&r���F)�.3\%�܃f��K������^%K�V`Px�K���$E�E�ъ�Or�{W���h���,`�/3 ��ݣ���ګ�7��B��s�H�U����ܞ�v�il������D�Y������ ���h��=�Ƒ ��K��#,�ɭ�p�)��
��}�^=���Z:F�Y@�-A_]�3a"R�U�f۸14R����H+.S���F<YJ�p���CSSo2��3�b���@��&=��ip^�==�%�՛�3��N��yd�������%/ޒ=�{߲���i(� h�U5uS)������Ό�ç�]A y�-D���qO#��Ee��wΘ��*w�l<�9y�lTj�����K]6"��5z�c���x<���u'����:�&8,?-+�駤�n���V��4��?7o3����p��*��H��)�����#�b8\%�
C��Ďhd!K���Su�
��z�u���,��z w*[��,eߎ5y�J����u��2��}�z�wX����a�@M��(89�D�����ą�A�>_oX�Q�5�i���VO��^� z����ք��D?T�f�n���	):rN�Tq~,�X�N���*��>ļ@y%�?���!�d<��÷W�T9��EcVBd҇�"�ZaitX(��JA��q���m�g���'�"6V���:~/��E�PpEPi\{�YrxDD\Q*V��<7O�Iy�U ���^.%�%�zeu�B���ߛn�biN��@�v��\�um�W��6�������Y��b2�|�w{ퟢ:��3���=icc����V��O�����7.k,ςJ���P(}ڽ_ eC�[�d����P���tW]8{�T$���<)�tx-=e��'�R�i��w�4�3+=�`��|^ FU��4MU66tj+\]6cT��Aۆ3㜩G*����7�[V6I]�V�DF��-Z,��ZѬC���#��S�P�ѐ��������� ��l>?P2;��.O�� ��rvh,�Y�k���/�ͼ�~jl���������x�k�P�$��4�I��%������wL<m�����c0H�����i�����_0�܀#uL�B ��0�:}�9X.�1+���Ҧz'RoN9
Cd�ܣ-�G�b
f������eѹ�I��w�����H��3��N(���+�E	��v��$�z����AK�VD��xC��
�UC�M2Q?��ys=�S6�j�{T��P������n��X�%p�2xgO��P��jOIh�X�)ʈU/�e�a'	�%���lB��,es`W���R{��fh�����[	�I7�_Q��D܇?�J�v_����rN,���d �����J�Z�TZ����Iq�J+to	,����C�cz�퐏�138kI�s�]�?��H��q���x��e@�	�Ϗ�bW@Ƈ�S�`;{N��R� ��7	U����SA
g)��^'Ψ}c3%��3�a�+�GF%�h%<2�3w��{k�Vzi^�
H������,n��_M�^vp��^��tK'|�Z���ֶ���8�~IKzt�9��]�G�qe��;�n|3�9	���k/w! ̭p�z����1G��_Ы*�`�B��ej� @Mk�B�D��H���Aʻ��HR`
��sx]S+3o� ���~W��.�i�x��\
�s���J��2�U�~����H[��3��i�2M^�g��`0AP�JV���Wβho��?�l�nȽ ��"����+Jz���~=)U���IN!i�{\N��C��:�qO�h�l'c�1����%LQ��(�&����̿��6$�;�Sjyk*���wUy�hi�.��^�K����~ă��E}��� V���yr8ӧA��f5�gcd��ʮ�?(�.sxhH��t�x������P�DF�]}U��]�c��q��}K�E�M���l��,%E!����1w��J�P���(���)e,� �D�}i��	k�+������6>����G�N���<aݞ-���K���L���ĀS�\V�/�K�_�
� J2�1tż��f��Pۆ�{)��W����8He~H���@�[d�[Zm����Q�@�@2��ݩ��E�*��|����mHi
�$:���E�*(rn��g���D��_�&�J�7��hF�/�{��������z���B���% �t��~���ɒ=_�_X��WNA�i��^�A��{�y�}�S!�J#�|I��,��3���?+*��{I7�< �Lo����-�~�)���(ِ��o�I��0�"��,�BV=y��0TW��a�o��}Þs|�'Q��Y$6x`� ���UC	�r�&�٫Ƨ���^4���<�S��M�&�����$���t�c}��������n�r �w6�����y[~=x���-����������-�-WU]�C����*"�9�+�TT�kH*�Yg���C;Ņ~5�]oX��
&@<V�m[�y��01mz�{Ȗ�U�Ҏ~!��M�
�R��\�FF��7��pVf�R
T����Ouۍ��|s�'A�ͱ�2�[e)/p��^�c�D�5v�cp�Ï�3�j	�����i�2��aӒ4ĵ��% ���Q��Y�'�D��a�8c�l���hHa�s�{��p8�L��د����;.fS}n�K{��6�6�i>h�s��W�nu,���q�s�>+q�p����J��5C�f��q�»n�ҫ)-�ͽ$���k�lu�#v��`@�g�>�$1QFgQ�0䂤���L�]h}�ܞ���;Gf��e<s>�_��R�L��a^�{� �QL������Q�����r��a�8�*�mi�Gw��}�bR%�A`�ˑz��l�k����]�Kx��u^���q	�ά�IS�ت`c\���^��D#�����_��$�����9OH�SʡUNʕdy�ϻz�����QA�<9���'�.^�OQ]��N#8D�":5>6���{�	'�$6"E[а�VU��0T��s�Z��չk���5�8�!���B�٦�L0G`ث$�q�����_�o�*���]�-�+�I�R�m�/��}ҙ�R��&é_Y�pfi�����>��G�D��Q�@�e^��H��3���㦠�9�|��#v�*�V�!@<���lg����`l(��vx��\opދ�F�:���Ҙs�O�EGf��Ԍm���`J�?:��a=��>+�Q��4.����a*��_鵽��UoK�~5V�d����#�{�i�i�3)5!3D��xJ��>����YIA-e?�B�i����RA!���>۝�Z�hw�g�Jp�Ny6���G���Ԥ���DZ�����Qs1:]ng�M �ngD!��Xf=��N	�:c����eP��Ċ$�/���ҕ%�_)*׫�L_R�`:�(_�ڱ�Z�T��'��ַbs@��ŵʠ�VAGf��9btU2���Z�dhC�0lK�r7ȡ5 ]�I�����X� T��]��$�Q������M|8w9��n�J�@5�X��rfK�Cz2--i�OIeV^���6�[�5���g:_�ҪN�	B�Kh�u�A8��sM�'m4z*��8}��1�,8�4��)&�9Y�h �3Ѣ��|Z-��o$T�I2y�,qD����n��ܡ��M"�7.��qi�ww�'��[���6,q��T`?���w��l2�^��hs���Tj�|<e�0�-�>��ͦ��qz�c�B�t���T��y�l�V���kh|]pF4�Q7�y�Q���B��zybonTG�D�}�AX܌)���x�+z *e��Y}#�x{1�Jj�KS�.�)y{�9���a^ϙxiH��A�YB������R�
l܄x�-b�%h�k��S��c���n}l����ɓ&<�p �i��Q�PG���A�9ۘa�5��}�}�O^r7��x�B��x��w`u�ɑ�b�Z���<]-���Շ�r8EAP������R?���ޚP.�z���R�e4�G�\v�����#�!�ڙk9�z�p���������"�\il$4��uC;�{�Zo'����"�j�>��g��َU~;����F1���A�!5�&�R�G�I2wS��fm���O��.�݄+?q�G�f���u� �S���[�8�9�g���ϝ��"�Dۯ��q�>��N>Ҋ���G�@�d֧�Ќ��x� ��q����n%�b�ulQW:^�&�%{փJP�Fւ��wf����w_�"aKQ��*�@%0og�v]'	��r��E��f���m�i�u��&��O}j���ɿ��Ĭ�X���O��LC`�b:�*�#1T�bXv�Y���8�ݨ���0����l���ml�}��L��u���y��sc�`K��n�,J=?y7�ie��B�'o��,��D����bjpDAI72�����Z�%�m(v0q4��������C����R=f��g߉�����P�J������c#�]i�j�#�� �o�]�t��:(�nT�MFY)���>(����������	��	�cg��/s���M�I, 3�W�,�z��S5۾}!���?1A��]�x2�fox;.�Z���ʻ�A2����&�iqM'ܒ�f��%N��M
d=�.��ݪ�e�ST�H"^�[�ZJ֚梋���EP�=g�ᨃl��j�X�}6���YY�z ݨN%�U��|�?�,\�h8n�J���D'� C^�".ش��ڑ�N.;!!�񸠹��G6}Gj�l߯g7.i:�ZFO����XPR鼷����H��E��d�j���>��18D�����R5!�;��:>��NI���٫�r�T`�~_�),YӲ�4�rJ%S��K�q����n��Ӊm�m�,Ԃ��¨���2�	�[>�L�
B�ѐ �׈ ���B#�I`�C���1���I��c�9����mI����Vx��'�6|r��l��g������s�*:���!�E�ap+%8M�o�(M��%��ĜJRB;��O��-�?( 6=�Ӈ4�J�~���{����璐��&w(]�����z�3���d�	�0Y|���v�eX�W��U��z$�xۦ w�!�oz��;���!0w����P��Gw�՟�'�&Ӧ+�S�̤A\�D��:
� ��Y>����+/���<s7��{"�(�F.���zw�|<eF!��v.�0�d�u������;4	f*�m*�}��_����U-��k�,�g怇ܓD4 (�d�D���|�;������TJ��"P�W�许9����"�ѵ����v�t����"p�)�8���(X8���/��k'��2q��3Η�xo:ƉkVc(��}�8?�I^S�ˈ��Z$��J��r�\[^�{Eކ��O�9�q1�	h�A��/c�}5b�-�� ��*���.�WMy�����s�ˋ�w�^aŪ�-�o�G��D��&3����U�#�1��t8�k[h �Ao�I�����ɬNۊ�OH�'���ke��[��J�,�X�b��bwy���چ���ls��7owX��P��^]�/�(".-��H��x�ax��[�8!�i�����64yo�x/�r���6c4�P�z���:`��� [=�k�
�����*�k;.��T����]�e��0�:G�uUg��𭚛Cv s�i�����o��j����IP��#�p�ј9�#�ڰ$A�Dْ�{�����!��`�H� �� ��`�h�����"�5����Kq7�$��H�#�Í����B��:�D��k�<�C�Z��
*i�>��/�o2���9$X0�-d�vi����L.���5���mh���ʟ�'�вBx:<W"�p�aR���,����'���_�~�4�a���עPL�Yj��*}�?`�����p�c^*(J9��m�1AS������"|�}2�=qd���'p�:D���g�x�@=�@�/�j<�ʬ͊��mBc��.�L?*Hk��B^���Ă����ft*���JYԜ����iɤ�չ�>����9�n(V���Ū9��F���������M%�`~�j�Շ�6rّI��9��`T@i���)�A��>��p�vb��߸b�۫0�`�=g�AT�G�a��4Y1��+��1�ąX(���׷�a)Б����Տ�nf-�|q �}��l>�z|��^xx]d6���	���@v�+ɉW(hx�G�B.����?uyo���<�C1�(bll�C[�>#S:$��]����`p�ϠMI8����ڝ�~aU�\�fZ� x[�/��� �
c(�����Y[���F2��5R����H^���;�p����yڲj��{v�D��&"/9ɨRS,W}5�O�K�w�DV�	Ĭ7�[�n�����T��R���[����*)��~<�`���8��R3�ݼ��^j2��-O���OU�ʐ�n��<���1�Ku����!�����'�a�0�� �"�(@�{7����Y;{{'`�hM�}��Tp�ܬ��+r'�xڤ� ��ki���@��r��>]�eEQ���,�O+�g��W+���K�{�[?�O~� ,���`�}��]U�8�?��S&p$w�ob��s�b���/mh���?G^�x��JS��{*�`��i"���g��A�EDA�kdx��Od��h�� �R1�&�a�µ��0��z�F�~n��?J%�3}} �-�)({V�n� [�����3ɕ�W�P��؉��X��L5�bV�/���i|�w<-X��e���6�8:.`��L����4z$j$Z� �2�E��#o&XR��Pq�g6��:���_\�ӕ���<谭N�̺�O1�[J�bt�?F;ZA-ZO@��$R
m��S��+�vYf��0:x��o{���E,!'4�xa�;(]�(��*�:�?:�b�8���e��hh�&��̦���nܧ@�'Nl7ް�B���k ���������y�܁F }�Y%�_�#���N��k��٪�W�]�r�8S��q��z�z#���4�!��0��Z��m%�K����9A3�d����rk��{���I�$6�v��u�V��3r��q6Ŗ���H`�����A�0��۱��>���Z`z��?YR����N
g�?�#%Sngi_ή���U�x��!	�.TC�Z?�{N<�K'��-����[�(���B���V�9�j��Jx(CDU$���F&b��9y%
H�Ze���B{��f�K�ż,�,��V~ܩt��g�?\��8�Iڽ�AD�6j�����Hx3X��!H_�(&{��4����K���[����r����ŊGA�L���'�m�V:���@e��:��[�툭�t�7JA�R��4)��|�IH�l��&LV��~?_��S�M�u�~�J�5����@��`[�6(�=6��F^5�t��[�5���$5{����G��:�:g���d.�I�^H��5rv%oHl�d
��Ȣ���J�����$H�qR�3}��o �iT��t�x%m_n�UH�nr�'�<DB$�r�e�zPF��Ֆ�Y֜��u�����"�-J���%P����������in`����� TQ�4r�ǥB��l�d��X%*L��M��cv,������){��,(�:����!KX��E���+���#r�i���� !#���i����ʰ�x����vE-���$�S~Y�H����su%��!}��5b�߷=�}	"�D�C.�R\��A-4Zܢ� �n�F��vh?��(J>��&M���qg~��z�j������қ"^E4��H}�zN(j�}�[d���O�������d,�
cc��� ���e��9E5�7<���Ɗ�T�줇/uL�y��%�+p�Tg$���~AM8�dk������J�����G.��u'���,rvL�|��7nL>�����0`�1�L|��4Y�o��c�KP~@��Y�#T�X����Z-��Y�k�q����ATb�^�>˹H1�>��(�����Mq@�=���a|���YlSk��33����)���!ء�����2�֊��c!�K�_�j�@W2Zd������S� �����������R��A%��|�-�yg���Xl�ex6��h?��J�1ek�dC����;j�ʪ-A�Up)I���]��7���Rް׊|��A��1k90"io�28�g�����$9�L5:�$۲�mE�S&S�%t�_�UNiy!��1ntHZ��kb�ߴC�&�a@�[aa�B	��0��茗�mX�v:J"k4n�e��|R)/�i2���m���
��1urJm+^0�d�F	�$�	Fr��t�% �M-NtH;��<�Gܼ~pxK������׀W����ք�x�ZJ�ߣ����߾��4n��w�?�,���Jm�e[���Z��÷�"�@����� 5e!ȡK,�� ��l�X����h�Qu�c��a�R�5�,��{T�S�61�}1�.�eE@ ��I�S�)�獪�)`G"���!F��鈆����\5�\�g�����2�ՆH�T���h3�݋=�k-��]1H�G�L$�̾_�Z�n�JW���7I�//���6o*'5"�>Qf�Y�ӳ�i�U����>�&�{`�D8�'���G�J���z/���W�Zs ĳ��%�����7�#��"�u�����jĦ�ƫ�!;�H�V�l����3�C9��8v��.�Y�x�:���'.�Y��H�Wqd�)v�"��$��U���@�~TFR��jM�]����m�;7	5ϭ�# �s��r$)b�U�_������S��	�t%�~��+���v���^�,��i<R{�͓&GBn�.��z|�B�!�������K�tIyˮ�k��gˆ�J���b��oD�@U�����|)���Y�^'>�����-����E� m���7����YB!����&an�@����r{A�$e��H�SЮd�Kݺ�M������F@H��{2�x�԰��[��nA&�[�ul��I���h�ˁ-KW���n.߀EG��Z�|�Tc߆�Ry���h�%�A=k���2��(:帢��q 1������K/�&�}��ݎl����G����k�mP0�T��[=l:��N����aaێ]���$���Au�f	����6@�m`�̘��qAE���؞�԰0$��>t3@����FJ*y������y��l�Ś���j�u˒V`�ƃ(��i����]� b�r����sw����������� ����OK1H�|<�����ȕ��A��K%h�H����)��6��fsJ
k-D�j�WXYu����UQ�dBٕܷ��*���g6E�ʇ�_��ˣ�RG���󊍦��׋��b��>�8�MW��.ag��L��ޥz�t��
k�����1��cZ��B��1���ț7��Ü�S�U�jp 7&���ҧ?NE_�s���i_O��c��Ǡ�5mm������/_	�C	8��������7"
#%����<LXa��'��L�JL�.�f/�Vx��t��=vaM�&ř�Zً�}�
�<���n��9,]��(+V#a�6��*�0_��.��t RH��c	G	n`��-�@����1�ҪO�(K|�g��/0�?<�4V��m�o5��h�� $�鉰�
՜��:�r�&5im)����>t4�G4�����@g��.n[Y�5��w��ɯ ���!�9û��pH]��wv��Ԥ4\n��C��n^�q0��[/�x:�Qr��n�8���z�iNMS��h7XN�d��.�NyWe���J�N_Eʾ�3��Iu\���*�&�(6�v��Z�jT��(c"�!�ph��7�Nc$5���b:cC��q��:w�*�K�]	��Ň�9[��'O�x�Q"�R�!���އB��c�*t5�D�U^z�+��[�FY*]��D
V,��֮��+H�N�S��Zp��x��x�� ��c{_��+���IN���ԟ�~���� и�$��z�F��~���n0��:9~}�`Dh��k+t�(���ǖ��C��<�t<}�p*�W�EC7 N@��v�+��v���@6�"�X�`�=i��*�_׻l#�r��9��1���"��@XC�)�ձ\T�OH���l�'t������c�SVI�����H�����Zt��&�|�� �E����@��v19y�>a���1�,!�οE#3A�"���C'۶�9�[���i���[�W!����C3��i����M��>m�H���L:��w*8�Xw�e �'J����w��K�Y-�SK7�7���@��g� u<)�tX����� �v8m_^G�'�_΄���&EZy�N*7Sr��;�IyR
w��/��'S�v�Vy;�}��f��G!�E S��֋c��?Uc���Sڏ!�p�4��f��;q��t!��q��<J��o�7=C���b`D^�D�,���5��/�X�ς�J���?j�7���tlb劐�����Pu�j�0�J��qO9o�=��.�N9w&��ü�ᷝ����Θ�y�Q
Wľ����Ө.���!��)��L92����p��kx�^f��B��~��s��ly���F�!��{�O�x�f�ȸ�9�'����\��U���3I��%$Ķx@�U.`,;B�xI2M����?)�<�)�Ʀ��+\����qz�'�!�:����ΉE@Z����b�6�������d��}�v�v�|&?����t5C�ؔ��
70K�j���>8�tW��-}RK�-Ѽn�je��Gt!t���0e^�5}�����'�@�[x;�����B��F���w��uu��� ѮO�;�;���+�wG��2�(6���ݾfoC,Z�e*gc��7��;��/&��a�9�������kw/����Exc�����5C�G굝Cmz�,�������i1I����O�V�xD���t$��2P������jFa�Q��2$�9�v��iib��Ɍ/_�R�����H�������⍮LIy\����a� �~�{�"X��B�]:����L�'��TdW�5^)�M������lY�������>fq��脲;���(��ǜk8S�1=�Х�E�<�Y���F�|Ȇ��+	D&�ᇽ`�E�.Te���~�*�}��x��{`׫�f�P�7�|��� .�h���lV�z�6ե��Z�"���:a}����X��>+�r���h(h�@�2U+���a���T��H�:d3��r�.�rZ�۫����Yc��B���_f �2�ʊ���i^qh���k7��B�L�6�0�i�@7)VG�[�[s�2�܎�C׊�51�4��ض�uA׈V���l_F�L�Κ_�����6�s}��H;-j��1שA%�>"��s��IF�J:O��7��r�����[�}U�`���Z�.��e��0���ؼ�I����	]���{U���89��L!��	�-I�U;�fa�~���o��/C��RK&�sw�Gb��J�����1�|���@HWj MT�!q���f�=�6��Ǖ�j��ny�9
��s��PI�����_�/�c�w�7�Č���B��*��ƪ�w��&BV-!L�}N����)���J��}���c�PE�[����I���	�z���G�>D'fn��;-��m+�0�:���aG`k��� �d��@�J_\�v�+ˉ�B<g�̡݆����JF ��җ��'ʠ�W��L�i#`E��x,چ	=�����fT_k��Bc��6u���;����@��i����d˥T���Qhه��P��{�����t�O��?^� ��C�Lb��B��v(�h�Jv��,�Rt��1���t��4�{-Ŧ*�G�e]��u6�Yi�k�H���Ӻ�N�y���%�1~�/�l+��mbdj�%��	�9"�y�i 2bRXgۮ�SކN5К�6�)M�d_W�m�#��/������C���)�9k�l�N�q%1]��`,��/�5
�cGb�#^R��R&�_��@��}w����I�`�n�:���� i5Nk��X���β�=(��q*�άG+pX�J�x�Y����VLA���"؜F�O�c�HL���78�0Q����1r:w�w���P1'��|���]�)6Y,��?*���0�	C��g��bǄ���R�?57y��a>z�3�@Q��#���ko�s ������ N^I����q�A�X ԩ����&� }�0:&"A��|��Ǝh9��m��(����
\�����MXfk'��v�9��<�r,��1�!���Ea:�[���;�,����K�pћ���<��%$@N�{�W�3�U�Ą5�6l���p��]��"WS��
j9eC�fI�v4z��/�/�i�obr��g��'x�{��� �#�sI�-��V�?�*�P�BԂX������?��"� Pn4l����R�0�T�x��
^��+�B���o퍃�+_�^
�y d�x
2� UI|��#����qƁ�⽌� .`d Wk�T�h�§$cb�F��#��t�1��auX�	�7�8�`��V@�?�H)�U���X���jt���O��W7�7���#�0�\�y�k�x=�Q�\@�i�V��o����&s��QY1�6��/�/Y<�pDe�p�}*jm����-'G,D���p���7�<����9!--MHa��F)?1���f����Z��z���< 4��BF9�r+d�	��$&/I�vm�]�!✝é�C�Q��ͧ�'���۶M\�+k����o�C�6�V�{̰t�I剪����� ��??]ڰ��\���^7�*:��Q�QYQ��/�=ɂ����> Q��{�kh�E\�e�ו��C�E���x�>����3��N{*���N$^H`�g�W*%a�2�D"���ۺ�<��XW�	0QlU�cVu���]�w(�y�('��@����)���2�/��or���T�8Z��������u�E[�ZP�q��<!�ܸ@&��)!��q���|SW�@D6��k��f��n�!׎f_��F}���8F���;h�̸KN�*�B�#�����=�y�re��RtՃ]>$xa�0P���k����9"I9��)�9��Ϧh)To�ď�i�\�T���ʸN@?:,�M������8�,z��[���R�S�%�M�yM�����!] *u������يmg���*��<�9�~�?�)�t���k��֣{d��������w�6��7�8�/����t�:����'�2�=���sթ�T�O�� ����!��2��J�T����g��2͏��@��Ul�1�,���R;�E��W��րN�ZJpo�W�z���� ��RK��M���E뇷��4���gd���uYۂ)��v}5/�;�^a�m�9� n��E�=�g��~��������b$�7"��m+ˤ=BF�����cLՒ�C�
���|w)�̼��f��@w�E�Y��oZ�o�-QV���g�ݿ�o{���i����my���j캒�k�"�P
�aqp��Ğqm��5 ��&n�Z?��=N��ږ��^��\�O����Y��&r�EKU�ӭ�q� ����@
�8�
������fQ����&P���\ͥ�vq<%��Ɔ��fb��d/�NPy%'V�~����	~1�(�hN,VsH�Z�l������j�п)|���N�̿	�r����a�FC1��Ï`�4��s���KKj�S�^N��]=����W�5k�ʑ_�V�n�5�V�����4c}��\53Vۖ��f�loa:V�W��
E1����Due�n����C�[5M�&�j��YZ|�hg&X��2�$�	�(��m��\�	n��|�(�%� *Y��V+�/S��yٕ��� [�@*���4�@c�I�p�E��M�"�����!$��<H�"�/h�O�U��w�m�0��;b)ZF����m��M ���9���\��o$����C��ܚ �����b��6��]�����an��|�'���!��6�9���GT�F�0��B�X�{Q%�
<L��[�@����ʸ%@� �4������P@���Ћ_^�I�ʜ.��BJ�HK�9��bq��R��Y�\��O� �Z��i_���W���Ҭ�{`C�p�5J��1�f��ϚV�[�>Í���
���9a^�}=��w���d��{�ae�-1k�Rx*��]bɎ�-�hL�{�����]�h*h�1-J�]��\y�Ĭ�X}��H�~�7�d+Bw��ƪ�6�3������q$s��"O3 ��T&^�f��L�Z�����>�Qjp�������>3�M#y���d)��d
�9�-���S�f�v{���f���'����LIH�l��'����=���\�V�>n�����Iջ��On�p�A�BҞ�x�y����u�`�*x�!ˌ3�8��߈!N��9�W�>��nWo�f=�IB�{��FL*��2溩�pg��8�Rh�&�U�js��ڮj9��&I�\ؚ�=��ju6����78W�� � �+�*)�K6�S��j�a��t�xGTb�Z���~�lΎ�3�5M�>3��zGD�C��7p�ngiP:�k������9�b�Mv���~�FD�u]�����
�܌._�J�`�Р_:�&�}K��;�7o0���GY=��C�?c��ϡ��`WbrH�6�En��5Wڢ���%���=�畀���?��1OWk�8�\�=���M��"\p0�6_��kvO-��U�*A��A��r���N�˼��Ҳ ���]�RĈ����M�.�E�'��/���):��4Sjy��dU|q�[S� ��08#�ED���L��J�7SL2���?�Щ]�vs�����%W�垤{�8�A@��Z)+(ɦ[U�C?��V� sRB�� Kf����G=��g��������u+!������a�E���K�y�����\e ���\[xG�#�Q�}ϯ/�U{�"���[�L�<�W�G��+�&%�ؐ�D�ˢ�bړt��j��wD���X<�'���z߁�_ՔN����H�5��F%l�r̝����`���%��8�?uJR8
0uNO�)C����@/��i�"�C�I���L�Ҙ��;p\{>�+}�w?E�I�����\�����CXk�}�{�G�vF^]�;�r�������-D	��q��cH�p����WH��"�F���n�
E�уo�M*�*ˏ<��m������;x�"exuFe�uq���+ep�R�5�]�v6Z���q�x�Ճ9���p3��M�៦�F�)J������'�	�''��P
U��ħ���	������kf�zDza����(�������f>,�1n�/FE��Y7�)$��c�^����H����(�w�O�T�{�.�y/�椘n4�pw繊D�G�<��߿x�ޛ힕�r��hH��Yn��:��*Q���E?WhoϞ/���@e�AK�3�4 zO��紃1��2-����Mڌ�ڰ~�G��)'�z���6�:�ݤ����V*��1���D�+fH � #��X��� ��t&p��h��blg���y,�>�c�����`����-����������I_�B�ڞ�vfm�鰨�7�}~�K����P����@����u)D �ҽz�8��A�J���X{b7O�r	����+��mP-���v�O�0��~���9��Ios��'G�P�t����5)B\5��騡�r�Zo���8�����p�!�v�fc���L("�|	�����83W���� ����%{�m2�8A�����B���ΰ�=��'����[4����m�}�'D6���+Z
�Tl��K�� ��M�Q@Părd�N��!`�(�����?�Μ� j0��!�O�Q�+5�-vn�o��W�Cze�Z�|4��3Ƶ��� ��X`�,b���	F��kG>"^�4cܴ��X�E&�w�(/�>ٝ&E���#�e���M�ǍQ��eB���l�P�0��E�P���ͅ��N�ڄ*�#�M�^ẳ̤�iz) ��7�Մ^�$�F4��t6���u%`�+�	�m����(љW3�Y���ՠ��?���ݞ����C<��n��!A>���;J�i��^�r��Ym��8���=��M<l��\B��do��On�����m��±6ae�bL0���c�\f@�r7nI���N��htV����Q�B�#r��U��~���U~GG��֢�!�Ų��=#��ow����K�1P7Q�����Hn���쓹ְ3����q�PҨ���Iv�'an�{1�5����u�[�'�7�t�1d�<L�_�,4� �,�O��K.I��oŵ��F��:7t�DvT
��8�jj+��,�C2�n�4����]�Vyk�GH�8ξ�����-�C���84�~Y�e%5�Vvs��nZmB.�FV��oL��6�&-����p�Y��[C��"Z
i*�V�i����7�\��B���X�isk��h��<�IJ@�D9�x��`�$M�Z�-��eQ#���܊+���$�q�$���o�l�w�*�����p��t���F_��Q��?�Z��چb�{���)5�)|��$o���\�(�9,?YM{İ�G�l��V!��͏/48����q��d�����_|��(�H�$��,��ŝ{���jD)(N;XT᫧��k����~�`A���8R�RU��z؞�M�u2�v�~�Įq̘��_92�V��~�a�C�53�u���R�'����_.��<?�y?s&U�>߾� (/��ǘ{�ɲ3�Q��(�N�^�'\�G�8F�܆_.T�\D�:�.��8��Q��\��
8�΀��2{g�h�i&-��]m�.�����:�s��!Ob �|Q�N�5㬹t���K�^�¸Rd��ݏ�y�<y`&�v��O�X�~V0�Bñ����{3�>Մ�ֽ]$��{L���*�Cv�"*@��E�aw;IpҺ����g�~��iog������#�|m�a�T����a�{_�)�����U����w��'H]�q=fO����ы�� ͢��M����zw	F��t���}�%��{�g��=�8���7%������nT�wGz��Ό ��E���I_�A�����	��4�6�a�_��4MLo������Ԣ.f۶�i��+?��Ŵ���m�?D��&U��Nd`}}7��W����:�d�;7(.�>Jq>�\����SJ�4d�|m.���@�yi�����U��B���U�(g�6��O��4v�;"(8k��]�e���!��{��pppE�+odC"^�\�J'q�T��Q��O��Ɂ	5v�Zh�ڕ�uzAm	�#�aJzU�.xg2� ��7T�8M�&ES�/Q�Tf3��j���QwR㌲A�1;g{R��i<=�@���b�*�Ux&�G���V�K�&_�l���-1uN,p��φ�x�t�Q�MB�^t��m�X���Y�ݠ_%DM�0��l*�e4�ԥ���ȥuΰ�ل�v&�J�@��&u�:d�L�T��,s�`.E˲�5��ꐮ��
��Mq}'U`"2T�/���KP�2�x���su�H�6�����t{��R)�S�t͠��̵��N��ߧ��gǕYHzú�_#"��]�2�ӚvL��{�K��P��`��V���<�gmL�gOսw,�) ,�v��.��5���WN��=B��pivn��U6 "�N����5܆:�}�r+���o�Sb�j�z�ys���Q�ڡ�5DE��+6�����:��J���+p���T�����%~G�'���b�����q�f�>a���(Sp)�X���ځeS1�Af���{��,З���^|�ۙA;9�"�3S�����~�Q�T�1B��'^��:>"�4u _/Ǎ"B��*�ܦ`����a�{�I��x�x���4��l��{��6-z�;��K�͂^cc�3�v�߂������T�ӿF��:B���	G.X�/�r�����ޢ��5*<^>��LԺx�Șx5��P�:|�['.������M���.�3 ������{z=��䮟�}����Cls���Ș�.��@(��o=��M=��^�����Ќ��?G���GcLx/������C��9��f4�Ę�=@J�6d�W
ʥ��O�Kq]>�A�y����.���pT��rF7�j����`rv7f��{�_4iM��[��^����PHzW`J�I�q���)��Q��T�a�Y$� ��H1�˲��cbA�?��ۏ �%��JA(�V5v����
�,��IN>z�𲝽T��rJ�%#&�6$��D7u�;~8��5�P���RN<�����R&�\����S.yW�<^Aڮ󥾢��%�ĥ�_��nk���l�]�������p\��!M�
�c�}�����S5+�rn�Fhe��� (���f���7� ����.
�_~u�K�[��I�����X��W[������XŰ���aB�����j�Y*��ɉ�M�un��ì9���Q��'=r��ш�C3������%��/TT�>:�'Vkǭ6e��jNP�)�8l��>t��mء�H�WQ����-_hKVa3���zp�����
J
7�Z/y8�ܳG���]�%�x��XLTV�h�+W�	�3��4��ovu;���_/;!b�t��(S�X�`������V�p� ����'s�I�ޖ�l��������	��0�;=���R��<��oɱ�M���{�S�F��&�uY��YcH���� �\@%K�7��b��L�а��[�}� ��S��/ķ�Ġ�c�2["��Z%YvQ7�n�k�+��Z�U��A�1�	��؎��Rh]]Z#
������6���Y�%0��ʏ�+.�Z���8T�p.�J�Fp��xL#��B!��2�q�i@摲��u���KE8(}Ij@�:����g�@B�O��欪E�XQ7�/�3g�Rǔ4l���f�� )�6V~2N�ᇌ8���o�#�}�Lam����!Ll�j)��6�C�Wb�o��u꺮��I���j;o���F��ݙ��-yg���l�ͦWt��C�Ĩ��h��3w���	k�N�*<8�'Q1����>ߠW�W�� BG���:n�t�[Cb�udD�K��R���&�g�X@�x�t�W�������-�OX�Q��#���$g���>OZ�/ѹ�Fm��I�e��'�/о��	�D��P7ӴǼ���	GțeȒ�#y���k������"�i��vH��\؋�G�C�I�1z�9�L�����+����!�>HB�h0k�;0R�}��Ν~���/#H��A�Q��"�^�T�M�B
�d8�� ��Kv�4���<���(�T����us����g}�$���p���DT���w���{6\J�$�����9�����_JcD=��`�rیe8�e�
�j�-tL����N�B:z\Fc$�c���dy�o�he�҉�5K����qNt'F9�ʢ�ia��&p�M���e�X�*{�o��.-Q�3�V���� �]����������d�����wv�te�!�0�J�e�a�m��ҥe�P� ٻ�3�ON@ѹq��ݳ���qֵs�5�'�*�gD v�/m��+��,c,�r������ƻ9��1�6�ߨK8����7�!��2�T�#g-�'��1��VeM�zZ4��;M@�����|-�uc�B2��E
����*��O����au9.��"&�n���x[�N��Ԓv�~�3ƣ���VB��i!�=8t�M�z�5�NkK^�.M��8��<äl&��Y^'� �/��tv�	ʑ���N����@�] Y�,�Z?��a態�����:�d��B45�:�x�/^@������ؾ�1�x�||�W6�S�`�k��I*/C�]���\��&�J��f,���~7�"ױ���j���z��Ғ �i_���'k�vα�d'8`ߌ��
0j��IG��H�����+�e����l2ᖥ�M�,�v�n$��Q�|�4����"b���b���Nv5�KU�]و�Fhw�V��f�
q�.p;���RPg)F�m�'�f�q�K�B�}�c�hr��b����AJ��������4z�?��oY�uvn���@�����?�rW�j_����'�{C�����D1r�8�f �0�]�+˩,�K����-O��r��qVLup<QS�Cld��d@�����B�u?�J.#�7�d�zLO�<���pp� �Z̐u���!u��Ꭿ#6��3���^5݋�"[�0֝�i��\�(8Ԥ�v�m�}0U��M�`.�>Y�/�T�Rj6��{�@)z2�=�oDB�'i�q&d^Jp�����:20�7�A��P�dR������X6�c�<%�j��ӀP�⚺֚N9���W`�7D~��m{���c<[�S46/]�J��jE5���z��i���4��@	Ʃ��˾����t��T
6��C��k��v�/h�&$�:�`��O����>%�j@���5���i�ޏe��J��7���P|ŀ�KT�mm*+����4���eN�pً�X9Y�uLL�h���Ӣ���Upk?����P޹Eh�/Ma��Ζ�I�]D���T��5d~g�Ʒ���G���>�r����H�y�k-��-]`��}�N��I�9��R���Ձ�S��#����ݢ�!Y~��s\0���Į�3��8
�0�s�ף�r���У2@�Ų�U�S����(��m�8�C�����ZGʇ���0)�O����n)-�V��a���(~F ��7�-���q�-7��뎟߽��θ��%��]�W��
�P3� ��l�o�V)5������}��J=f<�F�����C�1���U4L�X\D��rk+��
`E�tWP�}�[;yXꏶT�-�:*�#Kf�|v��T�M%ML}����N��	�X䯟�a�"�)�b�Q�	$���mL�g�̘��N�Դ�N��~�h�B{SZ'���
���.����
��}G˚P��ezPہ�6����`�m]���7#�'a~��l���h]�$�"q��7�j��l�[&�]���>����	�
��4sc�x>)�@ġ��fQ�M�+\
�1�[���/����2���j�EC��o�к�T��%�v��FBl���R����TWص���S��=JX�-F�R#��6[��r�ܵ	��E�i�m�A�]�F�H�`4�����&0���Xg�q��}��֝o�BQי^�^��w(��dx�2�!yZu�W��h�;��X�Z\�n���]��W8k`ڊ�FFv{���ԂG/,Aۮ�X������Ǜ�� ��ڊ��}7�b/5�Q�7�3�ݓe�lK���
T��#0�w+���Muã�a����ܤfCǱض��C���T9��R�p�fFeE�i�\j�#�߾���|��u����X�!�R��z����C����� ������Nܮ�k�!��!&��i��#��*'�W��i~����̇â8
�p�
�ؤ���J��X�GI}��M��
�)��~4�B`*U��e�1�l�,Y��-��s#%`d�D���t�]_'um1�QB������q�LR�<���:�	:m�+4�+���^��.%"��osdA~d(��R��3<`�ٟ� ��Cj+�U�}��E�W��OE}} V'Dz�4 �z�
�D��_B��}�*�s�oO�����`IT$���NY�k��e���dV�Z��쳦��&���J�L�e��J�YX%���>�E�C: L�w,g��j�B�-��c_�BM�U�`�a����d��s@�!!7D���=2�Xc#��~b�(�v��� ���@��o���ԣ��	��߿)��������q��DT�,��-�G�C%��*講��)�^O�6�.p��	�����%��_t�@��s��f7�
��qd��#���#���x&^��;S;C1v���]cv2�⇠�IQ�r�RCq)�j)4�$�����g̩7����=y�]W�����<����%� �F�q5��Sy"u�����Zc[�NeSxJ������"�7��V|�No@�j�j��b�n9d%��X������"趭���&�;���D��ә2~?���=��0�����!MyJӼm.�2������BF��l�@��ht�1�����'o9y��Z�[8J��`��0c �^�?�O
�l�Y7'�k��V�3���C���f��0k�A�h�7�=4�D�L�?ָ�ɫ��x�]G�RI9`gkt��³-ğ�3N���/�<$�\8Ѽ.��;5���eC���3G��ul� l��Oq��}��
Y�D����RM�OQ�]�"	uS����)|��+��P2�Q��YV�}��ԝ<"wo8,��G��[��Q�iL������/B$Yx"O����qa�6��[�zQQDڜF8n��X:��Y^Ԕ�Y�n8�l���P"��1�N��z��C�k�eP6`�c	j�Y(�R�{,Q�����C��z	X�o�?0�����O|0-�&m8ꟚYo)od�����s������E�yqp�\��a�8����f4�ƿ^�_�}���#�@U���^���3�`�Y �&�ؾV�O��]8S�־�}՞�i�E��Q�e�_8�؋�~��'���)�M�$/qRY&�+\��C3	Մ�E�"��|�gH0��Ē�`����&v��\���w�4OHK�u�0*�V��d���ۢ�j�f�]y{���.���l��W�N�^IG�G�����������6�z$�h����@���ӹ���y�$�aݜ�q(����ν���^�a&4_���rf���D��98�8�s}B[	��|=���_���@���?=�^`����٪?:Be�&P|L�%�v' �Q�Y�<�ⴶ�����'.��eSk���>���Vv�e�T^�S�� �N���|ӍXNY�n�lG�X�2]-a���l��π��_�[<������7雛>��E��"G H*Ie'9�RU�qE#-�ԷNJ ��G�C��H²J(+�G�׀��y��ŶZ�P �|ɥ�cS\4)f��N�76#�	 ;��y�� [��e�1Φ��Ws��v}����vQy����j;���^��LT"ME ��q�zV�7�� �S#ʓ=Q~{ꫲ3����
c5��,*V`p
;�k�O>/:���ILRmX�H R��Mj;�q�,A-*iU�myq�aw����Sn���[}�� ��d�m@�K`a�N\�f��I
��A>���ɺ���)�4w]�KY�!�v����������%*�)9�p�b\}l.RE�T�.'��ɳ�9V�v�7�3�UCǊ�tfC�$��H���XA� ӣ�n�����6��}U�s���3������V'Z��.�PO3R�Ǹ������tMk�Un�|�$`�՝S��?�п�02��>�yg9=r|"v�`�"'�P���,=5�;U���Xg��9���6�e�F�L�/p�^�EK��zc�˞ｚ�?v�.���U�Q���w�!��Ŭ1{�.$\w+�>h��G�|�	X�ᆭ�A�z��C ����O��(3Y
HG½���ݠ:�'jn��;}�*�%��:�ߗ��2.�ϐ��cJwʞ�Tћ���#�Tz҉� y�U��a[��H�B,gBY�}L�`�+�k�*��`.Ldl�H�JTe+�Ҧ��f~�����?ɹY������V����7�0A�J�� �5�%q�a�{"g�?����X�����P��.�3���[���极��z��\�B2��[�J`��8�}L�@N(@�܃����\��)*��δhJk�U}�L�_4u�y9��QE��]�����Q�´]�T_^e�cJZ�ń7� �k���B��}�R�6c������}@���o��^���be��o]5��}���Q�i�<�*F��<��&Je_glC
�!�����pϸj�����S�J�$t�,�Jb�|�$��Z�C8�6��^/��vx��Js��8ғ*N��S���TM�';j>��9%X#?6�`Bku�չ� �k�o6w3���%��{��jRH־y�#�"��7�	�Jѻ6�KO��3+z�ԗڷ���b�5��R3�.�=��gW�@1-�kh�>^���z��^���) �FX	~���!a_�6�����y�Q�~�D�WA"�I����y��_?�� M���+�M��\;-6��������H:��oP�d�������àJ�G~�a[au+S��(�L�fg#�;+}�Y�]a�\��ѐ`w��7>�����A��5�n'�x�����O�)�@��d�z�g�$�!��k�z*r�rVIc��Ț�)�)d�h{�\���,�!��L�О?�86��ad]� ��yۉ�dw$2�<�D���-���Q�����d���m�%��̛)��TF�](��u�Qe���?�ZM]���T�54g����i��)F�����d %'�M`�l�cG�_���&��Y��X�'�78�'OEa��vJ<�Bڿ�f�������ㅼ�����+zR2n�ȱ��`�T�ँ��v���D��c�R�]g�HKC-�d���V��7�xDT�6k�}AU5\u"�H9����G�H����e�1y�b�]���j�7�(��ݴ���Ȩ�Q��-L ��}_C����Yi_�C�;E#
�1���/V�� b�����kp�㔗���j#_]�	7$�~TY�tD��6U㏨��P��t�#���ָ�7s�������$&w��&��r��M��*Fgcj��z���`�l�šd����󍳸\����b���
��zz���w�w=�H`%ҭvj���n����)S�C0������:,�����T0 &,�W~�%7�8X�^����Z����_-$?;��"j6[���*ǂ�7�C��b-��g(u+6�>E
��dzd��{��I��X�
�g���b��1Ҋ��^)c����[W__Y��mS	_ *�v8,~C��/ط�'� ��77�)�m����+V�D�2�dƯ$#_�D4Qդf'o�'t'��Ԣ��q{"�E��W �R�p6�d�01���X��
��xn�,Yg�Թ97�y�4�r��ͨq�N��<J7������]�u�řY��wEPԜͤ���W拿���d�G0�OX�����.I��᫷	�l(W,G�oU�D�$  =:	B&& �kj��m�@7 j77�#"�(���Ӛ��ؿ஺�#���5�������*��t������g /Ɨ<Li�j���z�����ި�^(�{ލ8�PB�~��{PG�
[�q�G�?]!=�^�r`k`��0f��-�?����P�@��r�����q�ԅ9��/�*"Ө%����z�*`��ȉ��u/eB9㟍7������ۅy��\�q���ֿ�8(`E1��}F5������>&[�΄��G:�OM��\	{���Fu����}1YC,�� u���J���X��xt+���{�{,δr�g�}����
X�K���7���KT�_v%au���l��;aD���z��,�b���Wb��o�>�d�OU�@�6��Q�����K6s��ɱ9�S��=R���� ���߄��->)2&�+��9�X�qH�tKq̛/C�����Pܗ�|zU,�u7�xԄ�D�U2&#�uxTMUCNC8���f͑��E�U�sy锼�c�ω o<e�7�X�I��P�d+���׬�����@��䁺�ψ`_�ƘEVj;��f3����9�צ�.=`1|�ȅLe�U��aIN%�$n�=�v9[za=�e('���-B祙1_��F��ϣ������I��{r�N`B�p���������^�����e]
�C�봱'����f������ja��[��z��\��l��T
�ʀ�j�A�x_��E>�Ě:<���&���T�ϯ��~κ{4�I�F�B���	��.$�����?.|<А�Ya�O0T���Y�GZ�Mtߔ˯?9��-_!�33�Ŋ�o��II���ޒ�����}�[�^/���ŏ�`�;3�[�D��T1�f�mq���~�ODC�1IY	�&��*,���?b�9����,GN�W�z~v��bS�2�i�oK��eU3pk�{x
�F9���Q�`P9���}�M���wf����K���16�t ړ�����MС�w�E�
5������v��2Wl�o��5�G���M\|��n!u=��tF��C8��y��̚��G
��>����'|\h Sn2��Q����RYdx�GS�� q9I���ɚ��m68�ާ?c��B���ԖԞ�PI@�ߝ#��D��V>�ݸ�0�!P*��+d��W��]b���k�x��VW����'����ԉo�P����wں��?�mn�H�W�P����ވ_�]�b�{���႑+����Jq�I�g�����I�BƘ[J�IFf��I5
�OΗ���V�S�y�u*⥝�X�E������Յ,����a_���u��.�����d�S�!
K�cYR,�`(zm�+J��[dXU\m�K�R�XsQl0�G�"��\�g�F�>���K�<���H����t0�����I6���b�c�6$�d-�B��o���;��8,Vxp\4IHVԾ�� �u@�p�R���%���#=UAK��!��s��GF=��v�:��-����ٿ��KZ�	�^��p<"Js�X���_���ě'?�Jg���6 c��a-���Q�$�V��rc@4���r��!ɘ�%�����x�E���
E��^ճ�p�G-}n}�TAj���fa���n�2�Y����M�5���*���X9�-��aMS�#kfF�c=�Fgh�>������'��G8F/��X��I�˭9נ�l�L��Ķk,A��{�[9�9P��Z��J������3�A�KB��ndš��Z�$�_�j�3����J�ʚ�ַC>%��' 1@���ظAD�F�,����F�h/� �a��D��KqB�8���}qv�%�0w!We _�3x	
��Tb8�i�op�u��'�^5�	C�u²q��B�����'X��/k���۠�����������ަ� 'T��;����M��
|�V�Q��^��vƦ�B�V���wh���őN�I��4�p��@��D� �����$eaG+�>'-p��bk?$S��.�1�ݒː^u��ت���oS��&˯����ɗ�h������P�ُ�5t�!�S���7�l~������*�0&�C�5G��$�ǝ�OЊ�i�O�Eנ��8��o�Y����s����q%�����Nd�s�Mڽ��A|�p.�t�}>��ڠ�4��'�Wq+ $�P�G�^�t�ƭ���)���~���O�T9�y-����,�WP��d:�y��	yQBK�E��6�mP��g9
�E�_D���#As	��'�<r'��%�$-�̧9MR�rt���cBV-si��N>!;㫢���cb��չ��yQ|M���򯭿�@�z�xi�������1ƃ߿�d�j���QҸ�4n��~r��\,c���;���>��%��- ���2|�Fe*�T�o�I�v�hTݙD�n�_�J�*�F�f�"}%�,��PXᏇ1��n�}�_I^�v�8���n�wd�2ɭm�o��42�i��
f����0���B��$�ޒc_�OҲ[�&�L�a�Iߨ�6�+GP���}�ř�I��� 	��qq䏙Fj�L��j��P&#���`
O����O���:
욡��w:+��TV����Ic��5�Nn^�ZF+��(�����Ѷ��D$���v�[����j*�P�^���h�	�u`��^1�3:OW?�0�y+�0C���T��ֵ����v.h����d4�O>� �z9�˕���P���5t�,��Z-�۶O�<-����R��FM���u�F�Y~E�l��w��iG�,�7xJc�����`	���O�xy��.1<�ls�m��b�m)��F�|�~�L	@����ԷΗ��n��Cw��R%���
�*` -�pq$ݵ��?Hښ,Jf���j�$�Yo���0��2��U�SX}�݈f�R�Bo������(C%Ny����m���]��	L������W�@�h3�=>��>�>�'r��|T��%P��hp�-�C!��t�e�Ƅ�5 ��QG��]�24넻2���k���AN])��yK436R�E`M%�V�qº�|�ϙĦ�Ú<�����{�g� �� �~׆>���J�V�����uL�&���[����Ib�j�jǛ�Igx���ԫ�©�оt��iM�����\�m�чu3:���$��Y']�K��粠��,��ᛁ�z���X��̉ ���sUe�7�H���c.N���!��I�yC��u�~�Zx��z��l�SBV3W�㉳iZ�yr �]%�����:#��?���4�3Zw�����G���y�GW����?dSJ;iL�Ȉ����,���S��V��&Hִ�:�k9��q(Ro�hī��{��50�8_n����y~gU�}�A��[,f�V 7P*� �7������1�j��㐙�J_�r����J���i.��p�0�����~{j{�y�������.��ϪO={� 3��U���-��V���\G�� ��v��"I/h*���~�ION��u�zr�+0ԗ�H���:�	��Ϗa3S��3�/�q$��Ą�O�=���pdeTcɰ�S'�8̑n�z6�/u�=�3��9���ك���k+������P�M�ڀ���K�&[��+��MY�GM�=�{��T��3ku~�aA�5Z�ϼ���&��I�J�L%�׸��#�x�=��g�v��]5ɮg�_�p�7>�'c��m=������2��Q{�[
�H!�̤��d���h�Y9�m��
g�|b���/	u�ɣ�����v����)���*�n��Wfe����7:�ڥ2�M=�CˀY�`
�逘��t�gb��ծ�
x�[&_�o�_:��a��6�瘆ZZ[�E�����]AJEG�٫y�U�,�y����ŉ�!�=�fx���z�y�؊�&+��v�z&=����#��K�H��[k��+�nwR��)���4�-h���^�)��,��E{}��k�M:mMU8t�7�)�CB~{��{p
i{� �%�,T��Z����*uWل��A*s&�t{T-�˒m�֥�N��W�G� �H�s2NSZ��aH@l$�4���_e�����2���u.�xaBL<z�hy�+/��0�,�+׋~�<�yHA��O
�H��x	K_�a|��#���a�E�\G��L&�ǋ���+י�����U�'��'r�ԮH$��x��{�9_i�������G�����q�4g���,f��f`��4n`�n�}w�0h!�oWE����M��[��=^�I��yp'N���=��3�	�􎾝�Xp�q��|wҗ���)p�6�%����fd�Yh���4��OD����T��l7�AS�0�^�\�@�6��T���΋ef��F2�]�	��R:Ґ��'���kQ,8J��X֚�L ������Sk�0k��+Z��y0Jjx�}�k��=�ϤZ�B���H�.}�w���x(Q�(�F��~mܹ/�G:Wc��Fز]3Y�[�:�t�V�.�/4}��٨��B\�B�(RJ��@h��/xc��$�
�&m���n�y�E@%R�<[h�=a���.(_�Ba�:�xO�c�X|1?m`h�� 2���.�f=ϧcݳ#�%qc�=�)����߫�$9z��4�zR�sƔD����i�����^p�r� ׼��0�/<@Ė�]\*�k,����$�A�B+A���p�����2ٱX�u7�;�A�x�ђ�s�'��EnWn-��b& ^6�y�\�� ��"����d#c��o�f�2�w,���չmR����»�3�9���4ck�Ь��hԽA!1`j�<�c	����JM�潆5T��!�"��HX�{������������#�ϼV|�m�S�7P/)����
Щ��?Ň�L�R�����9��R<�K���x��Yi۰%m#R�z�q+Ks'�^D���	��]��Wz�dߟ����\�Zr��� ���`��ż�#&b�ꯥ�m�%��˷3�~-�(F<��u��t�r��`w�/	4��~Y�{��*ِ[d�yI���jl�3�!��5U���+r�h�GЛ�{��q�,���i^��B��b��6���l/y�8�ģ�E��-tT1���V��T	�B�B�BJ�� �N}1�9&�Iw\`q���$�n+BKhc��&�m���9�'GX�������@_>0W����~E�uIcL��FJ\"w������� 4n;�~��1f��}��7/��K\^��<re�[��|��$��+�* ���Wl�����?0{)u��<r-��`���ݘѢ��d���g���p�V���#� �P_�#kn�����BD�;�F�\����d1�/|s�<�Ha9dfeU�ʩ�x������5�X�ޥl�>đ z4Q�O��	��,@յPK�u;E��H�Se�[u��	Ֆ�ӝt�� e;�6��k����a��NpV�����':��*��g
���\tH�TT��TT{�R�;�x�m�3;D�
X�8ɕ��H{!�gF0�GMpbL�ͥd�60�ij3��<S2&έ��۴9�F%u�s�08��[ �$�A�~���\��q��b��Ѓ:�I7�t�g:��ٻ�(����Om�@�=�����!lz&�\�oHT?�?���e�W����lF߾�3k�|�H^\#�}�h����9����Wُ$��V��N��k��O��r�3�-?��nf�n�e%|��Ͻ�8mk3�{d's(����`gzѣ�ѵBY�o����N���M�ٺ�$%�ip<(���#'�]V�@N����*����#D���ɑ.<!r�ȁ,ė	acR�* 4 ��N\��
��$���ݨc�M�\�P����i�j�+vI�̋R���	�4���>۫cT�Ah?2�6�&!]
�������J��E���"ҷC�N��ަ�/��v��F��՝�2ɩ�2��K��H��Qi�[I����xF���Y'�c�N�A����w�ډ��:��t7��f�4?�c�t˅S3��g�A��I��7�<����p9����7�d�{Zܛ{�&�'tԧ��E�/�V�'�Ă��5�N�ZG{P� +�?��f�H>�ٚCG�K�ĕ5��#NkU�7d&����k$:5v�^r,4p�}�e����Rk���]�_�,~�U�\}��РO�p�;��"�*�0�L���i,a%��Uڸ �yb�vAc�#H����
kd:���� (֩�
�a9���k8� $���ݐ�0&�0�6x?��/�H�E*A�i��$���gG�LMDC��;:���f
\���%7��KrR3�Zc�1��H�@j{KѴۀ%٥Z<�$�,/R�D6q�P��(=�A��A���S1bp]W��,i�1�)��x����J<�V11���cbh�A�s[<�o�愆v��VDٮ�R$�d�f��#n=G����aJ��Fř�zӌ|��b6-�@%�v__?��EUv���|R=`A�7HFy��o���/��Ca�9���K���6�����T�l�pU'���{](Ż��q��_��=Z�{���_�-�l��� �Jg��d���N��Q��Ԅ2�pIນO0��x	���%��\thYٳ����Э�vjy�U�e���jƱ���$
�X� ^P�x����Uo��ם��bo=��tz~�o�]���������O��U�wD�3bh�ì���;ZX�b�b]F(�R���#���g�HxQ�ݘ���z�+�Z!���DH�Ϸ꣬��q��i��m��C.v��4�$X�sY��w`mW�$@7��dB�Z.
�w5H���|�1Ɯ�Wpђ$�-9F[H�F���of:�Ы�{�6@���[�*���Xm�aW P���rs�����iZۑ4��-�_(�p�>�@~qU�rt�����.�(��C��i�İ����\���&�J{#��tyq�j�c�O�Z<��A=��F����W6���Q[���~��߈|���||O0Ͻ��I��P��<1�)[��_��A�Бm����=q*%�`8yb�H����yx���hSCʦS8*�x�}߁�%�*]:�$t�˲F���
��Vu~�j�`#���;�q� ,������:V84�Z�҈�������r��d�0h�ݪR�vI�@VyR1�(ʎC |5ϲ�$νbl.�U���5n��ݱ�*�n-`OJ�� ��.���(ڤ`Ļv�ƚ�c!�?�%.,�#��^q$	4*H����XR��*�ό��	�;�wޠW�C�N�w����`�Y@�j�{.�O�[��2���IO�����1����������!YxCoVOV�-&X���5&ρ���iwO��;ď*Gλ:\�N���G��w�z���I�7x��K��p;�?K��ۓ�l�X UN;��R|U]$�׫G����g\\_~Qf���l�꼚�nv�j!?k�5��-A�J�o�7/=k���0����nJ�`�G^3�8��Rȥ�?;�=�$4@��;x���c�\����� ���M˻�`�M����ȥSʵ ���+[K(�s��j�%фy�3��~h�d1!,�R�~b�M�Yn�&'�������*K�r|�Nw�j��J��6�ܩ��T�pB��hp��&��O�eƠ��Y��G^���ș]r�t2�&��g�&]:�ɞe����Q9��&��.��ۨ�ˤ
(����2X���^V�H�������ϕ��9R@̠U��rU�����<P�ό\�����/�++��ҧ��@�B��3#XA�߈"�P�;H��� �?���|p�G�� ��5K�N���i�<�����W��`��n�/5 A����-̽/A����0��Qm^�k�g�W�2,�;�`��-�O���,���X���oٰ9S���z�/<���h�zi%L9�j�nu�zYЙMH���
�\2��a�|���(��pl�gq+elw2��*IfMѸ���H��l	ϔ�iC/�����5���gAO��ł������$K���iJ{!>���Q^_�3�x��MO�F��sH�/�iS��
�aC����}y�G}9�K�	�#J����F���u�Sk�"�$�+�0F A`�����'�<�]i�Z��I(�=��QqӀ�A�Bi {�I��j���Dn�̢f͏.br�����b����2�`������S4�Ip�RA;F�u_��PBa? H+$s*0%�1��!	q��[�*��Q>$�,��	�y�	�=�����Ys��=����uַ`�f�tpe�bƹcj�xxQ%�_<7��9:ڦ�}�A���L�2��d]��!6:ȇKZ:8A萃
L%�n͍0��<���
��-��^7�;��}R�8t���0�T>�����S��Y��s�~<��u��Q0P�;B�䊽�{����T���o�*>3�[�[A���pn�������l<�QTw��Iu���5#:�Řw�
̢$ٸ�V�[{�����.�p5��f�6�֧0�y	/�u"�
=��q ������6s~�X9��D\E��/���e
7��b~���C{���Ŭ1�0;��@�@E�Q ���J��&3<�2g�12|�D��̩-��@S4�7��uM�=H�O�Y��������Zx9)�6�2�c_w�j<�@��mVκ�#�P3���|���Ƚ}�*���lM_?4�u�5��7����?���MH����g�)T�575�A��Ś��1bk���v��_�Ax��+�Ɓ����W��=32h�`��R���i@����,6���,���4��_��3TLT(ӏ=R^^5�GZ���S�z��z͢'���t>��"h&��_G��L�Tb�/f��ڿ:s���� H$@�p�jK!]Z>)�X����lF���j �&֙5���ƴ%���gC�As�()ل�>v�\����j�^��>_28���q�s�7k�d�%��X0�� �� {�2�;�|= ��>"=��/�=�@��5���X�V<� ���-�E�ac�(>}�T!����Ѫ��䟹����n0���dL�6��~����&� �pw�),&���)ł�)hj�`��iYJ��@.�=ry�,6S_P²�]��C����}��h���cv8�>
Ϲ{�0
�Dx<���
)�5�i���"NхIf�E
μǝ�D"�Z �.�b�,2,���I�f�v��,�c�J�4���4�'GB���fGJ��[� x�W�w(���Clr2���>QRy���F�x�a�+�ܡ�OM< ���i/9�M�g �<d�A X�%�q�+:	��B��|�X�ʑ���u���ͅ�XSڽ���B��;1=��a�R�[6�w	�$������ƽ,�_���fxל�jҫ�&F�zK���+�_�<��8$i+�^\8O ���4�b�(�&���ү�9�̊7w��	�����-�&���J�[��ם�M5��CPv��OL��� 
�A�%�)8������؂q�8^3!�Rx	�걪���c�%/�}-4�*[6��Fq��G�b��I�[� �d٣]H�ꁽO8{X�׽y"L$�����i<zzӚ���A^��},�R1;]�*TY�r���u�z�j��
pa0�/җM�^I�p~³����	�K��5I�S����uAM�!�_I*-5��&=�3��Hf>~�;WkTӴ�C��8��.t�Wm��i�eX���&��c+щ�^F(-Q���4ۑ��`��{��bLum]'��c���P� )_P�6����;_7l3V��+�p-�_S!�&;Q�X�.��n
�pW���@����''���p�[�]�`�Zȍ�,V��(֯�T�Ck��i�:�Dcԉ�����fU��]�ȟ>k�+vv$��_�$݀��w�ĢpA�ɻ��t	{Ïϫ�`�RR][�(�a5��RTќ��*ç� �t���Y,�����Z�`�{�B�#� �{"���=����������x��:'c� �F݆e��5��w�Sx�|ն�&�D��Xb��z��pM����L���yɃC�����^��N��� RQ=(��V܄|<:M�cV��!�C�°g�[�zŦ����qG�AE��#�^��Y��:2����N�khA�<��@���<��ˣb��R�kT���I���"�?g�(2'(��¦�(�3�)Ew3�e�r˥z
�X�9&5s�j��uIy,���'�|�[�ұn�6�z��U��	���~q�v��R�]�fy�㢯͝DzI���?�*������Θ�Բ���v�j2"Υ��FG<o��Ǘ��<f92�2ƍ��%�m0��'U��ge�<l%>����y-Ny��O��vݲ�4d(9�FP���c�R	�Hx{]�Fg`��L����YT��Zw��|i��D�B�H�_��?�D��blSS�o�w���Be�L���p��m�=U���­0���A			Бq��,�C�F�H�5��3�>@B�]L幞}��>�~U3=��0�-�]�Xӽcne�f��ꅛ�,S�;�f���i)�B F#�����"�xȎ�ջG}T�4��@�;����I������R����Z���[��Re+K���pF���V�1R���"Y���pzD{S��̾ �+��8)�bh�����݌�c�lU�n<��It�Y�4�$Lņ]��{�^a��t��&�3�����
e��FKD/ؖ�ZQ&Gk�n<�N>�P��@�7�"���Ҫ=y�?� ���gݒ�Í�^�9D���fo��%{Т����8������~�3_+H������JZ��rOE��(�+^���h	��hA�w؅�`�
�� ��S<��5b65ͦc�Fm`�F#�S'qR7��F#"��L� ��!�&�E�,�͝�agH�Z8�g�� �|G�������0���8��8��?�q����א��%M���,q�L
`z5p&�tqvn$���p&��~����n�h�5�������f!_�z�����Kе��ݜd�صf�!@�u^�.��EG<v��%�����[�1b�>�,��_�1'N�i;���M��N��j��լ����X�`��)��3
N����pR�����ըW#LG}&eڒ)��4̄�c>edI��SP\=����I�/��P�,�(�a����1���Jsg<�p�XF|3є s��+���?z���;!�>���'��
=�&N���v��a�T����]����nk��֢3?��c�}Z)|���yg�j���0�y��/����|�'��TċʻY��s��~�S���6�{ԭ�B������@:
�%�D��С��F���]��,v7D!u��Q	�����ȫ	X3	Ki�jD�����%�ŵ��&��������lT՚1���
 �0ɒ��`�������(�1�4x���է�������,E�k3��>(1ǐ��J��w��%�/�C���>�2:\�R�X��y����=d���k*S�B��T�䉌Nƌ�T�r.䪢�PE�;2����}ܿ�;]�~��T�%d�ɲ�:�On���)t��Ӽ@�~!��� ��g�o�'����>����ԞM� ��V����ƻ�n���42dЛ̏��m��y�[΋�$Ä�x�_7)!�����.�׌hx.A�٢��xG "5��J�%]��w��@������wB_�!º��xL�6��&&�����#�3�
H�Y)��4}�m�.��י���!Ǎr:E)|Kd�^F�S}��j�	��#?�e�S�Yғ��\蜟<�J�R�o$� ��k���F��5{��n|L�=��?��zmGG��!��8�$� X켷,=�u)|�<m�:�H85=�du2��a@�f��n����0��a����{J,6ۦÆ̥�����8^���k9��0����cd������rG�a�����;�l�&�6����K=!��	��I�=>4mD��k��nN�64�a��	�����ɓ�g/"a�����:�E�:Tބ����<��E9���;���2��Ҹ�<�ާq�7F����Oៜ�VM��oGb�ō�%��P�Qΐ*@�$��յ&��JU�7e%|���Q{��Bh1R�A2���p4<z��(F!΋~�Tk
�A�cx���t�x��m��.$c�-�ψw�����`��i�4��<�/�\�B-s���x�O�^a��e� |�d�kR�Č���/�0�.�C%��O������]���D���!_��y����E�ei�S��X}�]��,�-�l��D��ʏ0GYA^}ޭ�������c�}��PR�|���E�K궒�
����x>�q��iU��r�9�\�u w��q�����'��ILS���Ƀ��Y�AA�����-��E�S���Y/ٮ��I���d��R��8\hܽ��ʃgJG�q���8���ĸ�	��/�;E6p��z�����i���Y�����+��qrR���4�V~�ĳ���x���V�����H������.h^u�* k�B���p�=�3&�H2�xn�d`ߧ�z�����Ė���}q����(��rA`�1�Y�̰tA>I��q7�*�:�[md��)����OA+_}���ۻ	f��b���	����A�r(p���\3o�M���������+��*i���|H3T��-�̏v��JxV��w�֯.L�%�,ip��,EQ5��[ӑW��������p��|z5Aݚ)!�)+�,��_��Fjd�z�4�c�T��2dY>�*ʹ~���~=�8��AA��m����럊;g�w�&��m�,ٜ�r�BM
 '/��K#�'I��k��0�'ѻ6:�M�KT���V�ǋ|^��(BKʹQ $�&4�iL��7^���N=��b��n�9Q ��$+'���i�F�g�t�� �f��*#:�g��kO�W��_u��tP�"��=�ɰX�.���kKǵ�⾾��	>�8��#L�yU&���=�lHOzP0����[�5/)(� ��Tk�d�D�k�o�T�z���}�
Q�uy�s�ϓ�ݠ��m!sf#᛻��d��u1�{}�!�K'�bV�Ҷ��_��0bm9�
5�~�2�Ήh����
KJA���ُ�p�����Ȩ���@|�Eg4}t�
S��[b��<���j������_�Ir�z	�ؑ�jھ?�-���td�kb�DeGJm�~)��B���bQOs+�-[١��N �5q���V��j��s���ק���ĪH%G���t@��2.9I4j����U�������O�aBȉlZ���K����f>s
t�>o2�	�~��_�`Q�m0F��?�)p������C�K0�9r�Q�zz��z�u��i�f��Lt��Cآ��־P8*`��� �T�����=��Z��&�s����'v��\Ǩ�!�)���l���*��9�5k]r�a��}�Mʴ~S�P��3x��k:8�^Ȇ0Y(Ѻ�G��M�����Gr>��_Q��o�� �6�L�k���S�k�[���L�:�e���{�B�������n;X��4�p�� 	��K�
)v��j�����C��upHsJ��0�c_�//�zI��!Q�RrK!�.>\j��>�]���]]�j�Y��y�ݼ_�{�{V�����2��������*��^˕+R�n�A�9y�[Z�q�kN�2�G�߳��CX��[m'>~�%��fR��]ba�+R�B�qB�f�t�+� �左̍�R$�4n��XQ��p^����5E`dv�
�I3�G�� ����(y�Q����߭��-khe��cP�p=L0�Nޢ��U�~���@�~�o�c+���8�9�3����X&2�	���.-Ա�r�=V�����b�<��;�-��@��eրU8M�b��H'�(�c��V�^<��.s�+敓g�lvq�j "�Y�;tjZ"���Ԍ�1J�����+�qX,��r�M*gc�<`d�&�N�@V�a�z��&�}#��TG��^p-
l�EU(❭X~�e�P��+�J5@�}*�6��䓩��K��W\0���q��<����'�i>�Aa���	#J�e���Z�iQn���R��Ӻ��weI:h#_F�S�-��DԾ]P���#	d��" u�7&I�&��]����|&Z�~3^�[��(�`�`F=ꅃ@��[޻=��t����sP�SCH�=D�26l9;��"/$�iɔtpI����h��϶���u]���^H`K~z�/B#�c�ƴd�(`y���U�g�H���8��U6�	�Ų���Ӳ�hܠ�v��ȏ�D���71*ا:�%��WB5��<�[I)���3@�'��2���*��j,Y�lw����LfR��Dh謹�y��DY��~����Y�ֶ��u�_oi)�$���U0P���=7�KMq��y��,8^9��u1��Rc�<2��]c,X�0�}l�}������
�o]^l1m}���d�XE�P2ť����l�8ơ �]����=鶎��aSt09a4 ��EV�E��d��JB�\���6�m�ؔn��tɓ�Y�䑲�����x��ר�s�l�!�ϟ;�=�vb!�z&4�R'�.û�!�	���'��~$nH�K����8�#���E����:Ԝo� !��i��/��-�*�����+W�GZ:���B���5S���ե�DI�;�Z��R�0�#̝h�����b]���C~^�Lޥ	�kP$3��c=ә���������Y��8o�$�h@u\O2u@��u���j�/2,9���h�Z�3-􊌢_�UHް5��y|�~��Lm����,BeyC��y�ބ�ء{�-����3����@�J�����Q�Hm"G�����AV��g�A0�3��[R�,(]e�6�Wl�������)���+簙�����1���A��Rs(����G6����9�UP��I��9�x6�Y�+;�D�f!b-��Q]_����������L�|o%��v��)t��<I�괐W��aX���HҥG��ջ锓@\�RX8+�&��ǵ��P��ŀ��Aۀ�;�i�v�b�Ir�Bi�����@���b��oc X�Q�(C(�I��~e�z}qVZ<��v�>�Eb\͞X�?©��9��}ʄ���\���,GgC(���t�phx�r ]�	a
��B�n���6c�w8�-ꝸ)�pHqs.�1�����뻼S:/V�&A4��;l9���x"��"$��� ��J�"��'ʵ'��pr,bO`Q��R1�~^G��M
����LԪ��G�z~twt,�+�'b����
$ӉP`v��0�x� ���������)�B�[�{�B���a��U��/16����V����ZA��	� ��:��@2�K0O�s37�Z��P�(z�ҋn�����G�nUc׏��I��Y:7��y<�6�}BԶ�g���E����pf�����j�}�JF�V�t�ĺ��q8z����"�e�įl��� _�0�(��ʓ�q��w���U�`"#h��4���u���UE�pb}3�B���X���'�3Y���&����u���l|	��Ԡf�����;ޱb�8�>RGK=�J"s�y�Z�g�'�V�ޓh��g殮�G)Ü6���r$��dj�S~ oh�T�D��Q\TM��8j���4�~����U<Q���.\���(�!�d������1��z)�G?�m&��K5ˊ\X8�k���$ �~Y7ލ�L�.R=?��:frwW��fsU��ܣ*�@��E�M��~+��ɺUK,M�<:��� ��'�%�xVoa#���vV�V�;t����a��Y#��=i <��j3Zʒ��U?�r�~��í(nv�\��Ǳ`YTc�Ҁ+���Pk��'t��3�����H��0^�w`h���E�R�Gz��<����U,7� ��MH��>��\�d�P��*�:�Ā��
���WU��;�^�AYܵ��M��!W#�.N=�Vv��ҡ)��_��?%�K���c!@�j\��s�@���Pt��'��<0�TI�e��׿N�����%%�Q�����`�S���ê[���S����ǘ����U2�d��s�j�F����zŎe�-�`�is�sIr���3_l%���)�X��N�H��~��ʟ�R�P�tIm/�+�d
��w�#Pt�K���m3myZN8qD�9�d-VT��<��.6
m�.���j��GԚwv5?}/5��T�i$[^�Z�hAhF�YC��,��Κ3�DP�$�� ���9�R��W����D\^�2��:��X̡hY��������ꖩ@�	��|�� R�+ͩ��q�D��No��H1�!P��A�Y߬�`�V���^�eS��5q6
��^@����A�ɑ��윭JSH�-�MK�g����d��%��<��́�<�?��g�,^��F��I�h����V	�/JR�\9k��
�)���)5T#*x�D�..봛h��xJ�*qf�ĨPXJ� ��qe�DM˸�b�UD$7\�4p�ڗ�!��q���Q��-Ѷ~E�1���	��Qf���M}�e��c�6��n"P� �3��P�%ƥQ-<��[հ;+��B2m�V��P.>8���b됳��=�ЊOњ�L�O�'j%t �S4C=П��~����E �.����Û��0� yuew� � �R���\�����#7�p�6A�����w�ڹ��w���ݾ����ǌ[9W�m�
�
ɵ�=��80�\$�*{Z�|��s�9�z"��lj���6DQi]N��^T�"��wI����(�;�J�C
U�y��0�vZ��Xe�P�nay��Ƥ��Ng_3��c���� �_��L�K�{�o��k��FH��K@�UYEƟ���˩�#�<�f'9�R���brG��M���Ũ�K{)�'���rf�:QT�3T�L�w�#�1�[,f�;`!a[&�뗫a*M|DD���	�.���ܽ��#j��:�"��vތ��ԝ��u���;�l����������kǊ�*�n�m"���g	�VaN99� .��-�u�k��Z<ěu�Iz>��E,&bU�w忇� �48�W֚�70�3�'�:�<���Y>)�h�P��Nf_턒�L5��W����@-2�8�s�Do3��##� ��`.�[��jJ�/�����>����$�M�}%��WTP\X;	�����;�� �br��	�'';�st��	M������Ud��;��|����#:ׁ��p@8dm�����4/�!`�����&��w1u�ͦp����
��R�(F����i�����D5��Yf�Z&�g��\��y�
�j�iÍ�ap7�h,�=�]#-�н����yp-��j#Z�Ė���k�aK�,��̳��_��>+Ah�;>��vi��D;���,fM��������3��Ku�4.��t%ԉ���SY�2��D*t (��N���Hȡ��d~��U&e��my:]Aa�цj&��aG@ ��yh.�E��6zO@Ȅ�����?���ę��ܮ�2��8�[![�L=�B<�C��W7Ӥ~����$.�e���
L�p&C�^|��"Rv��%U�{#�-��W|Y��
��G�VU�utje^;��o����<x������%�V�Y?\,1��/��ԩE�t�KhA";�@z �����W�+�6q1��TVv?���ک VJ�CƵ�&]h��{bK_����j	�D���h�ڲV�h��
��?%����xe6g��0�x͍	b~��*<s.��{�\|i�v�j{�*Em��o#LS�k�C^��ݶ���Զ\_�!�=?��IO4�M/�����s�)���� ��~E�i��S��\yYW��V��N��ܒK��A8q�sG�jQ������^�9�x�lK#����<L��� ��+*�+�3�wz��t�����P�6\����V�`�(�/W��)�L�\九�C���Ӡ&V�(p�?�4>0�5)���� �s�lE�L�Efr��m�|-�G~b+B�`!�"g�
#�} e����sQ���V�/�%�>��$��R_��M���u07�)�qM� f%>z��xF\�k����h���p�[Gel�L�x1�AO��l�}C��#p�ހ����m��'l^}��nN}!�$�����*�>�����3�X6�7g����=�S	V�XM!��H�߸j��7q9A�ϫ;�c��2�z��RϤ��o&�|���?��!���~��KG�3��/�k��d��r)8}|;��\��ZA��~j�P������YO�Q�+������!%ns���#�_n�-�m�|_ݱ)�Pu��Z���`ͫD@�rإĥo�aY�n!�0��������W��G��m��w�be��iMZaT��q1�fr��Y������na,9c��>���\���Q>���乹#��&�h1�b�O�肵��-gA��I�B���AFX_�V���;m.rs6V
�'�Y�+GҽLI�7Z�Hb뱚}�V�4�g��Ax�U"������eݱ�>�GbO�E�D=?2Յ~�9�b������`<cu�_/e�tPHa�a�)_�4�|[���V\ִ,'�0�o�q"��.�K!k���0���k�ϊ�n��b�h4��|V�]�c���هVZ����~�A�:>��������(�4F��^}�<�dxB�{9��DQ��RەG��@+���e�́�n��f�I�c��[�ID0m��@("5�-�xg(i\Z ��S�,��Z|"5���.��'>ĽY���)9<'I���
��Zt�0��T�6���%<�&��<ER��=�0���B�Z-"B��I[�d���c���XI�Y��E��)�`*���L9�:���Ar�P��^�ð抉O��j�V5��q*�L�t�&�6�[�B��,cϡ*��Jϔ[m%�{��Qrx�PRp���U�6���DX(v�ƨ�/9ą��ڭi�b�fK�J�&�w��7��X?<�twA�$��+��(��f��ۥ��sk�xvoHK�k�4}�'����H�S=~=�������PV���j3�RI�;�F�;���%8����D"��7s2E���T�H�w�i�Jv�����0����|��@'v��L�ۚ8q��?����CJ���f�sH�z�h��-��v�{��.0L%@�Dn+��I��E�tD�hvI^,�wU_�I/p����{m��P?�W�I����������Ob��@&:�Sr��kn�C���|t��\�ܥ�J⍃\o�f����H��j��m���M��moBM���a�O����Ր��`��Cر�l�Qb��o��	,��n�DG�u<����MpˁD�Z9=�c>�cXgcD�1��P������D"����l@b�0π��n0���C�ْF���}n�]f�%����Z��#G��/�� ��f&{�X��`��:P5k$x� ����2��6B��:A'9�tU8�g����A4�N���tqk��Ah����ߏ���@=	s��iA}pƕQ�� �&�e:��".i�%�7yq�z61j%�\D��}�]؛�������F,Y��?��ɣ�`��,��U��o�3�)��?k����j������];ǅ�TU�7/�F����S�%Ƨ(DN��Lrd��2������qe��l�<�,��d����o�ͺ���E:ǝ^oq�s;ȣ��8�Tvh3�´m�§�d�I� ����0P����ڐ�$�O��*�m�ow溰(�,�f�I�y�b�.1Q�J�D����>��s��F�&�Sv��*�7d_2{��l��M�ɸ��䜭��?[@pd��Hf��J�[�s"�S�	������@���;�p;ހ�Fˣ��_k��#�*R���V+B�A�I����{'?;KZ,y@C��QcE��Ө�E)�T�����r&�������aJL��~g�����M,�Ij�҃���;5��a��^@���_� ��k��K)���r|�j�jH敏�����ݎ�PR�a�o���4�%֖��F1�͛��,9	grS z�����M{�x�� 6�K٘����d��ò��P�"=JJ�QZ\����ڗ�H'm��͏e�����yM�U�����tt=^<u;�³*��i<�^��/9y\aMA��R�C����cp�0�(��$�VA�4ù#�?�Jm�?6�,<1W��	���$mXk�v��=E�Q�沟�O�4����ǪOü��)�O���%trN:S"�&��|� qE�F{�zգ�緁 ��U��3�b��|�s���|$\��Q�䫁��u�A����N��/�8�&��\��YA�ͺ;�N���2��!_�I�L'S������T,�.��\L�3�?�i�O���Bh��i���H2�ώ�Cϫ�~�^i՘�iw�c˱By�xEW�?ؑ��.�6T�����j�bgu;q=tn�UWT��K:fW�-lh�u�If���x����!<��P�V�tޔ��൞!a�5 �2:<���2�:f��I@Г�xM�0g��^8��܏Ũ"����X�wB{'�^ b>�-��
��.�,]�7K�wy��ܘ�W5��R�K���	�A!&옿��q�wH����\���H����A�?�
����w�L��r�T�k��6g���fM�b&o�L��Gq�&�|r�'a���
�l(��¦�aVjm����m�ь�y��b?�\��b�8��vvE���%�>�§��~	ޞ�e��k8��RrK�PĳB���m��t��A��fH�T-+��DH�e�dW��4O��:������'��1���|X#F�.��^�#u�%ʜ���/%�za�*��3R����T�ΎP�[�L��C`���c�7(� ��;:w{mUu]��i,,�`,�k��A��ʰ�j���9��SR�|��ß}\/ �T��=K���UQ��iA�B��ʳHO�#0�#�f�?m%.���������#?�m��>����O/�W��,�����(Ls8) ���o|{w�z�/(��>k�鬒d��8ڛwLjzZ˰qy�g�]9���"[&�w}ľyN�vj�p�D�,�[mjuS�Jg�4��%���9���+ӆ���0+�:���./ �|Br�M{6���S��n� Q*�sfFJŷ�pצj~��ɓEY�r��݄.�gSN�E�����8$�����m��F�\�$<rֈ	���6h���$�~����2��1\;-�!6��d��A�P��<#�ͼ�М)�������|y���G��(�YCz�VY�h.�:i-�樂24@3`�_>cr�'�ȴ�%Ez�NS<28M�o�����p�t��/�D�\�K�` m���s�b%�ͼ*b��-bHP1P�"f�lF��l�{�M��^�˿���U���<q�pJvV�#q���j����8�h�;�<}����5��Oc�.ޥ�0���u�-�bw1����������ę�y��s��*"P��x���H����͉�)�Z����${U��[;��$�,[qӻ �����������u$�<��#Wa]r5r*u�M�M��k�V�@�m�,VdtV\�n[��M��s�S��d�%/��&Ԡ1,�9�q�-br�A+�m�~�M֒pl�[��蛸A�GgHjc�O
��Ƒm�g�J9!��b �N�Pc�k��|�ǫ�@�qt�);:!s��pHXȧ. ��L��#�������k*��`�sĿ=�x�mȷ�AA)M[�ǿ�Vu�ߊ�-�#WP�a'���=�$ c&X�oBQb4~o��:YRHJ!f!�w�_6�t#���h��T��<�����Ϳ	+B��剎��%��ǡp�:45u�e��t�G?$�u�/�Z-��'�+�Y����sY;������c9�����F���e\�Y���cA�H<�� Oݢ~O�������{
$}YȮ:�z�ҽ�p�B^ᦆ%����ٳ&���F�|��:}|m�8�ͣ0_rہ�]��ז�أ�|�_q����'_b*��Hg���\�;I@]Lh��J�@��o #JgM!�-���q�O�b�k�6�*��32}n'����^q�Rw؝�%h�AY�C!w��ѷ�E�<��+H+�sh�rMDpPx/��
���eea�J=�?/J�^�߈��=�'�1��뷿4r̯7;�����
3~Q��gׁ�YI&p7����8D8���Q?U�'�N�Cg��W�.j�p�ix��j�޸#��rV�
_2�BD��_��tO�1�~�>�����uѪޮ���O펽E��*r�J�+Z��Ɠ��X6����b�������|DqJ���d~�"W������}�2]����#L�*�	V��.�nz�8z�X�����S\U��g�
;Vs�2�JAb�@(���D��Ғdbԍ-[�դ
?)�@N���xmm�18��`v���d#t�W��|w:qƚ� ����@�&^��>�"*����.#;~F7U{*�W|h!����đj���Tx�y���-ұ�;e̅��Jk��y�C	��|�ԅD�0����8���0���r�ЈщF�Ў�w�ߍ�Bb��?Ӊh�����e�n�a�ê�����3�����`|��FK���7�\tJ)�}���^"7�j�����8�������]�mޔ� �(�"�U���n૷���B�ϩiG�)�W���L^ɫqj\�<�iq]�V9�m2��X���ĭ�Q��8�;i0v�@9���n����0�>���2g�w������R�
�x��U޼="_�v�Ck�x}T�D�_Z����\�aX|U͙ �p���`K�~ �z4aeۗ�>)���\ܜ��7�;���H#�-y9+�5� u�S��Z� �=� p�b蓈�k#L���j�n���ߤ|��ҵ|�lN�9д�4���xށ۩R�mZ���d#��i��%��a�@����U��x�?�j�0��2J0;�۾�bAA�<���	�oI�D�**"_�[F-i]V=fT��*y�QJ�וu����~,&�3˩�oʬ�|��x	��z��ﵪ\(��5��P0G���ߏ�nc��!��r��:?�N���H�#���cf<��8T�X�f��1K8��{���|	'/�?����Xxj����U�qHs�X'\�m4�:�,[�!wM=A�����)#zZr�;����b�['NX��-ޥ�ی��D:p7�{^�R�t>\�CU�)G�U��J�jG�����4g��﮵�R��<+�DX��\Ё�xu2s��,�+��
7K]uzd�Zj�	�N8l�Y��>�E !��k�mל�I���,��W�S��\��Y��Yh�R2+��тWu���C����Ұ����9J�*�����}A�㈜ͺ������aE����W�5��(��4'ΔI�N���B�g�B�'Ѷ	��㟓ʕ5c�rf��],�t�Կ�]��dxȀXk���?W��c�`�Ȃ �3.>m�ă_���}�yH���}G]sO�|�`�2�:�,�g6����DȬ~�jQG��b���N�]SH�o�10�g���o�����'�ߒ��ٷ sZ��,���1��y�䦚M,-`���^rt�T��ّ��۱��H�����n����U?tZ��$L
�ɗ+xO�B���옚���B'jF$}��X�ǆ��&@�j9,�M���n!5�3ψP�df9#����'��t��P2���y˲3;{�xm��GFo������v$�/ߛӧ��7��y��oO.%��צy^T;�jF����]c�DF�*G��*�S��bʔf�zc�'��~| ѱ����N�D;%q
.b2�#�Xc�-����c�ʛ�����8?;Zoy���|����M��x��9󌯭Sr�ܢ�����������i�Lr A�%Ci٪�"0��HA�wr�&?L��Yc����z���٪�YR�Q����Vv���d`�: zUd	�&�~�}�q|�� �����<n;Gg�<~�S;)1Q�����0��"!�"�Vl�y(ʃk*�x��tl&�\�W̽	�}X���b��»�:�B���h0<m���"�q�Y3���� �S9A�߮>'��Ȥ�����X6ɱ�0�2y��p����i�ҭ8ɼ`�������tFڇ���:�^�ix���\�����*��	������b2�z�\Qs�Mb�`�=@�l�+G���S}6+�â��oE>|%!
6�"��~z�Bca�i5�P�'^�!�)ݚ�[E�q��/�7I�jBF�+¶�� Zͧn�h�W�k�}X�������R��� �Kq�'�����b�V�tkS����N$5 )�0��8,�B�~��(6r�^j0Z�@&�S!j��3����K�Tß5���H��ݹ�R��p��#���j���A�8��л��f���^� ��ĄB���pM�/x�J�N(�d�=n��N�ɆR�� t�\�b�PY��!�Kv���ʓE_��P��|Z��^�xF����/}z�( �y7T�zNh��~�1*�x6����x�����`P��=^�(}ʒ�q�t�L��H9�Ҡ��j�
�V1�O����a�K��u�6��d�����IJk�y��e�L���҄t*
{U�&�B:A*%	*gQ*��&��aL#�������"�r庿��_d܃`=�3�v����?W��!�&=�D1����#C���o�J��T�������U��m�8��I�5������:hn�d��sE����i�x�]�C�۩-�^��h'h׷D��"��f�J;s8�Bu�7�![�=��t
	����m��R�6�����x�$�P ��v�-?���Kj�qqhf=�!�6�G��?��^zu���gwZ�/j���7dţ.L���Z�3���^���Wz�|>ʦ�.�[��Q�wIU�M�Z~�rJJ��D��S��K�gk
��J�3e5ٌ��&����jg8\@R�3��[� ��h�ҿ�B��zċ��9�N��_�`m�6� �5��wҜ�j�/��u;�ĕ�Ȳz�v���0�bW�� g>�é��R�N'�u	Ҍq+�����由�',��t�7'�@=m�6Lw];j�f�D�Q"+�@�M����K� �o��U4��Qtī�ͲB:y�ʚw�8��]s�O����W�ˤ��/)����ǅ���Y���䂯�hQ�kG�J,CǷ���r�2�彗���z���i6�j�6�>�����p�"6��%�"���^cY�����$�6��XjC�õ`!�C}hD�i�D�rr�ۼ�`�BGؾ�Z���#�^�*r��Jo��� ]���s5N�%�M�BY�g��\���E2� �ObN~�ҷ��l��'2�t�����i��3~sv�u~�Q �r�5Gq��F낤��&\��� Ŷ������C�Rn%]9ma������d8x�A�
��d�AP,��J�۰��|�Lَ�g��<{���� A���Ø�@,0K�>�q�㟸� ��j3W�i;���,��c�Fb���;?D`)`86e<�t�_�6�� �΢w�(l?�"�)��s��{�QL�r=aJ9lP 1|s���B��0`�@�G8����c�����x�=2��1�8�5w����C� ���rm=�IN�ӁԺq�9��>޶�}�,�X�!�T�!'Lt�ݠְMث!!#ݕL�]+�O���E��*Yw5C{�fo`�#�~E+��2+��">�eej�*�D�F��1��O�p���b��{�Y¹��T�R׈��0H�!��H��De���QL5f5E�P@�c�Y�{��������wY'?9wwvy���AuH�K!��i.�n���+۪ f�$�n��.M���	��H5L5D� ���ˌ%Y�[pjE��s�o˪��;6�C��n�J<��d��}����q�3����� ���ZV��8�obV�(yƪ+XV�����|����t���Ҹ�ot��Zn�{`B��g.ϖ����&E҇�����7e��<�~��-��9v�����L8�UQ~���>�+��x��v�7hA�\�]���Q=VduLw6DLٚr9_B���k�hpS_GBX@��W<#/;A��n��\(��\2F׵a�
��u��Up�[4Q���0��O7����	8"D��n� a6~��,�b��'=�p���G>�a�"7�I��?��7�"�4�1�S5�����L���;��E @��Ĵ�8i8fG�eLF�Z{ڎ��sD��-ힽNU��R}��wV܄�s��#���Eq�E��@vȦe�Z�r$�L��A�^�e
j-�]�E���%Y�OvbC�Һ�D��%P�{��1�����ܱ�4뱓���~G��zV�		� 3N1���'�&��os ���	��x�`��������g!���'yhaD�_���h�L�13�-����Th�0|�uVSť�%�����(�+?5ˤ�"|�hB��9M�mBv#\S��,�#��5���l�-�����fm���K�N�I��M^��a��S��*IU�B8�5�u`!�%�<��䈰h�-z���&=�Ͱ��[c����Tg����ި ͜�(�N�~���,oL��.�0�b�>_����8�w��(wLd�E)-�2^uL(a !�.Pi`��|(��r�L����ե4X�E�v�.V�'MSu�IH��RH�c�F�`t�.�:�����yH��t�t��y�ÂG�_
�ha�ѲY`;�%��Nڭ�k��lE�و�I�F�T������l7��G#���q������ �W���$�{�%M1
�)�9�al�%���v%ب��6�g��Ĥ��:��=կ�:@��^��z�~ldW}U�����vt��_n���ӳ�G�O%�pr�*BrsnnW�<�O����cgư�,W�u;�C�	U��F��M�C�b ��3�؀醨���="�:c6mdJw�T.�>����g�ٝ���f�>�@�9�:{O%χ]����A5�(-�fW�;��;�K�5i��1��r&z p��>��%eIP(N���2:�c�U�lwӒM�Gt�ij�B�6�hı��8���K�e�=�H�f�����3�$&�{�!dJe,L�Ρk0�A��*{)"��|�M�1��wF
Os��w���㓓$���Ⱥ��Ti�V��B2ޕ|
7&bF�����&�:,&�YHvyb�B��7���c�CiK ֊T��W��b��a����v�?D���>�<�F�!�9�Û6͞�	��oO��)����'�>9٥b�RR"V�%�!sV\�;��n%��;�v��)Ǐ�\)W�c"ޫ�UՕ��p�X�	YYv����i�ɣN=D�ϑ*E2�o�R�=�M���"�pF�5�����X.��ӆ�H0��2>��9���Gg�	c-|��#2��
�� ��($���Y��)�ŵÅ�n�h�,�`!�s��#DJ�v}�J����ϒ�Ө��kv>}��*�������E���)M-L*��Ӥ�יl����(*�{�Qz���B0�PAqZp��H/�pc��f��)�
�X�N�\�)�`���\%��qu�gڨY�0,�gG31V*x�������ḡA�2ߛ�����+97�g	};	���50�S>�֐+	uU�^I�H�ub
DK���[�uT��D�����z/����آ��o��ۻ��<���B�1u'
�0�3S2��W�c!6ŵQ�O�9��{���s��f�L�>�`����z�Hj]�f����{F���$���T�/]P�Q��"���^��5�>-p�R��"�½G)^Rzyjg��|G��K|LS�����=���B9���Y�jx���=�1�k�I3B߭+�㔺�l��.�!���������9��-�#���D U�^��y���5��/���m3�
�G��DXہy@��Y �-[W)��D����v�~�x;�����c�&�߰�����F7¡<�	��&	JWuF�&���U����9�͆z�jK8�:� Nоv��w(kDC�������^Ђ���@hHiH��J��O��Tz�5'ؾ�����"�X�ω�|:��� t4PGٵyF���_��}ŝ�1L�${�u�Ӟ��<����59�H�7��Ag�l�x���l���U1�b"��*+��G�����P"�ڡ� �9��OP4���'�'=�$z�'*��?�G����P�;�i�Ѭg%%z�Ӝ����A��&�����spV�\�>)��W̳�d��Eh�nD0B�����݋�_�:�D5�(>���g��L�W\nU/\-/���Ǉ��E�,m�,��Mq9���Z�L�[��6:C��`f=�F;*Ǒ�5
y��9Y�޺e���}k�`����P���oBOO����	��hLLcZ�>���r�o�4	�os�?�Y�6�T��"�U������T����pc�-�!5���j��Ho�D���4��K6qh�����+���l��`�Zנ4ţS��G4��3C��r�w���Y�ݷ�=U�{$�6j(��%cCmE��]Dǝ(g٢�`�yDX�"�/������H׳����@�8ف�-+�f��_�n�o�b��	�S�V�D��,D�#Z׶�1�����ؓ3��^�~��F�0&BL�D��&���
/ؚZ����ձnܓ������H�����&v�J�����q��C�C��A����HMޯ5��zm;-�����-�|w%ݵh��%�ӄ��&ҍ��7v��b���|o�Y�Ha��ט��8HL�$2#6�Z�	A�0�N縉�i�f�-&����X ��~�aLO3��3u�)�������כ����|�ꥌ�/7(�9�)#N��Kt��ck����X<j��J�go|�"�˷ƻf�$��r6�'�<�59��}�J�����9�5�-j���^O��X;=`9*r��7��׈>nXXQ	7-1 �>$=柴�\�V�����WK^�`�c��3��'; 6��e�fz��j����&87��4f�k�eV�N�:l��I��D�U��J�I�6Āܢ=��.�͌�F��}��zB|t�������Lb�!�	�=hf����Ƈ���wK����1�?N|8ML]�!��/�y��W�L;���'��,�I�j�rKD<ϗh\��?i�]v����;l4!����齂`��� �n⻑ж��S*$��H5ݵs�m�O������K�p+Z�`��q�+���
s�v�n7J�wXs�I�|��B1�.A��{��fl��G�jL� %8��W������-����?�H����g��h�l�� �^P:�WYI�Ar��?9���B0G��7�@��=3����A�Y����I� ��t�+7�T��s=���BX��j ��穣�f)zu7hfT�b(������q���-��586F$�^����"^�1��É�2��,e�
�W-9���n�2��L�B0���.�+�.��j���� f-�D��n�N5B�:�AV�ML���Q���S�k��k�G�t��C�&��(�@顾R�>��߁�Hӱ�I�n#��T������pop҇�����C���n�ZP)�Ǽ�ʫ|O���h�S!��I��@+��AV=�3����iMCj��HH�ヾ���(ND#hCE�j ����&��{a7F	0G��0�>��C\z�Ͷk:�(����1������4g7O}�fM_����}�?�q�}��o�x��,�F6_!���^dG���wx��5x�I�.S�Gޜ�>�z� ����-�p�V]/!��Z���Wo}Ϩ��q�Zo\$����GN��`|�}���,��*�C�\�����è���	�����B�y���rk�Gt�5�3R0 -�`>g�zATt�p_�bF(�9-�v�-�o{�[��S�\�9���~k���]փ$
v�G�� ��H�ۆ�0	Pw�C�8�%���[tjB�=�ˣ���#K���#��h�<�^`��b-3]�!��L`�&5���k��MN;��O4���V�յ�Ykdt:��MQ�4J���lZ]2�SbV��W�������URʘ��u�u,N%�.�})�}v<t����
(6����;i2�K�E�q���NĽ�Q-.r���!r��"G"C�F����s���㥠�c+j,�ɥ�dh�d(iԴr�z���Uy�����y']�SI��(�� ;P����A�i�&�S`����v��a2��4���I!�{�MF�T��^wm�Ļ^���tn�����fէv&��O��8�_��`��#J��2�Wv�s�OV�i��@�* I�1#�5�2l�ΐVp���[mX��9ƒ��3#hat%S�h"o)O͡_���O=��+�s�G{�Ԫt�C��ye�'��v��6��p�Z���[��7f�EI��@���3[��݅�N9��h"��DLadNV����o��Xd+��?:��H>C��g|�BK2�����.E�6��l����[�I	�����e#-tR8����)T�h��d=!�;ZA��^D���6l��P/{����&���:�p�������"�y %%}``R���5z
񚹟�?��R
7����?l���i|���x�Uw2\������P ��7[}@P��bւ�}�Zs2���"5��7�ĹBQ���t�T�Z���TS�r/�%��p��+I���	M^b��D�?y���I�2��Y=70���\ȷ�y�V+��X��"��_IhH��C�zƨ�v�~�^6o��	B�r?\��|[��x����)�t��<UZc�<eWvB������u�Ԅgy._l��?I��+�D���q�<������-���\[�Cn�$og�|���-��V��*�ϼBM��:�
���KRJ��8Szyo��}=<�����?�w�9]oH��f	?�M~t��"Z^�嵣RJ��3i��\�#/qa8��O�)0�����t�~�+�S��:�2��C�&.�W�=+� �<u$�a>)��������M���Y��i/�g����wۚw�#����2�K��ub����L�r�2=�",t�Z�~������b�HjJ����0ێu���~���J��u�?f��mY�v���ߩ��w��U )��7x��6]�͜�*�A͢�\�%)�ӝ�qe��~p-��:xX�����s�}��I�?�.���9����.�vRvu����[��Ȏ #�Q��1��o8O9���8,j�ej����2}7�@.ѻ�㾠���G�E�*$c\���G� �A�P9Q���Hdq��F�ov�!l�6O��a�';���A��0���:�6c?sB\��r�-��]��+^=`@¯��t&���7^��� �4�9���C ��`�ðm�P�I�g�{���i-D��E����l�G����})@q�1A�@�Q���BMU����#�%�xժ)K���0���H^��L�������� ��u�]g�P���%�i��g��SEwֆ�2��~	�`d��&��C��cD3�/����4���1ToI�'��]�Wj9R���.S��W2������#-A��!��:��.�N	z>��0t�ԓ������Z�I�Ѧ�^N@e3��0�ˋDl���Kc������l��_�W��'�4{Xj�b䰼Ɉ��00�n�H!�
��0��C�!��1�E����!C�@H��Գ��?'��p8�����k���F��p�6a��(�cϑP��u7�i�M\<!`��t1+�"��2F��i�g, 0��8 ���wm�c��'�b6&�ᱤV"�������*j#U��;Foi��2д�U&��RG�)ￄgOT�Pnm}l�h�����#�/ϗ�����U+�g��o֚�hD����X�H׏�ѩ�:�
�))��ݸ�}�Ď7)�&uϊu��GD+�o�+l���5U�q ����Y�t�Wn3>+���RWҼ�#Ԥ[އ�$)�8@�U ���3���M��d���%l��p�rވ�.h���.��s��0��uw��C2�Nt\r� 9�;IT�L%R����=�a���7�4�ب�����E��<~h����'�Q3w�{��A���TQ%<'!�71V�ČG��
�	�;��{0��/>�M�>�u/��J9R��ʈ�l���j) �Y�M���޳#������^��?V�oY���Op�qO��$���up�(���AO��D���;�l�Z�=y�n<v�簵{�h��^{whN��v}�}Nu�k��$Nh��
V�z�3_z�W��&ZJb�1���aMb`������ׁW�쁝��vm��5�rδH�:�:�3��(�����f�V-��8�+�m�^�i�K�M`�;�=�n6�����<�u`�t娻*��7�ⱟZ&پ�oP���-�p&^�����������G��v9�dc#��
鱂�>��a\��q)��XiÝ_파�Rߌ���x�C_/��P���c������ϝ)�hG��^����eI�:R��i�,�,2u\'�s �ӝ��.�'ε��nEG�u,��B� �[��t?.c�v��)�6L29�������K%W����|Cpf&[u��A)��6�挀HG6;aj�ʓP��hM�7���N��oq��e���P������z����8����MyV9)����x�B�l?Et�W.4u	�O>�-�P��(Wm���.���^9 ��B�����6��=�%�z]�ܾ`�>>-^"�=�i�۽N��[��Ӂ���e�9��f 6� Y�����$T�V$�ΐDW(�Q�D����͟Z��P�jJ=�%����؎�:�F�J�=���Mz, Zr$�Z
0%­��(��&�Cv��.i���n�{�J|���N.
����31t0n3��F�����7Cq��E1 �����h ^Z���EF�{�| M��Do�F��h�N��$+p��M�ڛ�0y.DQt5_+;Q��`^�&�Į��0F2{���ӡ={���5�p<����&��@Zjp�ʊ-T��F�S.]���s^a��܏�ƈ� �%�ш�e&��S.<�j������m�d����R�����:S$���?ˡg�UT�c�OhW�m�냓�U�$]۰\�p�~�L��sҸ�ha�C�q ˧��1��uT�.�b7��@����J(I�`�θ�y$���!t#9�st���l�*^ޚF����~&��V*�R�c��0���%���)�.�Z�y�<�G�CY�q�����U�]�0;W`Z��>�b���at�>���tP7 D��E-ͿM���Nh��~��N	�ǿk���Ý'�'w�P��nA�0W�ws�m�[y�h�洴ohݳ	�J4j?~B�� �l=�@p�����p�/e���@���e��i	%
ȯQ'���tL�x4Z}�[��1ŗ��|��]��v1��y�ٶ����&0����	S6�'��@�(�Nt鸁iKC�������Kk$�+��B�ۜ"������c�.,'�/PJ�._�g�ʖ�g� �K�G*��.��[wH�QiA-���9��{N�˘�D�d9��֣�46#L��?8Lo��Z�n;�H��b<�#�|�k�W*������b�� 2B껍I�ĥ`�ې�F�>�m�|�ҾdH�����AE��o�.$B�b<C�-�*b�l�	O��\Y��@i��ˣ*�X����[��E@~C��*���lUvm>��8��:R�euC��- ʺ�Z(���E�x���&��͘s��{R��h��\\c��#��A�M��@e�� �6��b�9ުO��ȪR��[m��t�~�g�w�y��,T1?n^�/��c@�=��R�C�\��A?�ь�.cZ�ơ��R�~����GRp�/�Wi�k�u���}�+��]���Q̖��i�� X�k����D�ktT6J}ٺ^��Ƭ�i�����=f�n�$�"b��N�G~_�ƴ|��A�*�W�5��v�϶���
�L�j�*��qP�p���,������ױ7�*���Ju*�����]H<���5�f����?z�]͊9�m����f5\���_1^��̍yT��)'�˴�[yrݝ������AV����:��Q�x1���o��UV�_��TZ�뻾U�6�l���9�5�ףy�r�p��}*�hs	�g��ꒌ�Ҷa��m�{|�3��*2�6�� E;��="+! ��W�C�=��u�~�,U����!w�5��UBD��,�;8�ΙH��[s���V�2��vo�a��+�k�h߲��![�H-�1��Ch�V�A�'w���B�_��k/S�ү����D;��t����Psiy�K�+?��C8?mG��k`�įW	�]�J��Ej�11�g!RBC���N.�%�eA�V���b����wN����*�0 �܃�������@{W�x����WC_e�w����;�~�������>�E�S�C�Xkg }��)���X��<���1.����tV�#������'ɹ3��Z�McI�r��M)`pMO:jj����"�J���b}�ԑb��`��ō6
�x�9�����9���6�W%�M�!�����Q�:�۽2˨B�g^+a�u�;#ź=��X�	��B�9�X�**�j�6�ɉx=�k�֚��[i<~{��Z�����{Yu�3�;Sm5ݾ�P�n�D�/��Ccª��ِ]?�c�b2�Սo�\�,G�(��pɽ{u�sF��n�S�&(��3���i�-�f_�?ب*Y�qU�'w���:g5��ta��%q�v���^��^;��88�������C(�,�Ż�Ҙ�iyW��t������;%��Lj�Ug�a�p��^��m����ߒ��˃E+����Qb�87�2�M � �|Fn�Q�X�\�lۙB���X�l��(�øu�k~	�A����[B�/�Yfiq��X����Ʌd�;��o۩+Öy`>F]���vX��m���N��=�2A���o_[+�_��!)��G6P^\�g�*]�EDN郂Ho�@��@w��Ug�h(�?��~�����;�?t�q����� ��#���{��D��vvDE�"܄�Ob���W�6��w�`��4�1��H*'�6H�/R<y��ƗT �ݳ��<���U4�V�~J��C-GN(���W��mD?��5��5-����-�Oz��H�� ����}d�#��	�_����	{(�����l��ɺ���@4P��~���7��"):0at�@��`�Q�WS��u�˕��Y���;����*�oئ������s��#�gI���F��U�%�=I�j�VT��5��v�I�50
J�҅�A8�J���ç�Q���n��$
�(Rץw�/����CQh����GK��s�"������)�z�����3�0�y�H�J�d��"��Q�F�E�����iI��&����R��C�O�冫Kҳ�l��x�1��Ͳ��V��E�8N�?�`���l)6�'�W�c�f�7gB�D��ق��'�5�jg'a���Ȗh��)Q�GQ���Nz�3�`�%�"�p�x�*j�l��lEa@���6�0�&2C�����-iȣ��(<=�3��JV�'���<-�J/voZ���%%�Z�����E�*A5W!��[��b�Օx=� 0A?��⒁�醻J��(��u.+%Q�MjM�F&���+��CV�8��B�&���;��Sݍ�E���6-�p����-)j�Sc�]�x�r,�UV�y��!�H O戻K�M7&�st�F��i0����'F��8�h��.��+[��{�����!�W(,C_=�d�h�q�K_ ٣3aߊ��"X�XܸA�4�	�_(_8 �?%z��E7Be�1��U�/P\?�v3o	]�-�M����`��Uz5��g�,��(�H��-	R���C����G�6(�Y(���Ц�g����@���}�*u�iۖ­~�ڡ�d���\�8�͔����)���5���?�P:�;���X����D���:������.�J��'���
s_p X�z_մקۓ�색Wݻ�s�iV��"قt�Ħ��xN�:ۺ��Q�nγݘ��l��ob������4�ˤ�My�lx4��n��`F �|C��9��(�ΰ�c��.:!C*�j��R�ml���ARj���j�������e[�@��A���B��qE�ͧÁ�RnX�n���m����k�-5n`_�h6D]!9xiE��BN�Kj��=>�0��{u]�O�҅	��S�i(��x�a�q��(`	m�=n��U�	�\`�R���C5�%�t�(l���:4�d�=��d*���~Q a�JG4���Q��Y�l� sxQ��'9c�w�s�<�E���d�{5�#ESξj/0�s����&Kc�5�W���ڤ����ʓX�m��ġ�P�0��p#a|W��h0?-�g���<�q��1]^^���k~w�&��r��������!���&�*�"{�5z����ܴ���n�}�f8��<�j��.S�^z���2�Hy�!��sL���P����X�|{�ʝ�米��Vb����s����A�6���#�a�(25������WE�i/{tY�fh�=Y�.Ӹ�&*4����p�1A�z���tuGh��5}>啵��ח���$��[�Q'N9M��w%�*���E�@�j�{Mc�`�;Ïd��x�ăXs����F@�b�`�[��9�<� d�sAn�'!�����/�* S��A`C���p"�8��,DL \a���P�i|�n����ϲ�.	�mD�F��t���P;��/J�Tu���NA^��e�-�KG��ɟ�q�k´�Y�:�Dp�CMsi�u�����sē�4Q�%e�m���͔�E�ǭ�Z�@����}n�s�) %/ڍw�m	�������7p�����ZI��FÖ�Rz��%�6����\_�<l���t~$sߒӯ66\笖S�zm����Ȧ��(��ipXDMF�J"��%��,F���B�ou|6��eKp/��MA�y�l��T򼀫TmH�mŖ�?ȂZ���B|��F���6����X�ώzB���.�ۺ�\>��>>BZ���L.�E�<K}C�*o��.���q�Q�sk�w.�N�#�����#��D<�a��]��⢻X��-[y�t�S�"��'#�9_�!z�6�d_3C9 7���t?�SD�-��Q҃��;���1HL(;�P@Y�o1�����l��v�V���~h>�4�d@&s��!\��1HfS��%,�i2��r��"&�7Ñ�I������Kkv+j�;��Jg�m}�R 4q�P�u���3���ZE�<��1^�xVX��*K_
�X��k�T*e`;k[`����&+������#�e'�7��P����;G��n�%� η��h�B��5n�E�w;;m�16��}�h��>Za8A�I���bk�*�b#fG�̉𮀄�_'{��m��u6��X�}>�o��� ��́Ҟ�������"l�-�]�y'��
yf�x:n��Dm�y�E"�$���Nr[�����@c.%��79�KV�ĚzM��B�I�\w����l{�������!���6��Cp�^gn�T� �!����L���`l������|�-j������dŠ��V<O2����c	0á���Q�j�r�<7���}�Z���82BE�F4��0H�`��Q) �0�������P���Y�<S,��'�����?��?����4�c� ��4�]m�jI�Juzj�!�f���J�b��k_����ߘ���S �?���*e��i�+�D,�@�2u�Z�&�v��5�����(O`C�J�c�K�P? �o��R+����/�5'�\���~mCc����;W>���T��_�W�'F��k9�V<�R��q��"QXQzеwRcA�lP�aԑ�)��v*�hft�B����8Ue�u�T�N'����!�MI���Ӡӡ�h�4�"k����8^t�ԮZU�ٖLf&�<C?�97���a|��`rX�wn�2���FW��5�^Y>�	>��K�N�ˬ�׷3ފw�Rv�l�~�^0m\��F���T��]��ɘ/�CԺ��m|&�BH��%�cx�hʿ~�K��6:䰯٤QQ^�f#ck�����g
E��,a��j�I����.�w� l���k��V4v�=S���F�t�4�ro
�V�e0<vJ 7����f)*�O�n��:���r���Ɛ5D؞��껶'9t{́�i}Ҙ �lȱ{T6\�҄jX�5�h��������7O�Ѻ�
����+j���gA�?�8�ߡw��6� M}z9wr�ĸ͡�E�C��R��	��Q��u���;�u���gh�8�)s��\h��z V>�AVDׄ�� #��9�!��uxs|����
��M�:�=KZTe ����JR�ҫ�7��`���>L���b�p��$�!$ ͷ�TM5ݡ�a��܎]�gW�"�q��f<��&w��L��6��!�]��󁓆�ͯQ�j�����M�/�2�Y�yd`*�aa�c����=�M�~����>C����v�������o�j�Zso�|_�ןPí�]1�ͥI�:�y�}̝#���R�8����S��/�yek&��T1l=���;R�K�:x��sD��O&q�(�1� ���G����:~"�#/�;Df����s�5�ZOW �K�ah��}�0�}� �?t��Q�}E���M��Tj��r��t�Awq�2^�_RS1��r7����X�o�w�o�7C��p����d�˝IZ�冏$]�{��\�ɣnb�w�l��J�$ qD�s=z���K�J[����ڹ:�i�+jcJ(����f�q�]�@�"��#�̦�5�����4�%}�b-�3;v�E1�P�p	^�|�ݐ̕B��!%�쫇�[�D����_��2%R�vNH=�L�`��xLl cSL~�p͡�x�MU��%�'{C)7_$aq��/@]�Ѝ��p�K�i)X�����DfD?�A{15��Whl�r�{����L�g˼S;.(�/!��2wc�,�`%����͟�>��N2/�CFX��h�E,��q��FrK���l��~q����U=r� <Wj�?��ԙe�Z;�%-�<z���� ��k��ִq��� 9�����۾|Tzbq�K*�������h��'>��Ji�}b�!�a � 	B?%���>W}�nħ��f���h&�h��})�p0_���̖'�Wz�R�(��ÐU��q��p*���	9�![k�3R��L�"ۭ*�<i�8Ʈl��8f�1!��eæ��M��C���}8�o@�t�C g����P�ۨx}������C�BC�.���U�k
d�'}�c��������<���x��l��9O�����p�0"��q� ~M�=T����4-�G!��������(V��+�"�۷O_���X�$B�ɔ�!a�����u����8�/��'�A�(C�<q�[z@N�і��sW�T�U[�:x|gq�a)dh2�6��ه58����M��}X~�?/��zk�\�1���%����y�j�_��)P���U������' o��3T|��E%�7��)m}�$��2xr�h��t�+�h�&5W��%A�3�<@���a�C�)gv�Z���"?%N*�㔈Ef����[!��J�����[XG�1�(���,�c���L��ȈVJ�f��pE0!z�"uI!�3:��n�Jh+����:8-�<�N\,��Hʌ��L�o�Z��LֶdЍ�.�T����^O����ox�\��H\B������`8xfcAfkF�ز�Lf���Nv�����$��,��,#z�I�M���K���0���k�j���m�%���ߊ�$\ހ,v�D=�I%)!�J G-=O8y�DOQ�6,hO��j-ާ��%�9�=����BI�.�)�� �Q�M���dE�gE=�1�ɵ;΍P1, o�d)5���Q��#[�l�9۔E�#���t�Fo�۫�E���✔O����l�wa+ǩt[����*��m؎�c�bخ/X�{FV�U�[��@�J\N
���K_����,뉾�V�i���kM�3�"F)�����W�������$�����F�Ҿ6�zR�Q��5�y�dv	����H�<d�,��r��-�F�mJdyi�z�
�R6d��_,�����
)����Z�%Я��dXھ��Dtl5�`V��D���@�a�y.�yՖ��s���D\���s�nS�hI�]������T�����sߗ��-��_���<��s�H��_��v���K�r&0���y���%K�㫷����о�� ��ou`��HP��#Cg����=����0{N�r0Un��7��ӂ��,�O��E�&q;+&0�3C �=UKXKZi�yԊ��{9G5{){���	���+2w��Z�x��	�92>m��X�-$К�W���yt���B��s^ ��&E��#�!���M&;��EH�����1�"�^n������Ne��m�yyH����6��s�oO3#���嵍����8���8���l!��|�L��-]�K��"�%�I�VJ��<v���!3�`�\(Ş�P�u[�t3팕8�-�7�]F���6n]��] ~�Z3��E0D�'˶����o�Yl:� ��4ذD? 0�:�h��f�x"������S��Yph��:�'$?R3�$.s���D��k�{���^��q[����QC�������F�2�5N�Jt�w� U�/A\C�d���kL��,�U^�G��C"(nS{r�D`u<Hk��G���Ee1R��$�S�G*��M����J��"7E;e5^Ѯ�d�xܿ��J��p6�� �]�	D���=���*6S�V�����x�,�#֒��z>p�p������N���Kb���c}D����\C�ɥ�QB~K���+sN�:�xn�?�[��{CnHs沔��'�P��g����g[s2�b(����6 ¨�c���<l�I+��ߑԴ�0N[���P�]6��ct�1��#�@������B}����-"�ݵk�u����`��C��w뱥^jy�/��O��8�%�QB�9��˽�܄R�&�M��oO�hS�����sy��ɘ���>��Y�J�?�������n�y�P"$�$k{��]������(��B��#֯t� 	 �/�b�Y������\)+}J����.����� E挧��jg�z�%oy�J�O��%��VŌ�(&���������{P��ʣ�<���2�G �u^O��ӗu��́M��~���\E��Dצ�D��
�E��8	�YGd�3�U:�%���6S����ͨ0u��Q�ܛ��=�N���_ƪ"e-N�%9����[[ޚ_V�:ʋ�}�]�Ko����cn�7ZI��fKWf�U�>"p�.� �^#��M+N�������ʨ������@����v�G��[f��f�ߠ߇G�q!zh'��ѫM�����&����쮎M�S�4#ޙ�G��y���tc7"�3�
���ͣ �nr�� �qkҥ�P�x;sK����t�0TT��>��n���-֎KQ!o�>R�;Ye�f�L?DD�(\i;i�O�7j3$_�I	?J"��-��!�U8}4ǆ�4,磂�?oHȚnVuq/�d���5d��2�Pu=Wߐ,��U{���};��jG��9��[=�o�FȔs��=H?{ ���]�N�+�5�˿~���)�E�=%yaF�Q�/,��'�Q��j������_�!p�,3C��E���$��hp�h�7���Ǆ|0W�a��ݥ���|X<�π��*����MC�X�'�r^����~!���>1��	O�������v��j3���9��R&� ����9����D�᫨J��qbZ�π
��H�'��݄����K�!��!���~7���`�t��:	_�2b�^Wd��\2D�Cн�haP�1�]A݃ui˝�]�_�)Mq�Tդ$���L_g%��9�o�^�@��J?da}gց�])=��vD���Q�>?rA��|�&ܓĄOA���/)�zR-Aaז5�<��`��MFav1[pP����Op�)���"RUx����*�)48�o�H����=u`o�P��}�3$�k��R�5���~��5ɐ�#�%$ޥ{+b�W����'�����cT�i�t��	���+d�;=`��6��`Q�����B�m�I��oǶNʘ�z���D"~=¿���v�M�fU�NS�����+��PU�;���zx�ґz<��z�m�S�ڤ���5�$�2.�]Ύ\�G��f<(X�b�R(���8��%�u��49tӱ\7��~UM�����z�j>�Ȃw��=����ѓh"�]�b�}OJ1�'5�o&U� ��$���A2e�kH�ފO�ҭCb��`7�z>���g�l������9�s�p����o��5�L8��_\�s ��%�&-.��3���DĺO��}	�;H��R���m]p�n@�[cf�і� a@�'�*��&����tzz���<Ys6ϟ�Y���_�ߍ"�,��|���Ve�B��s�ݐ���BN ����`{N2��q���� g�M;�ЧH'�N�P����o����������jN~z��d�{��8��31����r�����-��5��9/��p���� ���DIb��/�{�ǡ$�@%�ƾ���Q��^�[=���ǌ��{���V�U0��O|��
G����p����2�
�C,M��s�wN$5:%Ip�	��Z���%�9�\	��w�����c[�� _]8��K<<�����1���t^/�#�3�h��xp��7�~΀����m�	�'C�[�5
��V���=~]�I�Y� ��C�o��RgՉ�u6wV)��31�c�,"Ϫ��= {�Zgp$�y)<�&W��#ֽ��d�}p��K��Qb}n��q���)�r���Y� ����Uפ8�+��kIk��u[���}lK� i���hdQuy��{�C� ^�������KS{����Ԏ��}�É�+�z�� �9%�@B�/Nrxb���D�r�j�7D.�|�%���#l�g��¦��v�)�v��3b���<gQp�H���k�K�)�����X �Loe����eF�4!s�?�n��:��w(J0��'���BA�#B����c��l�]w�����p���Jc�u�xn���<u��3�њ�2���چ<���(ۯ���d?��1����_��_V���L�`���@�T��h��p�e�FS���r-q��} �L�Y��=U�B8)M�x9������J�^#ݖ��[TK�Y��ԯ���ib��w�5���[���%�xO���,'�D�x�Q���;B��\w�uz'<R1T��a�	ƪa,��M�9�B��s��Nz��A�B�����jG
aO[��6�A���Z�~���L�F~�N�Zɫ���p<ק��š���//q���d����6������f����� %�c�;*mg(��7]��֠���}�b��y��ʓi�QzPFk<E%�-�}eP��iE�x�~������Z�3�+}Q��(�>��4�u���{�xK �f?y�Z�`�J��g�3��0�em�o�x��ʓ��f�[�;�9����)�^��wO8�����`����%y<]��E��Uޑ�{�u���XRu��.�*,�0� +uS��P�p
��X;�}���i�;Gb�\G��<Pr�=qu��b��V����Y�a�}]Z=��E]�廘�5&����W\�����U"���87k��?�^�\�կz�r���d�fc���z�.$�����5-��jk2�Th�8˽��L�'=���䬸0�D�8v�j`2�O�%�M��dJ7L?�y�<�+6_�˩d3W�ۜm��SJ��EBt[��:��]ī�:y�΍W��W�{�~W�|���J#7��(�_��Q�Y8����攸�]e�� k�$�$TÓ'�u��Y=s>=�K6�$��S���?�����sǺ�X��L��܇r��%�WV�������]h��K%���Z�� H�*�b����G�I.n�PY�7��;i�6����١��*堄����nR/����<��|]�A)�&2`�>�sf��K3��o���69�}��v��B0)��ΐ�u���.�&����JRK�v�5؈����� ~!��fgJ���DC�͍�����P��,p�/����A��� AOn��A~r�0��`��b�!B)�~{�}�W��X1p:�P�Lk�2Rw_#��B��8����>6�ãl��H�� q�����VE��omN��V��V	�o���q	��'Y$y��ܙ��.4~�A! �C�/7Cq���.�{촴Fu�oCs��ShY��%��nq�e��1w�XM�,0�߂!-�h#��Y[cUa�cLǗo�� �ZJ�� �k�Tꓵ	����P.F�ɐՑ.�j�@�����xw�5k+Q�6�Y;��e�z�����7D�@��"�v��Hԭ��'�oA�AF�Z�X�C<�gt��p���Xs�Ν��5��dʕQ���x�����Q�F�#��G�V}���Tܝ�uY1Ĵ'�N�;`�b��G�Ti�p���u')��*�U�v;��ڳ��E@:�Y������@W{�u��"%�S%:��01֪�e��L�}H٬�+ i;�x�t�F=��%Wy��:4c)��$ j�f��nႽͱ��K�S��!sR�ܟ�/��Jq����vm�X��ɲ$�G���4�ؿ��W�G��.�_�ڒ�E�53`��yvqı+�E��d���`y�v�3Ùȭb�`��]��;!��^~`&h6�	�į�ỿL?���,�Lo�~��ّt��ʌ�a�P�j`�ji��3�GH�1*�T��٬梯-�	��j��wI����E���zpSK���8��wq���R��R�RMTǩ��Y�Vm;�)2͆yo��ϱ$��Ao9��@{�EY��n^i'�/�������"B�F.���&����Q��<�nvO��G��~qFL����X�%b2R㧙���<,���Ko����]��^'ے.2RǏn#��eE�W�q_�y�����i���-��x�z�É,�m�kO�LÉ�k�x�#� �
��܀F?\��D	�ܪ6X���V��ީ�Q��5Q�O�VC\N���I3��-�sUsT���K��\H�æU�ԩ�3��.X�-k1>�]X&[�hՍ�B��A��?�a����U���I�w�/�O(_8�&��BW���Eh��sZ��F+7�Az%~S~ݱ����(h`�l(��Sp�É�A5�ZJ	8�<0(q$ �-00���e�$�5�%������=	�4�^]������(� 6��qek�
��m�қ��n�K�� �Of�(��b>����H<�*!2G
]<��"#�����jNb�L��G�������b �k'q��^N2�jZ�zR���z�GP�w�mA�\�0�4�2�>u7@HW�S�{L��6�7R�a��K �ݰ�K�����������1K�|c����r��W{#;�/��]�*��	%"E��� ⥆�PV��˷�*���g��u��v��	DA��;����@��8�|���z=b ��o���E�o�3}���h��N��)\�Ql��VZ�S8ֲX}�T�W�G8�����?=>ː�L�Z_@VSs
�9m��$'a�B�m�6����|�c�4�1P�`�����P1�?�C;�B�N@���	���$H���ʵ@��e�o��l(1I�8:����:��T[�	����=|tO������d���F;*x	��9�
��%It���\\������w�x~�6���4�
��8"�*(��7ӎ��"{�N�z��bs��� EY �DGUk\�ƯzQ�l�0�� =Ei��$<ӭ�/J���ct�G��T;]���ޚ��s����\��߇s��nqo��x/��C)�^�`��i�O_,�����`~V��Qq�Ή�,�͊>j��e3|��.��� 	A�m9E��=Z�g3;7�LI �5^v����}{�T3�!�q��D�#/Ļ"-l\�&�񐎦0���w�5}�1Pe��$dk�[:�Ml��5lʔ�2�5P,�y�8K���g��/j���Y^����9^�u5©���hk*J@� �
���ڕ��$]��+�ѮG[� ~�ߚ[����,@��#VO�.L$��2��O�=5��exE���6��	����<!�Yux[ H�m�FX͏EF|�������%(`[;b96��+ņ��bV��t�f��c��9)q�ٺ��9xIb�	�L0��G�+(�ȿ��G���rFM��D4뽘�!:�:��Ƃhϓ�z�l��G��`�Ӡ��Ж`�]�F�é�⧲gI5Z����.���p��������ȗ\T��Ⓗ�)4-=;]Z����ģ=��/����,�5g������t	������6����^��~��w`��vR���[���3���rȵj���bĖ��
��/Wl� �š�R�T���A�������Fd�3���$E��|2���$k�S�G�qP:�tC�����v��_��'7�B��7;�`}���� �mLd	`��M.���u��J��W�s�����_��*�_}���0��E��zVO7ۥ/V�Wiqn� ������_�Fõ�M̦^I���ɟ%�s#��L:L�|�H��a"�h���;���!������-eu*ͿPإG�f�!������aDv�=�vN�������կ�-�J^]Q�!z�+�͹��H���f�n^� Oy6�w�
"{��CG� ��n�W�ۋ�&�o�z���7$C���E��\=�@Ŵ~Y{��'1�������
�kl�|�vn�,e��٨N-�g��h:}#.,��?6�������&-Z�f#K���2�a��i�h�c�P�D?�>���+��$ \�!g2��tN�|�7��E��lb�9�z�V_�x�p�oaq����^�g��]⾺M�Kg�v��-�J��ލ��v�{�s��(��K>X�K��f,@���c�l?��7����yd��i����P[�!����_��bM]��ƌaxX|�w���a�`b��:�B����@�9��¯���r5�S ���Y��QY�����A��l��8�ܾ�q��z%S��Z�9����2^�q�e=Ě�C���PY!����.:����<�h�bI-2��x�j}pW��<�
_�(w�D��;�*S����e�������i�w�<R^l;�3��?=YϨ}��2����q�!��>�Ft�˿�7�3�2�!�гƺ�},溱l��Xy�ȸ�+B�SJ�Å�~Eb)c�9�5Ǣ�D���Q���ρ����ɐ$��!�����Փy/A�L�5��s�P]��G�8�+��Z��]�ޅ���N��)�]�¥ݟ�����Y��Bs\ml)�+ԇw�����t���.�t����MU��ׂ֫�~U�3(]��X�=!JyO���w�;`�V�y�ñ�~��YL��=�A�Ɗ+�ur�0ۿj��ic�q��-���p�����d�뒔��1���W�r(�e-�V(}��pu$�J�U�M�<"@{B�k� n9mn��O
�k4)�9�umVE���'[C��i\�|�N�:����p����rX�|'�����T��pׅ��ٖ�Y0l��d!��'���ul?������hd��H�D��B��z
��3��j�7O���3����Nܩ&{�ܟ�?�?yfgN����c�����\���a��Wnab�f����-
�e?���w�F�ϼ��P�AW���䵿�?�+[PJ�����ɥ�_���p�b�Fr���lST����xJ�r�t���XII[�3�|��L�mP���y<�a���C��Yn������(e�pxvO��$���$Z��+��`r��熝�<��P�RL{7$�W���`d��]��i����a��O[�!�dI̯���@Z�����]����p%ޞ�����N���!�){�=�# �J�s\�<W�-��ߞ��|�eoܐ�*��Xn��a��j�ϒM5�*ws��Y.��=��Bd@�����/E�?�de�th� q��6~'��[s5�q�(�t�I�s�T�tA�x�G��/��)Z�r��+Z~��&�ت�,��5.����ܩ)ߒ�h����U�'^WKsW�}�O_Akii�4��R p��j��n
�Ĵ�X�N�w�+N��q�a��86�"��"�+�����,�kL<P#۫��݁V�L�����$nusWz�H�\h}C�^i����׿�EF�us�<ݬf��@�,1�c:���v�G*���<��9)RMᬃ�@���a"���l�6e�n+���8��o�%�ֹ�Xq0��DLJ�(�����p�o�N��^T����r	B�H�B��&FuU& ��4�ٮ���)��(���Y)xt	5�mQY�'����br9r�%��e���V�1�* �}�N�t��)�c��Y!S�V�Hu���D�݁��)��B4�7���8K���+eUĭd�O��JK��/�OP�D�3������ː�Oʳ���d��}*$��Mc��u���~u�c�7�Y������/-���y�>�#Xx�n��Z�Sj�e�2;��I(�9J����!֔��)��E�k�zf�&YG��C���,�:���}k���3���K��݉3~�Q<�!/�Iي(��WG��g�4�r�Fk�+�b�1�m�f�G�� s�W��jr��<}k� �#.�Ԁ�4a��`[�oyŎv�0B��Z2�h9�3��!���Ec�Y���Tyܪ�<m�ͺ}t���"S�9�N�6R�yS��RuԈ���2�����:/h�����$�19 C	�1���W�+�>�����o; ��R
ƕ��2>]����h@!�
��u�a�*���\=�Ш�Ε�:6������� �0�0HR��f��$-��p~N��ݴ�����eyZ`	M?���F~=��%�����R�+����(Dc�%��}�n{� �в�<�܉�e���§Wր/�7�Yܵ� 6E0��#��{��l�d�����Pճ*.���e�Q��A��a�������7LѠkU�7�繼��/F������b�k��[+?(�GG^�����_q���^�=����lg �?N�Y�|��"���O!�¹���β�Q\z�)�7�F{6�]qЬ|L*¥�66"1�> �r�*+X���3MĈW	[M+�s&�o�QL��z�~Y_R��=�nնo#���A�2����^�	.�KG�b�"{>	���ά㛣x[��M�+���@յ�'o����ۉT��_3�ij��CϦ$��(���"O�c`wӎW�Pc�|�C��YzS������i�dҮ&��tG���VN��k	>�?�Q/,�,P8S���Д�򵟾�hԡy�^J�-����'�H�r3��vwS;F>�;��b1��Y���H��lb���W��	:/��R(mʖ߃1|��
O�{��@��4 �!����5o4�kn��xJ���-�·�A��dY�o�/����@l5V9��@+%*kqQ��]����g;̠0�Zj�ʳT��
�N?lV���rӬŨ��[�_�n���⾨;q���Om㧘ؑ2u�SwMǉ#����-CΕ�A<Hs�){��������<�}���h(L=5%c#��k.?���9i!z��cݝ6k�]�Bqsv6K�� �T�����㗒nkC�0�/4�˅��uō��t�*��!k�� ՝M]=eC%��~�>�ժ�f"D���4�5��f~�XѪ���Ю}�f2h�H�5�	���,9͖}�o��)�� �h�e)mg�L�@���g�$�4`�S9�One�uw=���$�Bk�W?�#G����%=��\ȏޑ
�P;Y�����9���D h^�H� 4�7��^zF(���ji���'ʹ�C 9�^oI�̧2*̊���u�g`�9�	�*���
�?MXW�T�V�O�n5v�Nb������Z��j�FĄC�/V
��� ���K\̚M�e����c¿cO�M���w�v.��=����LC�m?M����(���;`Rrؖ��LCA�,�k��|G��Xʠ������w�+1�F\q_` ��|���h)*^��s/�T��>�k߷��Y�ο�������TEH8�tL�+��4�ˍ��<S��2��Uѥ��c(��0^�{@gu�8�5Ȭ@��]�g�\�0����a�>1w�,:��K��,�)(P��} �p(GRt�9c<MV?PSxE��!]�#�5蚓n8[��h�}�>�g^�\*�ϡ�ub�y���m�C�� I
�?k��5ǩ��"L��[7x��
�]�{���
��Z�?�2�b構�Z-�jzm��c��z�ݕm_�z�-ci:����ُ��UB���s��>1���>��b�U.LW�<�\��E��%e�$6'���Ko�t�h�]-��$�]VC�۩��D��#&L��W�\�jݩ#�M?��C�#�D�	������2U�����>���ex�gs@I�ʇ��$���Y�6R�)��1����Hd��EnL���Ų-y"F��[VL�ݧQwMq�m>���}�'ZY�)1w�]�������A���� [u�a"��b\�B"�`�~�[L���z:�X�Í�!���(bM��n��k!��?x�j�`�>Ja�l(cf'�Z�ĸ; ���S ���"�}3`�Ը�qXfgo����uN7��ٕ����Нt�r%=��Y��� ���h|憇o�E���w��HM���č6d�����hȞuo>�Peg�ӂ͗wn��%���>`����}��r<��~����M���L���}:wb�r��t���괃�@@�z���9�rX#���RB�|��[���B�)�:9=r򗱷.6&A�CP���@r�L"J�Z�&��)^~2_M���Hzދ���_}�F�>1�XO.#� Q$��b Ά�����T�X��!�P�g�ΊB�Iw	��_(����#���ZZ+���	��T��W��OXF���^F�<�eƃ+����3�N�tI�����t���G���$�F���X�dB��Z��gط�W�"4�.�nˤ,��]^?�I�/�7Iaܬ�QW��C���	֐����-���SG�t�2��a.�UKw76YB|�~�l��5�6�үW�_�aô�(Y�R�*>r�Ϙ����g�i2��c���ݺW�1$W�`�8��2!�#�E���Wܱ,I,� ��̿���1�9� |{��ߊQ�7���F��v~d�aZ=���ݜ\Ȝ+���>�����^	��.�_1������-���ѥ��-�觸$[p�����d���"p<�D��F��I�ӉaC����
T8��]����WV~�Td�s�v��'�����`�XFfqŚ�������4���^���MdK&�_��/wN&���%D�
�de�����O��Nܚk��#C���{^�B>�����I����;z�|R�_�i�p��V�U���6�~h�Ôdi�h��f�Ω����m� ��x6�`@7m�����]�&z'T v�X���
��!{����o/_Ge׺��3�����0��V�~(ڻ�Y�m��������(f�(B�������F5�W�,ݺ!;���U��
{E6}!�M��*Jmy��V�{t��mگ����6�@����ߟ�1����q8�����n�Q��ߴ 2]ţ�
��s�k��	6�7_��Iaj8Ey��*K�?ej��9�0=�CARa>���ͻ9m^"��f�j�.#��J�]eCy�6����ye�;���IsT��1�Y��ִ� �ܥ �I�*���(Z���4��E��mi��Oމ㑱���l��tn�s�y�H�A��j=��^��v���s���Z��:}'fHݭaP�H��K~W�n�8��"8+��� i�n�N�	���WE�r�/d;���m����?����9i�BQ[ͫ�����Gv�I9�.��� �sL,M�ׯ0�}��l��U�{.x�0dY9��"�X��2�"�)�Rî5��B#�zM�WJ�v�wx���X.6[��}�t�2`�8K���-cO(��%L��"1�Dj��w�hCQJ{1ce�W�.a�,}�����UGj��$.m0�k���?�{A��'�$�fG٨��x���Ͳ���ӎF ;ke�a��I��*�Sj?��h�"�v"2.��hbQUO6;(��m�gt
Gx��@B���gZ���U-]\���p��v7�_��?뇳0��[d`�n�3d��Ld���X�帿$�&aM%����;�!i�L"���E�:���O�D)k�9�8�ث�u�q��u,���\{l+�e���dsx���C״LH�E����.��e�cnK�<4��?�����;��t�82�����nZ�C�B��ٍ��jۮ�Q{)�:}��dR�Ց@\l���@����o ���X\J�����`�6�
�	@� I<ϲ��\(�}<��%��'�]P0��q��`���Q�P,Y�v���!�zY���T��i�Q������UQ$��7�^���O��R���]��%â����{�x��;	� �@ᷬ�ɓ69�����UA�<��;.ܫN1A4�������
­�6Ӄ"�:�	 �|��n5��(�
�z������#T �8Lb\�)�ZvNt���X-���砾M�)� 4H#�82����l�1f�Hs h��.���?{WMP^T�}��X��U4�BtT����6�h�D������������$5�"��٢��_��5v�h��2���D'M[T� |8TJDz�1�!�ߌǿ3f��g���m.$�|e�����R=c�-"���o��,�]f�&��V�u�>�u�K��?�P�AK��e��y<��H������"�]8���S,�˲3��tä�
���&/0J�4�6>����-���ez��0��V��o�/f�d��:N��F,x?ғF�X�$
���dM'_
�3�z�(��	��;�9<���2��A`0��?H��Ѱ�t�V-�V�].yp׍�s�ݺ9#�#�Q�M��-��VG��f���2���M�_���:Acރ��g
�X���*���rZO�����ѫK�x��2��f7�� ?��Cņ� L��M��d.�_�U�k� 虰w���G�(à��i�I�����V
�-�r��ֲ������lAD�[��d�(X>�(���.��}[��Ҡ!:�1-ئp��R.�Y��	���^
�PZ�W͓�g��:����à�$O�Ċ�E�=	�YR�KTcr�l�ri�����_;���f>���+:/G���:��vkЕKc�X�{."���	������_ٷW��D9Ctt����K��hd��-OI
�O4��Fh���3�ʨoX��T[�y0c`s���=���<�Ŝ���5���I$6�e�%�(��կl#1��\$��c<!J�y�c��àQ5�]y _=��n!+~�������>ϳ��`2�V����9��}9W	� Z�ȴ+�	�ٙk�6���^8E���3_e�G�=;�=��;���<�+׳:)�E 3����r����������SW;C�9Lj��oPiW��?�{�h�>t?H=�M'#��(�����������e�(`6I巔�{��¥Nq�{Ѹ�/V+���^Y���P�,�K<��z�T��*�cÿ��-N�ĵ)����Ȓ3}�^|�3���2�E�6�7n��E�t��H���Er��I!���/".�m߭:	���2���>p?@�,fM�Y�C���a�¼� >�;��*χZ����w[�t�˛��T:Ն�m"�dWL����.�ǀ�ny�(ؚ��A4�[V}G־<��������2��w�4�n��f�cc;���B!SUm�����8�8/���2�}��C�S9?�~0R�6��d�YE6��QZ�˭�q�Υ	n�MeM-��H�68���G3��&C�W�Ο�<Y� Ő�G<��nQzP����!Yt(�4� qKp�3j?\}#{�Ѽ��Dj$Pv����n�:��'���÷<ö��=�E��!G����NG��躻�pF���!©�Y1出��?�r��qŖ�]�D�`&l>ŗ��$�!{&t���� ���h������1�t�`������ k�+�����f�Y�ޱhZp��t�D�tq�x�cWr�r�8��Nas�W�"��c��.�pq:�A�5�#����BU�����R�#��.>����K���/��3�F��)I1�I�9���O��� ��Q:]�XQ˻VON�^�e�W�s��/��aIO"����oqE�C��v�a�F�ִ-!�ļ��,3�� ��ț��{�#�5ѭ�v�+��J�ǘ�k�1��l���_8jM�X�~A�e"��	^Q��j�s=o:�?n
�d+�R!��iA����fx�2l�� -$$�W/?-�.�ǽMޫ�q������1�(���l��=�2S&���L�f1�~��l�\C�N�ʱ��+0
�-J��^D�/�e�_� �l��g��2&����>�Ջ:<K���i)/��M�w�c�u�bw�3G��/�6ͩ�v͚�WcW�A�����.�<ѝε�'�υI)��;�j���/]��r�?ew��R��������N���W�}R8�Y�JqC���E#�O�ںS�0��-{�&��G
�*��Ϙ���J~�[�t������\n�VL�����oD͋_���Jr�ߨ����߿�Qn�k���R��ֹpY��t���o9:��j'��_��;tIU~}n��N=
�l6i�B₪�٨� l�Icqh���k�����J�����Ƣ�t̼گ�k'<���KxI.b]�oB�a��P��N8���%��U?�0�ì����bvLWk�;%��.��Q�?Ej��%�)�i1���GT��H=�O����d���NN��W�:%�-H�o@v�����#3����)����C�-;e������:x!~ �G�Yyɵ0�+�y7�����%��Zh� �ׯ
͚�V;����Łδh���B9LZ����c��,� ;����fcZ�5�7��;��17�y��� n�ᔍ�C��F��]�
�>ƛ�4rSw�p�T��[��+l{��k��c-쪟����$Bhpz8�
l���ٜ�����7����$�<d�)��~R�1?�엂P�q��,����)8����&���1q�[��Z��^��!*@4A�O�T���^D��^YM�P�/Cst�~���i�H����Y3�����w�˒���g���IUN���|�M�?#��^6�F6���)颃��4޼v�B��?E�s����q�	���(��R���.	\Z�G�{��Nh�`���� [��� ��)�fA?E���^�/y
�Wh�_����6�#~���yQ��/���cW7�A��`�Xj��%d�4�u����w6l(�<����[Ps3ޫ���j�o�����"ƍ�k9[�2�f���cv�5��:��7շ�
r����� t���t�=���;!7�/٣=lu�N�����pc����Ҹ�E�,~�ꋪI�?���l��;�EVTo��;e�$���ź�
s=��l~�/h�:��׀�n�_M2L�~_��D��5������ag���XK����_�D�4�\���
˓أ�4D�AN�F��A��	��]3#Jv�A��C���	m��ƿ�s�@F��#�%֏+��5����69�g����:w �V�|���W�t-�%[�A��,�h�a��R0�Shc��/Z���FV3$#0�-oҵSX��u�r�PjJvr�1���s����ٹ�I;�9�T���V����t�j�c�`���⦪�b_0s�4�ђa/���O=}�_�1|ϩ��:���P���� � �`�c� >��B��T��(;���~02����ka
���w���K���$N�'Ȼ�0z���<����v��|�, _�5�dp��iPcK@(B�b� ~7���R�S����z����N�`�7���DXQ��[�'���U�7"uV�^��bC_|\�����l�4#�4E�=h�-�yN���r����l��	/�$u)&IťAr.hE;Gvqie�伫(9�
�}>�`U!w-�p���j���5���Fa�i�����^���zV�n�G�����X�o�yG"��Ѵջ�}�h&��3��=/���P�8�`�}�&�n)�r�|ץ:�{	���	�-�+��RJ!^W�̀��y1��u�*����a�9)t�8�(G�17�����6CK���s���E��g��Թ��i�A�~�L�ug�,�h���U+A�Kwj�ǫ��IAjY��"��\zZt�'Qw��D3=�����&�
���t�8]��S���|K�;�{�+;"��3�^�>�O���\��x��`.��:����EK/K;K�*���.�~��'45�M8ג�\�]�x>�^-�E9*tc���&C0���E�W�N�SUY��N3{�xU&�+��V0+�uo9���s�8qI���B�x4�3	����͛�wyW	�%^5bPz��F{�݃���#y56��n��;�9QW$/�n"$6��S]+Zߒ�����l@;�K�8�e�@ �;/�e�W{�8C2� �6G�`w�h�'��>y4����m�~�>`a�[������a��E
R�W��_@,t�U-����1%�i�nv�DJK�=W�o�I�2A'�c�>���}��_��A���{��"���[m�@o�VQ����0.b�l�OQ���=}��xK�5Q�*!+ɣ�t�kO"+�"�/�7��u�~
9�Σ���gb�h0�x<]�J�@�.����k�x;�n,[R!���Y�ΐ����5J|��*g���v<0Tӟ�C7T�cu<$��� �ú�Ub�#���W�J��RflϷ$�k7�7�ׅ�C=u�
-j|��W�T�s��dV���L+��f0�.d���y�L����(�	��n�1�^CRw}��H'>1X�w��U��X ���m�	�<?���3v�?�M_"zLH��tA��ڑj��%��g��V�f��:E�D��$蜘�o������R`V�W9q�eo��m����g�rh�X���C�`u���!s�|&�;�<���Af�cL�n���}��%ʥ��(��^��)�0��b����dfu
|���K�ޙ,�I '̈q��ߑWsĪ��¢����i�ȼ1>�	�\C��1�D<��ݼfބ�� �c�����E���n�p2v&Uku}���H>��ڂ]�:�k�æc��Nn:J0߉��w�fxf�)z{_�2�g��rL�H?8��U݋�<��O�ὕ�9�:_��$}�Oqb��0�`�6/U�1tѠ�C�Q�r�?r*������v�"��=>s�K�c��?~�{$5��emr��[M���Ʃ���!W1Fn�e/�ˉ6�m����	1�LQD�c�-��ܓ�=�t�Z��A�&4v�;rM�A�:l�ƫ8݀�Z@�f���Y|����~�债w��!6����[���s�AA�}%)���X����dԛ��r��m���C��-8�3�6ތf�7ݾכs��3���� /�K2?�G.�/ro�6J�n��1�5J`� LK��~���H�0D��\OXB:�Ň�A X�yT�׸���M_s/��=��\ƎO������Vn8�_���:�+ʠ0�~�3���j�^���E��y
�:��Y.��5��i?��0��S��NNc�ԑV��Ag�kU���)?�U?��,��я�f1���:I8B�Y��w��H6����
:4�ߺ�{���([댅D�k�.�;�Zv��/�Y</�x��1N�������hR	^����2$��|%���[LL�o��9Y�p-�<��-�vV��[���<�$"����1�%�yzYs�`gC���e(�?�[K�Ғ���>%"�_�N>S�xBk$�N#�����T.�o�هo%�(�̐� ɡ�˄3��� ��|�f��C�6#�[[Q�{t���{;jB�1k$�5r�T�N)i ���ۤ�5��������;8!�<�h��mF�́�8��㾮���wlJ���U]���@�6+�@nk�+�/]�^�\7̚^R�Á�Pܸ3��7a��qj)�����o7������'D+�+�T�̀0ѤOӈc9��$h��/+��8�h,�6ӝ�ky�v�E};�v��Y�w�����Xb�V�gHյh��5�|M�Ru���'������8Ym�xd�b�!n��K�+��茁��$-�E����f��p��f^S�#�ҡA�^��V81�w�wuo��"l�?��6�3��yld2���;0R�}��(���gl�_r���
eV�>�~�W��~�gҗrʱ��O�\�"bK����l ��&sb�S�����������x��>6��ͷ:�@���r?`4q6���_�]f9���A���lM�Ss`�5"�b�y���T:�{�X�fG} sK�Cʒ�8Cg�/�<�v�5Ϛ<^ٓ���(�Wd�	먍��/a�d�p��r�*ySu�[�ŚF�Ъ>5�w��>"����R:�Dp���F����;vă���N�����i]��#��:�Ce�	3Ϯ�y���]߻����Y�L��)�	̩i
�q��k��d�i�1K���t�=������q]\�X��u��s�p"��@�����
S?��㠄��W��CҶ���e���7�b	3~�I��9�P��ZX�� ��L��+z��3oL7�����TQ.�?D����k�V~�],.�:%��h��������P�١��*�g@�������?�wM89���A8����5�3�FJֽѺۈY�k1hbM�H�`� ��졶���y=�v�[�&�e�?��e�6{�f�&���4Ǻ!�t��c_�c̗�:;�:�m�C�ˣ��M��^�F��IKȶ�H$�z{Q&K�"���`��,�����F57�����Lg	A�x�d���<�X��V�z����
���|�=��jNZ 91�@@��cQ�)-������s��k6�Sm��ۈ�i��aP��}S���b��a�� \�f�Qo� +�򓥲�r7Z�`K- ޵��4L�R�ul�!���J��)l�����;	k|�	����<�&�0��bw0<]�7pI�\a�N�5�����&xfP�)`NGy��K�n��f�ܴØ��'��N�Y��|=j�d�p� w�w�<�g
���W���[�2��\�6Cj�����ei�Lxd��-��fCG��`�������u�>�R*Ej_��*��?��E�2(g]�V�:��;�~�<q�j����,�;��P������7�0_��y_�N���@���T��	��N)G�y��AhA�d��LK��r�W��[z�d!�"Ӗ��Ab5d��=���1[[UU���κ1D�B`��tk˩dڿ"�:�5�ֱA��'c8!�R9�!�,!S��M���%��S��D>m^��F,���<*]f�}�n1J�����P��V��U�Mm��E�}��(bR�k������fk>)Y�cI��Eը�S��L�dJ\�B�-
m���P���MH��
�����	���|B�bj�JF��԰{���ʓ'"���1�f��;`Y�L�FJ�eH�1@ut�3z/�Yq�`��{#�2�MS4 ()y�&�O�-R�ז����^D�vp#�ai�V�:.԰,Z������C�%������ʥ"�hks�@����Y�����"�T�6/R��5�W�8o��_(@����Ĥʨ�j����jw�OT8�����-U�<�3�zF��A�͍ڔ"�0KJEC�p��(�V�_a����睱˚W4��$��].F��l�	����ה+B����\{pҘ�kX�)�%�����Za���Sm�`��R�V�O���d{�f^�qq�5�������u _.��6�6���W�8�/���;��Pφ]�DN���ص�C5�7����ne����"�X�v{�=qh��
��1���[��?��H4k�=o���D˶nc��0<=�چ7~� 2,�M�m e-��%r�S�c�w�!�r�PN��=7k���L�P���_l%7���'���hD��g[s��˧&�ne!���f?
� ��7�8,=��>m`�\��n �\��%�FP�3B�Rb �*��bDuѽ[�]�}��}���-S���;Cf-Z�E8W>���$��Q���C�{�Ǥm8��)�@w�Z����Z��b&c�M�����#�_/�&�n:N4�ˬ��t��)���Ɍ�`�u�ũ���;������<�\i/n_B	�Er~.�2�+�i"����)B'Y/~�H�7�2Mh�k179�������-o���9�H�����2��x���!8,�ͳ#c���m66`j4C)>������(E��4��n�V(�8ۋ��l���>JD����	�ے��FI�+�X#d�XR�!���9A \bJj�Y#��"�Ă�Yi*�+�7]J̰|��V��+p�E��S��J&�˕��ٻ���Z�EE�bq�c>Na�#�掠)rl6�˴�[Z�S��C�ظu�6l�u��Cx�G8^G�ۗ���jM���fE�`�+����X���o�I"ՓqA�zsڦA_$�=�g�,�(N6�e1L�6�G�K����/t
��w��o�J��+��0�w��*��l9�pW�+*�i3hU�My�)����W2u'��|��ǯq�7������jF�Y�o���aQ���;��تs_/>b�W3?T�<<��G�s�>���c��������V��f�h���`�������v7��_�R7;���N���^F�����~�%B���~/Z4�y��?��3_���y!&@���^��W�B:rC ��v�,�~��패�~�������c�%�.X��֘�V�I�� �eZ ��J���h�%�}I���Ѯ�)�3+2��,��!������ڍ4r�L�m��[8�5 x�!���a,<�s�cDVv�Eֶ}�pP����'ax�8pW��bcW��-f���2!DH�B�<B�s^�y�ˣX�p�@�|;z�$f�榗�xE*��\O`���/b��"Õ��"L	��T��v�����_�?c1��^��S��0�vO|
���o���8ve+�� Pz�qg�&R>��9u�5�XG/����3�����$��01A�K�^+�dnfh�+��
ƪx9�m��pY`L�j�h��)>�{4�˶�_/�M6lQ&fF�2�/��R������V˸Bd��٨�
}x��à��xsH5���aW�q���c<��K*z��B�>��prxI�	���.��L�td�Л�H�֒�������BeK�.�7)�gF���:Ł ��^�Y9�/Wo߿�_By����Z�Ӡ����#�F6{:�w��#ې����-j�N�)9����*|M�l@��[4)��D�P4I�jD���8S������CD�������zI8��>	wd�@��!���#�x�	H"�~���FO�����������xQp#���DA�:��ľ8�O��n�Cm\5�[�k,��s��U�̚x�اT�h�otN+Y��a'|V���E�I�'w7ZA����W��	�B�I���8$+'��rg��3at�M�s�z��B�Q�+�'w�ߪ�&~�xE��5P�q�dm(yo2��%�th.�j�rt�~����~3>�e�ET6�6�kM~��~J��rժ2�"�7ch�u0���
y��d���%OM>Ya�og8C;d�,k4!��zdo�3`�e	�������+g���{]]�g��)��#���k�"�u��r���*Xb&X�_���N���0H���/�1��O�ʽ�.a&�����[k���� Q��J�O�����<<ێ�Jy{����I@^��&3X�l�Q��Ԁ+�m\�<f�5�����*ʕs��,��X.P�w,���_��,ܺӁ��L�_ZvMa
�#5
���W*-f�_v��\��q<���ʦ��%c���	�"�F#����8��Q���=��]�-���:M����E���=��\�
�P�� n���XD�t�=�$�^j��( u[呈ͱ`s��01;�$��.Ħ?��A�Gԇ��V�=�����P��d��-F`p��)חi�ύ����Cz={殽����3��!bޓM䝡Gs���| \�O5���L�#���<G����8vCu�[!�,T��d���ȑ������A�*�A���f}�yt�23��}�@}��ݿ&st˖/��u���Y���s���ߕ�"�Ԕ%u����p�6�L
Ȇ��I(G��=���Ñ�氝0O@�F;�������e��1
"I
.�K�N����D1qF��(S��S�5�&D
��EDId�c�b����M�|@o����� E*َ�A�����\yA=>��!��� t㸒�|5�'6�����52掞!�)�נ�[yK����?`5��j�F�]'�U,����nqu��6�� ���Ttc�rF%�G��F����M�<#7����+3������/ޘ�i t��'ő�:�ƻ5��+��˙�"��̆���m�w7.�l0�xo�_� ��d�h_���;	�X�
FǂX�5��8�֊��e�7�r��H��#�[�br�#ΔB������@7i`�x���3�W�� �̪�.6i���Vh7���\�V�e�.�|���2�-�\��?�jB�X����@'�׀8�������R%�Cɸ�b�!]&��b�x-����$<�?�����#� ���t�$v��îRX��rZO>`kqK2Y\�nN��_X&�6���*e�L�k@�g�@�!��3���}�G9e����!tT�>TwcCo澂��:P6P���ޅV�A�G3�޶,R/�o�.�a=������m���)�)Õ��w�<�a�-K��f�|	����[���O�QI���R�d����I6�M�1�)K�hY՟�2FA�A[�V�k�?c��k�I�"	i ae~�WI����D�#�\;/�6�»aEs�u�\��!k���io�c�0�ٔ)Ć�S7�lAYi�v�����E����.`*�-��h2'�"Ҙ�!--�Ռ�� ��Hm�;�-Aj����R)���(�����4��a�Sw�또.��/�&��yz�����Oj�5ϙ��rާ����������w��8 $��iZ#7>FO�kÐ�	�M���;��c4�K�ӵ%[�.T(�T���t�����<w�����P���S��_���W�C���:�"�V0��M�;܊��i�"Oy��,��5<> o���kߞ��\�e�=��PU6���w�P��rY���+w^����ZY�Fn	�$�;XfYBa��(*���L*|�A,�O*.��Fmr�G�K.�Nv/M�B{�ý}�[WX:X��Ч�����gĆ���h��*�B�������x��*G���G_~�]�?�-���D�f%~�w�:���XfE���E���޻2����<h��z���6��QG�m���������*��و�ta j��&Hd��F]XB��Ic33p
�u��ڗ+z3/z-\ ��@�%dz5(Ko�B���X��i=��FN|&�'��㌣�6ZX��G�@$�p���̝�b/Pg��8��4X�ć�-�=jl��1�V����z�xE1��h!�/_	 ��l��KtR]� �D�àտ�Jz%�R֧�Xj��J%��O���@p$��_�(�JƔ��Dp���@����z���b��gB	�-�� a��$�<U�=ٵ\�x���z��^A��ta����D������v?�%���{oHw-���O/1��C�1�5�2��_����9u�o\�]m��A��0�H�wa�u���U�� )n��?*'����C�zF\u�7TJڷ����|*�Ň��R��^��P��#+�V�qV@
� � ��R���GD�z.1>�����)�(7P��L`~`���P�Ǉ:I:G�h�h���G����I��!���!��T�6
�C�B��E���ƸT"c���m����j�҇����.�btS�.0wH�6m�����@9���_�$E�8|퇂wo=�RuX5���MR�#����3�
�����nS�sd��u�
؆�� {�U(݅� �����Q�V��˒�;/0x��Ǣ����,�ר�B�	ރП�}h�pźR�X��o8��6
��\'\�!��Hs܄L��b�^�+�?��E�!}%�Z� o_�rƾ|��%���{e�J_}��!�*9�`��J���<��ʓM��m6�-�`XzkR>�zj�0eySa�k�  �)s�:(�Tzy��ώ� ��@%[ݷ�~����z&��}ΪhM$�/��	�L�-��~�uY�����9ywfN�K�ə�]=PP���o�Qu���$�x{o�SlE?-���<k��0�!�a�t� �M��*~+-�v����j�
�P��0y��!�S�ȸ��[;�M���́e��w�ީ�p�A�S��ל2?&}=~<�〞���=�w���F�8�����=k��ో���}��ʌ��*����ߔ�s�HÃA�V��W)]k��)~�E�������&�%���yRFt�}�۸4�H�Z��t�O�J��A)�,�!2E���J�l?��a�)������a��{_�LYJ@�.��%�W�Т�K��H?fuʕ���zS��N� G�ܠ6u�p]x���+*����[3��+���X"bv��Ē��9_�����Q���w��ͯ�4���J ߠ#�wM�ah�}K.����~x��)V3�qGd�u�%�'~76P���!�A��u�j/4��V��^L�S�[��V<$�~�����;��BwD}����$�RMCd�T�d���W���4׊o<��O:���]�E�c4���Z/X�NW�aq*�s�xݴ�Kh�\�ڪ�L��q|F�Qw=�".�VR�j��>���P D� � ,�y9�a:h��HqJ����0�A3q��/b����I�B�'�
��i�7PSi�m?�:#\08v�  ���I��҆
�+�	�H�i_��mm���h��f�w��^fg��<��fl5]8�ZT�Z�%��J��	��K���6Fw�u ���f��^�;�؁r����������Lޢ]dͦ�=Mc%�ZH������J�c�f�8����Fǀ����!��n{6��A�l�����x�%��LFS�Y�5c�I��9�7�J���W-���-��:�j���{.\
*.,<�]�M�A�rF�n�#5�"�=g%T6�g�"����\2�~�T��T�������^�Y炬�6������
1�w�8L�������#g�<��j��F�(����4���so�z�{Z�$I�y[�1N��G*��}R�U`�,��/��͘v����80������7����5=�Kcw�<q���[$��"��y[̿T#��_�����R.8� �0oLe.��:�UX'�3D��o�V-9�T�?�J���=���`�|�M�R	\YaB�!M�,:3뜶�Uޏsͺ�#M&�����Vt!����.ͽ�3���{lFX���3?>"EM�K��r~J���a�'�["���qXbi��I�\�n�(N�:�ӓ��$�<����B1¿W�r����BC�����'$���匼s�Q<�r�S��/���mM�s��q;�u��J��L�3�����Xs@g��%Dpmp�D]�~�(�RĤ��e"�l+���4�e4$������!�������R=�R}���o�<N>��cR��UO��`�a�%��dy�8��"�uҐ�vw���6f���m���Ц��	/<�ja�� P���T�����! �jw�g��?q�(RI\�Ic���u�m�E&�ff[�q&�{-���W)�H�E��|��#��l]9�r,���ȷ��@gd�J 1�yJzt	���j��_KF07h�%Q�"B���O��Ă����1�N J9b���8�jq
���DBt�n���.
�*F��1r��Kp ����:�*RTVO����d�D������n2p��r� �e������|Kv�4=���ut5�b��cK��e�Ÿc㉎o���T���� �=`7�'�C�Ny��Sr�A��"�Q
ie���9� Ͳ�;��?����f�J��:�u��.WO�f��m�`_���l+�R挢H�F:�{>Tj�a,���&���a�&1[�s��H\�UOz���!-t��|���(���m�[=�&s9�C~QT��eK�����}����M�+%�m�"2y�����h��r��Oo:���s�0�qXvbnDabE�Gh1U-i�͔t�X\,eǚ����ۃ���y��x�֎�[�ib��3�`�;T-�qNѩ�W �nI�:|A0(K��w����������$:*H@'�(�lF�w�Q%�1� !�Ԥ���W�?� tMaI!>���#6���_g�)�P@��U�.��r��U4��:���E,-�Ǹ�����;�`��f�\�s6�u��'�zC�q����7�~�$���{�)=I���8������,g{���\;�=��������݆�;���m��I�s����^n��lQ��2�d�Zţ�龑桂�PR�G��RX�M�p�b���[���]�<�RG�U�?�>P��o�x�m�u���RRgu�XN�X.Q��rͰ�0�����Iù�O:~@Y���r���z?C�ܜE���K�=T0��y`��+2�=�0�,yF�:���3�F�Z�;�,Ic��I��Ў�m(����K��Z����4a�5+����*�?7wO�u,���.5���l�sMH�'u���:+�9�%�A/8b�F˷KN~��RX,��!Շ��|l�{��
"+0<1��:�Ab@{I]Tp$ZYVׇuW��DY���_��=����������z�w1��M���}���L6��a1m�k��S;�%��䤐�EA�����	�Ѫ���|��3��a]�f�5�7ڜ.�?I�p�"� A4�϶�.X�9���pwkʸ]_�ą���g����^^B�M��udoQ�uwJa4s�,����kI��췝P])��&�!ncyx���o�E���ҵ��j��	sKIB�y��������nuƈ��uM���A���"���\���I=���:�t\�t����E����r�h4���LW�y�3T����`�l#�_�4n�S�³t6����G[qW������Ə�|pD�JE�?a�j!���ub�yKT��b�%
�G��+�x�)iWxe��s�l.�k5j �w��g�0�0�\w=�Q�]c�����ah��n/?ӣ2!Cŝ&�̹�FD_s�g�p��h.ra?v���fjB��(C�wC�y,�֑3��P���:!?��V���ܸ*n�K-�~�3SYu:aP)��I�"�u����y{�[�,��ߝ�cR��K�{?�
��- ���s�k̈́�z�!����Q�oF�Y�>l�~�;u�+�u��d$�jhpnÿq,�5�*���ϻi�?lh�$�{ɬ����)=�GG�}&�r�P��S9��>pa�i��@y���K�<�_cP�k秆H�VL�t�	뵵�ͪ�A�҄���U(Ҽ��N)odŋ���-��Q|�U:(�!�3H�;c}�&??��a@�ۈU�d/����R������>G���,�� ����pϑ�@�!x^DG
�`ϘM?�������vF��Sv-��	�l^ٲ��~�9�.[�(s��"�t�nq9$N7��
Qhߦ�Lw��;=���
a��oٿS|��oE�Y����6	
z仐6�a� ���l%��P@��N�%�|��xx�P�7�)rg'�i��	@c6ۆ�*6����WK��������w���j�j����߷8��Z_�B%����O���dN�ĕ
�v!���HI�:}�/�[6���h��^M�j�E��Ԛ^�7=ݰ1���Á��bZ��,S6k��n�J�:��=<(I�U�d��6����L���V_��Ix�f�4a*�t�����-7SMe���O��:΋�X�Q�:c�%d���|eg�j�j�^J�ݳ��<c��\?UjSF���ED�e��G�R{�@݊�sX���e�qFӥ��6CP�>y�uYl= W�3���C��RgU��.�j�hG3�KdR�L�O�q�N��jb� 0	�-�r�>��G�"$���RKu��DR��a�l[0�׻�]L��)�UH����ٶ)���1^�k�	4�X2���6��+�-l1�U�<w;�m��W}�0뤬���Y�R��+	��D߻���Mi/��RKmڱ)���Q��kc5UM�߉P�V��kr�e}��04�1���Í��9��\�B��0��a֥Ss?��zQ�h�G����Zٸ��n�(S��&)6V�͒h�|�P�	䬄A܉H|D��� � H�>�n��p�k���T"�B����#[0$`���Ϫ�L�g�
���W�"W��w��Yɲ��:��>�p���:'�,�f:��sh�����'�ə;YG}� C\H���
	�֧K���S[S�G�
S  �غ]��b���㣉��-��~������Xז1�vH�;��$A8�����Y�P����W��z�Lv\����L��f@h%Pޗ�-�K����*��:\nAv/� +:�VIclt���b�<�� �v�Xr�L�֢w_[2�ȸ5D�C������CQ����s�Xu�f!]��Ư��%���pB�����S��|�z���C˶4�<������Q�.+��*�b�f f� �L�?p�����!ڳ�pa5�9t���Z&�(Q�uvkol�y{3��,SW�(z�gC�A]4]�"�3;q�P$F4�L��[;�HU�"�~Bވ�2���ظ�l��~����Hq������x�T��ʉ�?��9��k�����L8g��B��B�����������z5�c�"5/i�iL��}��O�f3u��⵪&-o?�?4h�C�r�h��xk��\d���r'b���H�r�7�X�!�f�q��Cd<�Yޕ�Ժg���|�����hR���5�pF\ғ���͵��H9��w��@S��5.�Հ�$v!����%I����tT>^����Bwd9�i����:Σ�:�[ʮ���#��߈���1S�LMp�Ffy+�q
���* 3ċl�V�_�w�hi*�ywa�)��\���,^��fF��L�b8[~Tֳ?U?t�H:��@��[���U4���ڙ@�3HMv��k�e玝i}&.�\psf]vąwN��&��QX�B��7-Z�'y2����4J t��(��@"��.M'��Ss����_Iyv�ӥ��3̫��c(jK�+���� 7>�ɹAk߱�����'���iu���g �����x�KA���݊�C3�/|O L.�	��t}\ ��5�:��m#r"��r��,�; ��
�N2Ħ
.�]x26��?���=|�}qsK��U05q��Qhh�����n��=mw��~^,S#��+@��0���u�~g���:;EJ��h_&����e<5}z�������6����\HC#RD�e�ٓ�Tͪ�n�%/���_��aP�j���$��)���xo� �8��=���t��C$����&e������&Ϗ���a�Yr(�?���i�k�~"���_��d�0�W.���Vv��B`+DC������m%�u�*o�Mx������e�[�[�-���^��-�PX�"��w�FPP��$�z�t��J�o��)Xp����E���Hz�3N���HC>��Z?p���t.���6'��TC��e�%��ǯ��3��#X� ��BJ��P(>�Thp�,:��_S���&eI���4r���΀��	��a�,�$�4�DM<>��~tl�<e�?�9�~�c'��4��n��J����N��^TR��#(�9(_�}e��T0�Z0�<�k0N&��f7��E�P �F�(C �A��~h���E�'��'�M���6���9��?k`#wB�V����U�a���Kxԑ�+�����C� ����; ]�'�DED�O�����(�L�wP�NRi�����W|�R<�KBT�Ґ(�`��gegwyV�򠱞J�ݷ����X�.x�����{�w�W$��y�b��n��Y�j$���YVƘ#��C����E5��O�d�T��� a��^[֐�e�M=>A�$�>�~�X�(oy��7l��N�m� �^߻O�V�����C�YJ��i5Q��wی�@Hʂ3��4�V2��<b��nԭ�ұ
�n}/�HqO,7<%[�yRjEnȠ4'���X�?�3f�V,#�D�����7���8s�)M��(�_�q���Pܽ���J��%i7P�2�V�W"�>5��}����uv����p�#{�����	6n��b�"}o���{��r�`�1v@X#�	0���%T�K�����a_p������P{��|s��ΚJa���*���� �t��N��Ӷ����LAN[b�������VV������4��H��<^�Ѓ�XD�'y�=����/�H�?�g&�!T!cR��)ˁP&Sp8y���B�@T\�q�c�'�$�ɻR+r�%�k�/	K�Q���w������6yw�G�N^�z"���+]�v�oE�������UwS��D_J�*��[����=Uz��t�]���ۋͧ/��LeA�����%A��O������ǋ)�Ćإ NPfsǹ��f]ߛ�t;�6�bz?jz}In. r�
�Vw)��X���<W�l>X����wA�%���$�BC��?�j���e�����xaS<�PIx�_��8�ˀ���/����-��.}�[�������jO��֪�ѱ�qo���I��f��d;���{׵�0T��@V�!�v��Ȅ�"٦�^�� ������C��W�w�yŧE�����x�7@�����yjm����XdF�K�L�_T��Q��O��U�M=y�9��W�7����s,��������27��}����B��5����V+�`S�8��-�k�jcL�����] d��B���/%"��äȟ6O�$G���(��#K;=�q�M�xs=��w�i�mDX]l�` ��xnl�!�A�4;}&)to�5��>D
˃�hӿL�7\q3b�W9gZ�/�H�s���'}ߌI���R�d"-��=gGF����YBHBlЋ�O���9DW��ƔH�%���p��$��=W�:����V�!�n��l���$,�Z8\�ŋ�ڰ��x��^
�����)R�č��{>'k.0�LowN�i_j>���/�Λ�����t���BL��l�ɺ4;�}���1�e�7y-��u�~��W��eJRT.��PP A��5�����+&�G�{�-b�b�Y��OT��uI���y��`��m���Nu�5�t�y��le\�گpf�t�B4�g؎�Dԯb+׻��X�	6��[.خ�ah�]�[�P>��%3mP%�:��>C
pm�XM����V'��f�Y���c��Cp(��vw{��Z�ϩG����6��ky���y��ի��}6����}�O2}�3����@ѱL�� ���6�F�(J��W����K���߬�Shuh S��"�&�G�P�]t�9D<W�כ!J�wF�a����ƪ�{���)��R}��`��:�f�޴�e^t
�
3���WۭF�%}��"U!�ű2 ������,�}٧񡠏�r��F���森�������P˩�=J�B�y�M�6*�gs�f��R�
җ��"EtpRA`)et5�澠m�;h�ٚ�gl|w ��wu>��Y+�x(R��\��\4��L��L�溒#4=*2Q�αJ
j�<g�C�hhڤ�
�vc�\Ȏ��B?ux�>�uq���\���"@�e(m��ȭ��3�j\ڍ��%�(�� 1xU�Ì"`��>L��,)e�pM&:���e����7�@ޢ5���ᕦ�n�w�|�՚�zZ��H/��kF سÒ�"$��*��p_��v*��W���5�����/ɶ+�P
CT�����M�_�?��о�8T���{��PXr8ި<#��G�j��$,g�6�Q�?Sq9�N4�OD+ըX21�����}"�������b�~��|�L��%N�̔I��	'�CFx����eH-�Е��7W���,֊jՂk���;!6l�5�@,��B3���ΒRk��:	`����?�m#n5"�]���Ȟ�c6n��	P��8���tp�è��$jĮ"�$���J�J�WU��!X�t�a�E�Hp�ڰdaOR����K�?��t�U;v+�	s�[>\�&�x|�P>�Bׇ���D���[U3��u:�2��U�ӳ�Y�������h^}����35)���P1�� �ջ�BVf�}!A/NP��7�Xe�P��+���:r�����[	����{.�9�w+��v��?]�/`N+NO0���U����:�D�M�4Ԯb�ґA_����VWr��!'Sڥ �_����b�z�"A�^*�VOHz�6�ӷ R YI����6��h����uf��5{���%����D����Vǖ.7%�����n�<��	�sQ)���r��=	����+��!��e�w�z�\��]���

��ݎUL<�x����,��<?��8!
o�cRG�dIK�F���翠P�I�E�]\��6���k�O��+�.�V?�9�(�t0n�R�$�R��I���r����"�PJJ�u׉��\[��`��8�Q�7�ؒ%4J�ĹO�u�q���>�H�VxoD߂�	�ѵ��w��
�<1�i�s�u������T	�a�2�y��PX�2bN��H.X�N1t����!��NYɔ��9��4�������}�%gIi��P���i٪,�S�@x�Ş�,���F�j�J*oP�Ğis]�5a��]��%%<����6��C��T��#1k�vf�$3 {��2�m�ZH�-TCq�`?��Nj=�"G]*�# ��i�q`�߾0M�F�Z�T���e�[B*S��A<�`|�oKvo8�5阍3���!5�Y��;�5w�>ˡ��P�}|����wP��]ǗÇ!�,�}:S��m��=2��A9�i\ēw�;Ŗ7;w	ג�+�H�����&����TG�?�߄"mK�'@����4ou����~���c����MY��&s����@��W���]���Dd/7cP(F�,S
�C� R���5KR�^j��h�*$:�b�"D�'(~�,[E��QQ�T*��8����j�����W����B�#x����.�׸걉���ZE��ǆ�t)-�b]7%4��Ť4?�����rR��M'�,sW�������L �r�iۜ޴��*Y��W�Q�2��^0�GEPyV���K.�����/�F����%��-n��Y�R�ҭ���Ô"I�U�������
]�?��c�J���nf,9=�&<�%��e����HP���$��&|"�X���z�'�V�@�>�����ߦ�L!±�ԣ����S��{ z�� ��ܢS��7��}erh�k��G +bX&���Yw��f�ߺ�����k�Lj�k��������k�d��Ҭ�2���vu�٪��B��m�PJ����'�m��qYu3U	�`<����m=�y�b����ް9�!�ϵ�p��y�)/�[���Jե�E��-k�=��v'2jF�W{����a\��|��z=2ͫϳ/~�v�19~2����Î~E{�o�<�%K�Kn��a�p���bе#���_w@���l�d>����Dj�	�)��=��%�U�fŪ�3���+X�Yu8s	��K��H[o�!�ݎ�nn�H�!���S$��%��-���֒��m-d�Di��xY��ï,z�MrQ�=?���rf�&1QOɼ���rc2�EB�~�k�ˣv).|�*���2�'�2�=������e���R�ޯ�Ž�9���Q�'��u�Ҩ�$C�s��$���X�����^i��S	|�ϛϪ�n�2�A3�CJ 8	�5���O8]˪��X!��3Ѭ�S�JeCȻ}D�z[���}K�Nȟ2m��1�d�noЃ����]�'�F�Z!�ُ�W�+S�6�=�m��K�� �j��\�OA+%.�|��1�޷N�J���	X��J��|D�N���'�Ny���(w�J���1�����b��}B=C�<O��j3�n��2��瓭��!/u$E꟦�S�I�꽼�
l�r��S=�]%�כT&��^{��p��h`c�u��oa�» ;��J�WY[��rn�2�spߩ��B�Â��e:sG];�֤g^L��$Vّ~�W��m��@�XL@D��WQ;�i�G���4��}�o2�_��Ԓ�XjV�c��m����[Z�)3��W��d8���b��Bʅ� �nKxF�C^�Q�S4e��=��DA5%���3�&1G���+,�Q�AuX@��mco��?Y����Q'�x3�:�c \����Ԅ���
p)�Z�pR�Qp�e)Q"�Gk��[4��L�vrۅ��T�2 ���
���'���q��z�f^E�+��x�F+�B�ڳ�U�y��(P�}
��F���x�]�c��T��S~�=��o��۵�������^��֢Ԯ��4�s�K+N:��D���\C\:BX�Q���
�٢}���|��%b��BL�#�2cڽ�\F���)Co�{��;�ך|'��Scz�w�Y$�ġ�,�U��2�����-C�1��w�&�`P#�(�LPd� {t4��F.���w-}K�[M|*L��
���&T���4�r�K�o��`N2��T0X�b��m�^�Mz�b�t_��X_�K��nJ�3�7LK��M��An���%������W�۵{D���˺3�;H�9֐ȸ��!j^��2�qZ�)x��n�,��uvY�9"
(��E(kbH\m���Y�$"V��¼m�ZCmr�B�%� >��ƭ���aA�{���Z�b�/҂��l� ��-]��P[W�t�a_���������^��1z�3�l3����3*�GvM%�������.s>�w���nĊVi�+)����Ӊ=�$�%Q�?��̓�+�:�*PV�r[{��
En S����y0�{����󂕴��`�����*�/��D݋L�?�Ӽ�R��ioR<2���rd��r9��իs�rV�KيW�^Ⳓ��XY��|̶*��{RAq����-��v���{9�����d�PJ��Rx��,�$�u E}�OT�w�!_������L���Ӏߗ|�~��I�!-�Ӭ��`��S�vdOk��n{l�3j��z�~-+2� ��39X(F�@
j̢�S�ZapG��[�OtM����敥�Q(h�rf�kôr��]��g��*2S�(��c�A���Ȕ�5��3�o��N���rT�uœfnո�Uvί�w�*vqL"[+���Xҳo���D��6�F�Zĸ_�{D��$����]dm�6Φ{�����{-���� �kq�_�)	�gr=���M>��ȩ[$�I�������D�#.RdE�4�B��̾���[9���$�~x�d��Vډ9N��1J��?k�ߩ�p_�L�IMD�����������v��W��8�����zӸ,�}H�����n���{��(�P��rH&h�嬑_�o��WV�o���~g隑{'�霊��*�����?\^���l�����4�{(�G\����,�n�ޙwA�ͥ'G����T!-����Κ,�O�;�",m8��}X�+�H�{F����,_�t�k唌�'��0���.e���yt&�.+t~#��]&�΅m����+0��j�H������>*�!��G~%6/���g���5�l9"���CW`�ϫV@tҔ�jw%�h���{7Y{Ŷr|��BY�����k�[]�s�!~��,ܮ6!{Gy�)��+�l'��	�X�_��1���љ֠I���^X��(SN,�����]}��$��E���S��v*�M�q���g>�����LE��dwt���t�c����z�N�vw7�z9�;�?�YZ4"�0��F%���G�3�%�xS��{^�7Qpw���#!Ƅ�dra44ʁ/�y�T�:����GL1�'��|5��AH�+�*��VÙ3�YXY��]ZR8���� ���a��@�3����K�����!n/w>#�(W�I��Nc���1���a� Gp_�9�A�^�dh��?F;��j�"���	19�.'$o�{a`;$S2P�
���&�ܵ)Z��x�c+*,���������Ӻ5"��|���`K}������68�_�8��O�Y�M�R,,$���[����%���89AL�#Q⧨�Jw��M�,����*R!gl�\�������B�Rp!��!b��6�L�J��>KĶm&8�~fZ�	
�䫇j$ z��n;IQ�ʄ5.��L��Κ�v�R�u�ʇ䔟����¹���C�eq��I9ˉK��1~�?6�p|
_����/����f~s5�Q�4P��T��-P��'|SY,sI�i4A��I��i�
L�o�լ��Ը��
ѽ��&½Fm�-�� 	��	���D�3�g�{��:M�֪S��Sv��=i�(1�64�����/ �iFE�O�`{^����"��N�>-�i|�S�eT� �ޗ?�UUgp����;��q��j�.���H�i���l�ؑH�~PH����B�<��>MhN	�(�6�g�Gk 6�=?)C�a/0\�rΑ�i�VI�e��zE<�������<}��Wn�;���R]?=Q� �uݬf�����3gJ�ŕsp�Y�(3c���ɻ���y���'��|�8�ΐ��� ��{�xƒ'it�9�#Bl����v�e�q������	Yŷ/E�pN�o����w��6l!>�oB�����R��z^�_(��9L�td��&c%	���֤'����V�6D��FY��a���;�T�
�O$�JP�~о&����T,(�%��_���zՅ��)�yn�%��v�~{'�rP	�ݲ�jڃ_
��W,���8vC`>�������&.�rEU�&�U����� ��`����W�,ǡ)f��I�`��Ҟ�Ec�<n��k���}�㐠�^0�߽�c�0��O�vٻ��>�f�5�M�ǥ��м�ׁ+��6�:�R����$��ַ
�,�57蘘���ڶ��mF��/*�P�S%	?}�� {��z���=	oO����a�B�U�׉�����]��S�Pg�^�M����v��@������ꌑ�;�S\����J���A��0�Z��,���t�^����A�ZՔO��a}��Om���c��J��k7�r]q%��6��c�ھ��;�{����Z�4���^�r�XF�|ta(Ot9\��T?�;�Kؖ�B<@�%�}�'��פﳐ�L�}�4�xB��� �w0��k���̂Go|�U��桮����v�8��z�[�1[���R��o%�=����jݷM��hngf����;��]��8�~X����J݇j,�DoYb�?v�"���KE3g**g�/��jF`��Ϯ	���f�pp.�F�7hd�N��9g�/��>t�y@�k����)1�S
���B������ ��mSR1~�Q%���1C���g%�m��9�{�D��y�4�W�]J�Q��&n&�|��$�<&cSa:�w�.y7��?S��&��)��Y�ZI}ɡ.� @�B�N�?���V�g���B�FD�Y��K)Mm-ޚ� OѮ�r���1@Q�*�ז���0����-�N��?����U�5KP_��Yy)��D%8�u�P��������q���tBJ����+�?�΂fȜ��Iv��W���=�r�8;��3�3M8{� ��*����g;����P�)��b�M�8�ݍ˃Yw?q4����An�g�:���c���I�ɵ�jD}[PˇK��y��*C�ל��ZI<q�!$��l�:�[2�̔��"�{L��6���Z��n֖j�����ɂM�
�wfG�I�2B�d���n�G�Ę�Y6�v�WT�0:�ALzn�c��V
���K��$��5�5��{�a}{�P�����~�,�X��XQ'���<=|f[�4Z-���P��!P�{60��dˏ��o}�N�-/�m�,�î4h�%����T�(k��V_.n�ń7�� ��SI(,'�D�|& ��"+��)�������0���{53�ehә� �e�2��_���L��,���<���L��3]��.��^
ȣ���
��7�Z�gB�`������=��])��U�h����E�;��v�9�w>���.�i��������6:��z ���Đ+c�1�C�n�i�HP����	�AWD�{�#J�E��T�lZ�	�3���	���ğ����X�U6�~�		s"^�ԭ�3��3$s5���J�����r;�E�j���jb�_\xt���*�Z7��.⶿x7KM7Cy�3ʌ��!z�b_1>����0�k���̓�2�|�=~J�:�g~�wb��mZI��k_�)e���f��Ҵ4�"�IZa����������b�$�Ƭ�fw_���A,�	/�淩!�Yx�R��r2��كF]R����%"�>�'q�MJA�[}�����8V�C'��$�"�Q��gMw7�=�-nyp���S�D�,Ŵ6��g������m��{�i�+z�<k������9k�?�k�p:���\~߄��h{�ȽWa�A��aE��GD�7M����	%�;��q#�au��u���<BLXW�qn��&�1���)���)�X�����vYg70G����������4ٕ���\�-
��J�+H�
4d�}�1*=��-��ۥ���ih)�gD�~�I6i�hG̝K��6�(8l�$�-Ľ8B'�P ����R�xrm��Q��&�CTrd�Gc���?_��8@�pP�Th�3Ő鳀��!j?�D�+&�P�F�-ԭe������b|��3�ԉ!����ӭv=�	��X*���t���E�M�C�Y�)��Ӡ9d�g�F�F_Ӭ"���Z!�DDXڻ�isA�	�Q��[�[:"��	z��K��t���-�������}e�omY�`O�z�Ϊ���lP�햛���io��p����@8�g���ϠAV�{���.b9^���E|����Dh�3��h�!��^��v_a�X�m�]w�PU�П�8��ȭ�"zL��-����Թ�'MZ�s�j��ƿ�Ot~(P9v.B#cX��&���L��*��L�0�G���M�R��`�|�/^��k8Txa�O �%�������mxp=�*�b��;S+2����糄?�GR�,i�N���Y��nZ�����Ý��rm�֌&J/��w�'����,b��I`�Fb�����Ek\7|b��gkQ@��n��I�������B�$��f�`��W�$�DW����� ���<5GߠIv��i�}}��L�6zW�{�m(��B���P�9WԄ���$�+�B�<$*���O0�^Ӿe��̒~h��e�l�`�*���~��TR��x�E�?-��dָZ����VU����C�W��
��}﭂Ύ@�U���d�+��Pf�tm��y�.~t��T����'����?�\��Q%��F�BD�H�UU[���.A���O��!�G��S}���u���/=]hT�/!3Č·���6m�  & ��s<�#��2rh[>)Cp�
s��ktЇ��S�'r�ANB���՟s��tM�Ǻ�J��T��|2��,-�X����/���` �̏�e����r���G�r|A ����
cQ�8��C,-���'e�Ǔ3u�Р����(�#�G���_���Uf;��Cn�@V(@N#MR̡�Rk���F�|7H%��zw����?��Ҳ���-C�|��9u��eSWdR�1�5bQ��Fs���: � H��Km�Jj�E�pͷ��v�z�{ �-���3�1U�Mv9��t���3T���G1a����@�2��خ�	f	8+�A��H��JF���'��`L[s�.�����cA�cEF�/=����jfB^L��e�T�[�̰����� �hE��y[�9��y<�U�����^`�W��i�#m�J|�4��E��'zV�'�~Y6Z�y�XE��Q�ιqg�Y�	tk�����Bq�_"�Nv�Y"��/�blH��Z809�����O��5��Ptt��f��x~�1�8�̇����u�<���$3��'�����E%��ף+�MGo�m���`u�����
��1�"O�Gj�M�ORY4��C/�-_����9�d��,6<w]Чݯ�?7u�����{��{
3s.,@���|����oݗ�n�H���[�mO�-�NO������{J�-P��͊е�i1{k0xI\g�A���r*�����Ei{Zu�c/E:�0�s����� ����'bQMl�*��LH\FV�V����Yö���T��6�:�4�+�@i"�x�Qpg���V�T~�B��q��
��#�dl�u��[�XB���Xh^�� X����¹����|���H��J�ɵs	�Q��]���\��g��$L�)���O4�	�k٧mJطJR�}���O!��8��=xy��z������N���)\0�)�N��Ԕ*M��a.[�,��k�=J�������B�鿩n�4˪v���.��{�E����H�u��	�	���E�	����	�ޭ��C(��2��tv�տ�[���ɀ@�4�H�gt�j�01i�P`���9Hҟ���������'�I@��id.�_�	��$�C�n+1��Wk��	.?F���RТ0�̲%1�4霃i���RI�J��&�rZ�� �щV�e�R�U�w�N���ذH��������u����M��n��A�dV�_`����.m�c�}bP�S�����WJ�i{[�$[�q�A�g�Ϊ�~��0䃟�9�"u�}�.� ����Z�G�,ty�j�ê����]��4lE�d���	�`K��(�H��P�:��H}�5
�G���c7���;��+)]&���W$��SO�`��,��4nBj�]tZ�<�fI\�w#jJĠ�%�Z$ǻt#�+��\�=�����SU����-��~3~ 4S��F�ċ�|玬[s���k�eި,�����>O��t���]�)��m�̱�4ψ���d�n2	g���$e�ŵZ�ȩkd����m�QJE2��7�)�E�O����� ,��M8�ep ȍ�I��(�����$���aEf_٬9��&Z�{<yD1�r���!�
`��s�|#��h1�olzJ2I;#p��}�2� ��@���ֺ����G��+�?NA��)϶57�{�y7��Er�Y���iz��#�� �3��<%�C�r����X!vo�/EP6�X����R�~��u==�"�?Ȫ�c����j�wb������F/�ur��K����Mx*���s�UD�	"������Q<R�e.���-��D&ݺ��y7h�/�c�W99F܇�H���M��T���h�(�N��X�fRFV��R���Ÿ�/��Eǫ�,�v��V��yɕ�����>��L��^������H���j}�'�c�@��"�w]ƿ�f�]wƻ�� ���	o��0�,�_�#n4M�)Ja$�w�\��� ҿ4�Vom��h�w���5��M$��g����ަ-�v�hsؒ��8�}<+����HpMw��%��~���wP ��Ȯ�lݭ�[+X�	�,.���/^�+y�QF8E�z@���t��@Az��Q�A뙴�v���Ք#�p<�4lm��S]/�&�ޖa�<IN����s'_��Q��K��v�g|,Jx���*�7$v,޴s�����ew�Ҹ�5��Z'ٞ,B��\�Р.��i�2e})�1E*Sx_��Wp}��"����?�;Wy�������~�^-$:�y������L�k�E�S�L�'R����B����"��6��Nx��#�e�8����������Lh��O���<���	{D�&�j 
�#S0�bS�����=4�6M�?k��w����VȤ/�zrV;����AX{d\ \���|�޴i-����
~��A�M�B#�FՖ���|4Xy�4{�ԕwj�d�'L���a�
��N�(@*���7�+� ���w]5�O��ˌ�@�� pd�����O������O��~r`,���}��:2�����ʉ�,��5cҷ3��>pa�A��� ZaS`��C��% T�sx�b����>�4bU���(�����^������I��r�y���2��պ�8~�/��Ю��%y�Ӌ_\��p�����r��0��.k�j�ǃ��ר��)V��ʒ�]�I?�0ls�Y�а��L�*�M�x7��  �S��m�X`�m9q��~z;^b�������?��ネ��
�<\e=��3����H��M�E�qiq�/_=���t�*�j!��Ξ��:]?��^Xp�I��u'֓��|�l�2��d�SkR�8�)F�m��٠X.M��20A� �^�Fi ��u�"��_�fi韥����4V��J��Th�|�, �;
��YԀ�����sa�}�髓}8|*��e}�$W��(�b�3�#�i�ri`�H���V9B_k���Zg�vV1�=1��~������ll	��lIO�����}y��8uP��ҳ��	���	�恉KR��q�k}m�/s��(��|q\�����{�_�s�+e������eGe�B����)ֽ�=�l����������{)���1�����t���*rjL�V�Z����������e�9�?�4��s?J"qX��-��d�#<Si�^Gc�����lv���8������b��%�~�S�Pa? 7����׵o$����X)IB԰+~������,�>��QC�vy'�: �+�`'~�pxy��L\����lh~���飫� H»h��2R�xŦ�KA�i\�����U��)u�l�BA�>�h�dÌ&/�6��F|.#����J�K���r����<Яz�SQ[cR��X��Xy��ߵ0���TO�wfe��&I�'�c59�I|�d!ڜ�@A���=3r�{O(�Z1�����BS�VR��~'�e�[���Ą�<
y<���+��;��h���5�/f�1	?U���2�~����/���9K<T���Џ�c��뭭n�ח��+2��ȁLԩ@�����O�TDT�����?W�T�O�5N4~�G�D�yYĸ�ϫ-��6��k����j�S/A�����R�|��-��H�[���]�Z��*z�i�>45 E��ڬV�o�&���`��e
�1*���+!|И�	K��5�fI���i;ţ�͘\e�G�=�G\�HP4o�u��}T'N<N(�О�,����N������H���ì�P���9A�f5K�{��	:��P�Z���K���+����Y�p3B��,8<]��*|��ZR<p ��8bCј�.�1��*	MU��H�Lz���inJiGDɵ�P���L�xt٘��~G�}g^��*�����i
m/X˺Z�g]�A�D��#,9�ٚ5bl��Y����}})L���.�lf�|�RY�N�Ag����F��|C��b���W�5���ʀ���XE��o�j�@�[LC����^���2O"�����s��G�N�����H��j�����h&Z���Tz{�`W8��|Zj|�2(�� o|��(��L�����j�)��'�R�Rvd��O��'������ 2��1G��k��_d�O�{vj0�zW�A�v[i�o}�I��6�a�6��"�%�̂��\�A�@��I�.׉�p^��UmͮϞ�?���Q�^��*@�hGl�D�Xkx��F��<O_��X�nc�I7�Ս����Ȅ�k��������HW� ��$Y�:���c���z�o������GƂ�{��.�}��� ��`�����6{.������-s�]'�P5o��U^�����c�!S����է8���}�V3�����iy!�,���,�(ʘ��a:;�c�� I��+_I�8�Ɂ�;.��I�ݾ���cWh�7���LA�����.������v9�6�����2H0��ßưQK�ݰ�5M��%O�Y�Nga?���rRME��D�j6��v(^��>�H�!Ǯ켎�4V���g9��~ KQ�~�K"3�q���O)A5��~���Ǎ��>�����&7�vr���f����q������=���'"uc7G��Ye�� `1�e0=Q�l��.LED<��Vm��z��* �
�c$�	���v�zZ��J�L�/�`�}f��F�Qp��c����G4��Nvp���k��(r��[�Q�������Պ���
���*I�%�D=��]�m��y��TxR[�S2�v|ǵ�����һ�Ӏ{lN��D�o�
����R�j�`<�G	L��x�U��&��yy�x�<<-�Wmf����t)eiPp���*�D���Gy5�B��)�xF�
��.��Q�4��1g���<��W@.@���[���+�;h&�>�8辧~�Lt���N��#�:B�=�Yצ�qf�_Hz�"�P���0��9�[C�o�;j�4�5ж7:�B�?&m5��������*��h�)�\� ��w�;�I��.%m�p
�p
	t4��tt� ��T�1v��vg0̝Q����K�}7j�:��������\@˱,=����bB��t�gn� �^������6he����MQ[�����
����J��j�����RP1Ƣ�> ؾ�I�D�#;�j�����{��85f�;����=�	��R� �LѸ��?ƃ�#�O$�h�s�jG�y�]'4;�#^�b!Tc]�1�+�����82 ̊7�p]�L}U�g��4�-���\s��,��+^M	��9xM�{��y�+�,�|/�P��H��ލ��g����H���5;.���\�{�����9�D�eX���cH�3�D�A�zο?*I���H+����N}�[U�;(� ��D9�R����cñs�`Lה�9%�x�ɠ�d��]�*�h�쇆'MY���.d��ӽG��=gn�-V���Lj�kǑ)9ڊ���/���'s�'a�p�IGБt�^�������M�w�Y���<��� �����K���?Ǔ�6��_���YO�U*pA�1L>�^��x�ü˯BնN��F�x��Mn?�H����|,��נΦWR�34�\��r�cz��!��'��-��	�!:k�>y#i.j�p������Cs*�{Ao���gyn2H�_�� J��3M�1m� #Lsג�_H�\�3�\��E/�<x�e&s��;7�	�{>�~�t�Z�{�[UM��\H��9�^��8���=��$�ʆ��`Le���j�>�c��3b�phk�W��m��$Wfm�h� ����H��8Ӵi����o���OԺˠ��OA�QGQ�6:�8ܰ����4��<Al�|� �e���G��:X�nT�D���M�i���BchOK����^�8���(��wp�|يxI�D�MJ?i걯:*8�T,��2��5E��ao˂�����I]����2�/�b~�<��sv�;�+
}h�O�yK�Go �ȡO3���F�%��w� �P�T�_z������ue'�.w�N}��2HcV���֥��2��i��J����A��(-*�y;�Xwj\Sy����N�[ŌF���kh��v��Sݶ��L��ݱ�[�o������<��]�41����W �L���
��I,��M>w%�=�������BpN���ݧ�Ͷ��/ㅹ�rmTl���t�1Xu��MN8����M�Cv��1߂X^�RX�`���N4��2�x�6H���_2�d0;�?�{�d�+�ݪ��]X�)�ӗ��>�-3G��^�/��4w�����(�1�������BsP��42��P��w��Ą��@�?����,9���$F�����s���`z�k��J������t_�-{���&��V�m�:�'EI�?�C)-�hk�lK�w����<HVf-7���2�Hh�ͨ�)���t��������|�'C�N�Z��.*D���"���#M��t��E����X��%��mS��Uv��Ό"d��p�.�ԃ���l�k�v����~��"JA�dx���#8�A��w�r�Sx��9Ge�%+A�P�3�?��h���۝�)��k)*)�ӗ8�U������� �:��
��K���������G����"��\r��,K�)[^���U�<v߀���Z0e�V���Cj�>�S���d1��dg��VF���/ڰJ�֪�4�����=��MZݯ�=@�e>sIP�,������߾N�8*_��$V7Lz7���;�e�|����@p[�X4r����r���{:���%�
ϑ�VuM}��h���F�������[p�Ιڨ����#�F���2���n@?)
��=��
䃾�d��Ė?��zG�˚'��Ī��d%�C�`�u���\r|��-����|E�<ZU���Y~O�Avy���ͫӲO�`���ު5�fe�Z���F��ARF��6sS$M���ڹ�.��!�@#�� Z�&P"�\F�l����i�gA�E�� vF�A��Q�{j�X T���5�`���Vh�{��7�u������^���M'�j�*����=���
�o�,*;3��I4F�[}��T_���{p�6����B���Ld�4��R�H�`��y�h݋>���f��\Y�E;��yp'^�{�H���N{�g�ݸ!��7�������%>~¾�F����a�?�t�/(������EY��i��/'��p}0LG��g��Y���>����i����vյ��T�A�Ծ��>�� ʏ�;�6+�T>@�Z=���1���ϘMY7��o:�MT�5���F)����D�m]2��#vm�C����^XT������9��&|0^~X�����;z�@Zh�8ۣ�Tʪ�|����I4���.m�<�sV�ۂoS�/���E:e#֛���g@V��#�U������nO�5F�W��īn���O��Z�c2��n�21�]�^�����)/4|��&�̆� ?��y��̹��)����XD�� %����U�m��� �"m�P�ORm�Ͱ���ˤ��r>��k�nC|k��Q�|���4)�:R� (��:�����{�m��O�����������۔/�(���48{9�R��b�V�ztx�����Z�������:�3F���w3q�KB+�%��Q��&lDgV�zԓ�E�[����=�s�g[<��=z�x���.Ĝ=^�0`���T�Qo�S�=�"��»m����]ݬ�����j�C.t����m[k�y���~FYi�����XE��BWF�>�o;�mvgD�A��U��s15�n�о��e�~����.���̯D$}��?�`�$�@ES�QO��5d�WW��C��2��ly,��u`�||ɚ�_}0j�ޒ,���{@��8{�
��$$��'B��[Em���9׾��]!s� \�qy��;�D_bXg�E��8�Rw:�i�Yy0��+�5��<nj��ՌWP�\�F�qp
�<�O$*��7��. �QU2�]a#H�IGE	�pVl~�RsI�H�6�Q�W���Yl�p0;�@$B7νM��
��-�����J�L������8���x��O���&���Y?����bcm�B1 �F.z�H���e�W��.v�3�԰�g��^�[f�Ôcx��0�t��Tz�	F��H9q�]����*�aQ�:.�(uj"kPq���v�J)MqP�ز˚��O��,��:G�%9����O�\���iBY ��p�w;�����	�kt����X�sߤ��|�P������ῶ�Z�S�}�䍋:w�\7���M �L�7�1��Z�8�ɺɠ��,0ˢO�
����J5��5+T>0Vd��F�-:���u�#?}�>4Zf��$��O>�<��Q�[e�~k}�?���/,��~ϖ��NT�a����)�\���},��T��4��'��W񱋶�/�U]����w�T���iz�>c'���^}R��e�=|L�PV�p�z�#�s\���|�빗m�ĝv�b����e�'ͅ������@#��B�Z��CԢ1LP����B����u�VG��0^)�v,��Rr��������L������ID�?x!6�"Us�]�� �����X2������҃�ZS��� �YA+���	,s��&�sҭ=�qqH$��g\�]k&�q���
�=�0��4�S� ��Ƿ�!���V�1�j��w����֦z��}DP�|�`8j�ߒ*��a7++v��?�TѱH8�U����x�Ƹ���a���2}Z��(1AF�SV5Zҽ��B��R�q�\� &:l8\ܻs
����u�b�|���e�R��Z����z*�O�V _��k�tt��9%1����-��-o�� "�ؼ-��2M}d7HKd8��Y`}���ϑ�s�����Jfdu�* ����~˿��?����ࡁ���i����_wX����_}���g�4��R��Q�!�
����~^��9mEȮ��0�?+�D�3����1�V_��-��y0��\ԥzc����
���i����	�]�O�L��[��hXOH�)�P ��D��,t�h{����a�&�(!i鵡�$A��}��\m�f��p�9%|��G��
����e8rrF�@�R�����f�uhS�o��}����
@����3��@A�����HHw�w-U��Byݷ7�Mp��8W�z7t{��v���Kڢ�;xb��>� 쀛
;ۭsU�Ɩ��ڊ��䛲��W�2%U�5ZXG�Q� y�JFyJQ��Ԛ��I\:\��d����WZ��b�@�������s�b�����u�{���E~���s�E6=3ǭ����wQ�&�ԝ�S�QQ����`�۲�R���u����N��6��|�k hv�͗���1�4�^��)*C�hbfOQ�ɯ5�
~��+`q��Y�-�����J@�X��
�.jݬ�sP��7+�����	�����{���+w}ދ�̃b��.TC�®�8taXǏ�{�,�4����茣��Aŧ���`�b�6�+�>Mzn>uJ���������/�Ť��Ѯ�I�((�Jr̼���|�
������Y���轆 �Id��h*1������+|uE�c��P���O2�T�W��W�z��X�[�3����M$�~p����'?Y�l�� ( �3vF��k�8�*;���G(H��?Q2�(�)�	�*�:T�z��:��gy�9��y\��c9?�̷S�+��?��Ŋ�O���@����r�HC�vH*Ҡ̖�"kưw�%4��(��
wk��:tV>*�c	(�����U��RcM-񴈀'`sSW����KIH �uÞV��셄%��0���Fj>�1+$���,��F��m���l�d�n� ���v~Mi��EE�� a��@=�����'� Rf�6I#��8�s��8��+���wq'n��銯o�N2��D���J+����h�"/���&�uv�,��$6[��.��}V�ZXB�J����X���=��ߖ�L$��Z4R
q��	�*"�O����dpo&�;8��tG�^Q������ys������?�mD��[%A��!���<:v�-]�S��}���w�~Q��M�[I��?�{�	Yȅ}��P��2Ƚ�� /���f�=�|R�7~-y���'�!(�G;�p���4���,�V��漪�N��X��T��-@��C�q�*kB�����YW���0��uuY�_Tc\V�Tcx��W��R_SI��e�5.�|H*dpx?���+�։r'��<������G&��ͦ���~��(rT;�%�(4��l�ۀ�m�.V�iy*v�t�8S;�u��	��vEL��}�rSk�+���TXr�cU�T�
�it)8c\O�مD�3��P�Xz� �s>�Xa�B�+�_�e�������P�aќ�'c,BZ [�w�h2m��\D�q�q��9�}���ݩ�.�6�L��]��`���N��
�bB�*�_�~X�a�ݗ�}_חf�_��L1�C�[��sӒ����L�!5B�TΒ�g`�H�/�8�H���]�m�����Ѕ��Hz�Q=�퓋�ߘE��w���rn��Y�Vo���}�����.9A�@��kWF��� �*�9�c�@�Zؖ>.��ឞ)��͆��1���j��W���B��;��s�0�o�`�_�ga�vm{(?��(h�H{r�������oFD�*)V�M-"�F�WXw����|�]OlW���oi}{�E�9׏L����@7�9ޭ����Q�>���Y��S�j+�P$e��W6��1�6�I2�� �6�Im�Z��,����;��'�΋�9��檷����M(�4��(��Q] ��&�:��
;9�S�a7e#(�nF��nូ\�k��avB����fS�%�Z�HřTK@��#M:4�y`DX]� �>>/k{�� ��K�P���ʊ��_����W+�F���tǾ���]�6�P��˘���a��Io�f�����Tv�WH�Ê�/�4> G��k�-T7Qy��tҪ�;E�""��`
3�'�}E<��\�y�8��W����2�y�mr �����b?!�'X�n�Q��E�g%���qqZ^�¬��0����@�����SD����G���RK)��� cU����;��,om�ʮh����Î�����MJ#�����Vr��۳����F)���#��U 8q�H*��u9���Qg�P�0ٻϭ��f9n����dD�3[����������]H`��;�e/�1���L"�>d�ۿ�+�S2
�BʋzN�
y��1:�ݠ�z���M\��m�Ji1�i�_���,"̵�� ���/�W�hs�)uѷ(w�� u��)[�=�	�5����VN�E���e�R
1�i�ȃ��{8=�:ӕ����>��J'Ki���mh����0?!;1�P�{�<l������a��}�����I��ѣ�6`P�:'��L��Ǎ�S8ъ7�\W
�k|���4�xn�~����O0=&���I�ZD�T,4��P�W��rW�7�B�3^��j�^D�"(�]d"����*���)_��,�dH�0�| ��O}�e>Ս��s�;�`�./�������
�ĵ�B}�~�S�2n�Õ�����eI2Βݖ�(���s8���F}��V-���I$Y��#�(L@�:��/����`��p6,�vf��q�>^�;A�hRr�o�9�FL�P6�����+.�&g$�5u�,9���TJ�0Cm�"��(����ɵz�����Q$Y�X��AVܩX�s����e�Р��/@�c�g�)	��Ь�+���,���
Z�}�t�x�=yI11�������A0M\���5����S��������
J/��/����ֆ�x�|D�w���ey'�kG[�m���F��f�� ���t|������JrS'��� @�Q�=��N�Ո���+�3qz�)9*�v-;M�G�@��������%�ns�W|b���������k�ȸ0���2��3e��Ŗ1D����!���� ��L��U�޶ޗ���v���F�6�a^�����0&M��U e������KZ@�@5��D��?PUq7`��jD�Q�-�+�օ��D����,��,���Ƭ�Z���^;����MX�f�7[���f*�����,|Tx��h��~��i�b���^�S�ԤJP0ԏU썢���$�lҞq6���۾������$KV�$w�4Ĉ���T*��׹~u����w��V���\�Ժݸ5�A�MM���h����16s�K��pN������$U�����Ʀ�SA�|4^% t����Q���Z��2��ߨ�c�D��[ �;�\t�8�E?W��6.O���=�����M�fn!V�������X����lǅ�}L��|t�����r�]����'���X+�����!ܵ���<���@e�����-��A�@�&�:���81������%���u��/�F�t()��iD&O��oU`suD#К�/Dl�O ��5��U������N��-+��M��ӕ��β$���D���kld�e+����Mz��~F�{u��0���8��H�~gW'�xj�kE!q��K���n�ӥ���g�-ri�2#ő���,�nǋve
���̭%�jV��hOQv�`����PE�d���q-��I�\7�ȭ����Q����c�/��r��(�3�E���)�Ժݲ�
���q��n��-�\uڪ���ta����p�{�mu���o��v�N]/�Jc����7�����Z�핁����YI��}�0�`��l��É�$ >o1��D��8p"�%��6�L%�<U���34o ��醊o��u�A��TX���G#�1�M5�N��:��:�fW�� ��!�`}�!MY����4�]��[��pbte>��t�(WB��TܨXe�.�E��P��oQ��G�����jc$^E�9��H�=dF�5Ao�b���Vo�Uu`��1�l�P��9ՙX����e]��Հ�=�p�K�޺�������P
�DF�UMX�r0�>ĕLW��7�]X�y�:!w����gJ��9ۓggt�Tv0b��U�<�[4� �|�!f����,[�͎�}ia�����������Ր���:�l��AG.���t���B9+$�)B����\����ʖ4�E��1�o�:g��nr@=�����7���+{�G���N3w��������:�c���k`=�6�T�݀�6�<�ߙ�t��;��s����|�M$˹�Z�o�J��7c���X�5���-�5��J*A��"J�k˝�3�"�ƒ�/�G��t 
���Ѳt�U/�jE�}f,j�$Q�Ux�ѭAY�`\�����g�����]��u�%�~}�A����J�������ۆ��g����F}�3�	k&�ȂX\D�íZ�,�'��;��9�j��t*PF�p0��37!|Ъ�^nX�h	������fj����l��a1W�o2ݙD>����/���[�,��VǓY%ʚ1����J��ו{.VLwq�����G
����&oTڢwg�I���"��H�#Z̶�����?F%��c���n@V߈d�fL	�4��N�$�]hA��4�#29���6iG*0�t=��2{�\���\��|��}�|c �[����"��7�L�t��;I��[>�',�b�kw�t�r�B�=�c��Y��D���K7{�_�ޏtڻJPE�'3�	C��T�0��1],4�8��U�)�M9+0�9w�� �B���A�Ǟ>�=�B�JeQ��'!�O�#����M�*��2E�6,a�[qwJ1T� c�pS�>�����KY����>�~b��ܟ�f��Q89�W�5e�-`58��IBH���y����
w���{�����$���X�|\�/��=���ȱ2i���\�E{�2a�A� �Uf���s2��-��
2�O \*���_` �v���I���O�3�����2����PL������ep�ԴΦ	��(����iR��+0��.oYVD
��9CP��3�X��1q���������NÉ��G��ɏ��M\Dۙ?�"G�$�G�Z����?,��Jd�Oj<58sC�oq�RrWy�=-��ǍRԵtP��~�?O�
7E����8��6R>5T5�ݢ�����g���_kG�_�ڠԮrK�L�-��]V�oW����f�k,��*:Y{3�,#PT s%P�g
]�i��h�?d"]����9֐ù��	o{.J*��R�a1|����C��q4c�w�K���������B/"5�K��oEV�0���N%3Y�Ե�>�r"w��޴U����md
l9���"���@hv/ ��X�E=�<Ƙ���1�.��Pv�#�="A�CwS����fyqg_�A��� @��yXz)V��	,��0+x�,9�دG~�k	�d�1ኒ��g�����J�&l.��J�N���ɰ�=��#�n2aU��É*�& Ǌ�#(Wx^I�*���Ο�~U��������0j���ɉ����[jJ��{����d�̀��R�f�����F��䞨�� 3Gu
��;�:�P�	?�-�}��`�$#�A	kC�!�O�@:4��ݙT���eC����^z�Ϛ����OY*�B��˯�پ����;������)xJ֙(߅���*ZG�F�/w�4�r��J�~����Us�i8|�T�ޓ�h�$��}ʲo1�v�0�4��eH�Χ�f�L==������WI�y�T�xAn�`77$���=#ۑ3j9�Yrf���x@H��C�*x��sf+�a$��f�OF���]�7�����[�;���Q�P)��qj��@�
n�ϳ�]a�&o�1m0KD���������kƂL�X���IW�|#O`��Z�@��.�^k�(y~�-ݾ�k��n��$Be�ˀ#��gb�uL��`���Ĩ~�#*�����L�Y��&�������'���M3'�za�>j2����T'�N$�GK%��� ���R��h#yb|}�S�E��Y�%T|���"Pr^8��-3}	AX	 �o7��#�.n����N������/�J�������hʗ;!i,������0���v��� ڢ����!�'���:���>���РF�*���]�Pǌp2����I
�4q\��;�{C�����D�W�Z;���G��7���7�� r[V[M:��m �����:T5Y<�ݕ���$.��pL<>�G�DY�@��OyiGr������T���o�R�f@�x�X�Z!����*?�夑�bd�|��Ua	1:z�3P�� �ORE ��*�j^P��_�X�/d�&	ɸ�(~g�/���/=�5��v��u��%��1ca���:��ݚx=5��	��=�TI�TDƙ�L塦�1a	��it�dd� �Uw�tgI�o��0�S"�#;�ŝ�%(�T�Ai�ɥ���=/�0[��ۮ����ڞ�!�4���xHrZA\q��me�� �˦Xk�zUy�?�^�m��?��N*4r��[0� �a�s��(�h�7x0
� ��NG׍	r]�Ȩ->��Q��Q[=>Hjd<�����=�t(Fm$��jq�R��)/�C���H;Ӣ�-��L #%x��!Ы:�7=��L#/P��y�X��=�ޣ���J�`o������MyP��(އـ���S��Bӣ!΅ᛂ^`{���{���ՎM��I��Oo��vJ�ڋU4?R7�*{����LK��� �k[3�.�Η�['lo�B�ע�/n@��a����7���� �t���OOc�`&w1faB�>����5�|Z���5jʨ�o��&�,��0�ݝ��MAH��x�>�z5�7����T���(��T���feἜԬ�v�V�����/�t�C�,�j�b�g���ѿ�L~}��"������=�5ow�������g�8����H������%X���z/�=��l��$}3P/���[�$�!��FTh/t�I���� �Y���Q�}�� g�ˀU��.
B}��}��xyD`Oj9�c�Չ9�,bW/v�L���g��_o�Wj�w�N�p�p�3�)k֧EP5�disf��{p�I	*�?x��IqF��P�J/���z��2iY�ֱb���ϱM+�04������� ����KSm����b(�2� �"��=��'&��N�M=X�+cA��+7�~�qR������Z����2.2�6�FnK�g�=�") k0�K,�	Get��,;u��Wm6��"n��"ҙ?�F�,Y��t��4ȡ1"oI��(��7�f~�Y�u� ���$�j��ʡp�e"U���34C�|m4�&���$#��)����g��6V����'��wKꣂ亣Q���R�K4C�#�xa����HD���MZ��*(�X���[��X��^�f��~T�{.��M#��z*e*�J��8�I:2�+x����	8 �:bp#���~m�W�QB��6�O	.Infd#��e�ZW�L�����RǑ�#ୁ	���)�^��y/k��AG𴹑Z�Ftϧ�����4��MY��giS��tL�N�U�c�V�'��BQ������ֽ�S�.dS�
l����%�����(���}��*���w����/UR��z,[KV��1�?��M��}�n{�#Vw_M,nH�����6yG��Ҙ�13���!�áPʠb˟����b#�!�y�
c�_tl|�wOg�u�����V�X�+��_vo��g�5����(���U�v��࿌��������O���'fȴ�H.`�ոw�
�Wf�)gU^���bcn�;h�:<��t[�(.;���e4=US���zJ|��DL�i���㌔�Y�W5���������>���g���U��R\��{���m���˜LZ��|��5~櫩��5F��#p�z����^�	|鹆
a̒�Κb"ȑ�ǟj����#&�6n3w�0�:��]�q	W'��R�p:�ܮ��!u�ʶ�����B����f���e�< ���a�9����LޝV��s�ha!����'����˒��!��:*e����P5���-m%<\�q�A%��+�W6�����K��NׄP�p<$S7 ���<����I� �;75b��c�׾�%-���Y;�T��FkX_WA�d.�tXiZ�#�1�J${��MN�r����������D�����
�3#��'��QGx	��=X����/W��ӏ�}����FYߟ$���]F(�Q6�x�ߜlcB��#�5�!U��iJ,I+�5���<c�t��*�O@yj.E~�����0�O����j$/5Gyvrގ�OE <"7D����ci%�J�G*��:�ra�k3Znr��<<UTG��qU�y���vL>����q(�X8Y��4`g�ԖEdܲ��ˑ����j�^A�d��4�M�`5��.���B�J�!^z���sI0e �� G��p&D>8��z�� �s}_�[�{���iy�f��#�i�i�J���iv�Ǉ%.HHΑ�Q<�%��� 1��YGW_X����H��"Ƕ����&��!<��=ĳ��3�GI�$�D��O�K9�_%��LY�2�ڇ�B Ǿ��Y��Bu����T*Gl��x�QKH4Lb����B��K^q�5IG��ښ�.��v�%�E~�gq� }���S.٣��3�ZU�.���uEѻz� dG����c��{��Z�vc�u�oe�Y#��G�(��� ���D!�����\b��o�V�aT`��*||C-j��O��
��)��f�����2�F�
�/s�V.	��%�FGc�O��1�N�
��u�K�y��BG�-)V�������՗�����8�_�?T�%��.�C�?um����g�lBQ�m��m ���%lʼ�u���=�q����Ĝͦ�A��y�<��WY��M�����H�:���&/_�QPΏWD;�W�֫^-U�󡌉�*�۲]�O���~�?�2�X6����qG3�'�
ګ}��z#H�{J�L��d��`F,���ny���g������[!)*׽h]��v��S�Ug^馫�s��se�w��՜��*z _��yҴ��`/�+��mSXK�n����=��)㙝�w���F�1uE�XM�z�C�(kFS�Wƞau�A�{H��x�d����Sؔg�B��Gn���֚?i��,�L`�Q�WI��w�%�O�=�rl��%��k4�{�Eym�?M��W�����W����Y}`�Z D ���9��&,�z�ZEN�uIJ��cG���cj�j�P/���I�c�u/�Ux2�])$�<�	��HTx+�XqY!���q�K^/]��Y?mZ������U�1��]�J5�uإ��S�FL����;�<o.��IA�8;��3�q+V;`<	�@^�{*},�Wj����?��ҹHd�A���f�7?-B�>c`�@���|Hm�
C%DD��"۞A�m��U-)"k��Zj�r>���;�j�ДGLn�]��e��i�=������j5|F�b���"��{'("�	�J�#����|�>$�[&>���a��f)��qH�σ�y�>�䶀j� W�����^�A�{�Ǌ0�C9��w�g���b��F?�D6�u���p���΄�)K�wB=���m�Ee���Q��V��|fH��NU6� �B%��>V���x�&y\��+���e����^
E:\�<��$�`��j>�� 44��f�t�҈b^,Ȳ���݃��֥0�,>�q*ř0B{���_���E�{kG�\5$8œ��I�")��j�"VU\��_�ZKRWv��G%�Պ4'�o_
�����nƹ`A�|�)Ɩ��5C/"�*m��H|���݋�]
�I�0q�>� ԰EP���+8$�m&b�/��T?�4��GL�m�/��M���v������.�����,i���{�yF-��c����tG�2���*D����hs�2��L�!4#6� ��?�y�,t���*���F�2�|;Gݧ���@��|�fq&�9��>Bw1	oJ}�#��sɿ<V�Z �o�)����oB��=H�Xw�%��W��.7���7�'�?fջ���=h�cj��v���e3藺�����?46��mß�b� l�������q���FgͥZ7���m�Q~���K E�lrd���{�����.����%��t�S\��tt�	�z�|�;7�g*S1cV��=�Ƴ�%�f�z����您�6I%����%X��S9Z��v���C�x�|��^�v�*~��I��kj[�K3��4̊�_u�(���OF��p�c�������S~8F� �as~S�)�T�I�_^�ցǡ׋�WOf��@{�<��x3��䶥�z�����7⣷J�)A�G��Օ`	�g�e\0��m2��?�H����ǎ4�ӊ-��jCx4õAT�E���VSj�r��\qv�K/r��u�Ep.�H�����������OL���$�Q� �1��!��*%��`��G~��j��f+e�S��->���Zg����2%?��YÅ��	Q��g��2�΅�?`4;��~��f�>AO#!!khy/L������9�I|*�o��H����ԁ�2��j	&��1߸�R����)�y&�]$�	����(��1%Nv~��L�}&Е; %9��]\�Ib��3���{�hI�CY���<-��$�3�1��o�����s�lU����i�0>	���l\}I#�(��92��'�y�zM�A�+a�.j����[dI���3��}|�e7��p��꾏 �Xz𴹊�5��h%)��FG�R���فj$��ym3�a�V�\Uݚ��E�5�7L��� ��.��b�`��@��'M\�f2I��c�'�W���(�s�&
�W�W# ϕ��^��ǐA����A+>8��[=�Hg��{�Ћ9�X�5���6Aﺈn����Ў:�$�*�E�.�9�1�!����T�v�s��]��6(��nÃ?9����8���)N_h-R�Q����TW��ZZ�t���`RNY(e�+j���_W��*��	���Co��/+ m��c�l:n��$�-[֒���?S`�n8.�٥.� |� h�v��P�ܵ��lW|e�Ho ��
D�#��M������}���?&����wN�=R<�X�"���$k�+.�pO�<z�*�F��|n��K5�db����'��	h3���t0�2Y��ú:�B�[��`�UP�^�e���?C�^�KI� o�!*���#� ��(m=CmÃ|vG�������)T�ү,�>l�?�ҠA���m��f��|v>��P����W��_NE��U(̘��L��p�:����G�>`��4�ma�w�h�={���hz�	s���k(r�5��~�E(CP=�����lf����8�W�-U����@�jiV�+�dQ�?Fӂ��+M�2siN���e�3�t]y���Ah6�g`..�9��S��53�(h(x��$/k�Q�lz���U�p�P~���]�)��6��w��S��S���D�A6\9E΢{zU�ͥ��ا��4͎��*`Q�Z_g:Z��I�WT���Y{�r奤{�8Ӂ���r��Tʻf(�5���Jnbx���"��o8R�����Ⱦ ��$Fj��|�}�J�w=`��#{�-�:�й���+ƞ�%MJ��H��Tg�-{x�*˅-�'�<��}iáf�i�.sQb�k[��*����b{�HƧ�t��"���N?�?��M| [��8fuJ�_�_�C�	�����=���LOl�WZY]�$��*�*�~�����2����26;�8��+o`�2v�-���	tu>�=���}��ɕ��FhV �1�)ٽ�	����	��[�r����)�*P���uJA�x&��"[0��v�V*ϜYe�'��7���S�;+!.��<ri�j�)��'����:������q���rޢ@�O_$6��������X�n��%9wH�LG<np�C��Y�Ĭ��ex��	�O���SXWQ���AZm�TCp.ތ�O��|����@��m�Პ��$����������^���@���YyO�v3�T��#\\>B�͒����߲�S��x:�.a�֭㸷e@��������7qO��L�@�ݬ3E|m��͛�Y����4'U+�i�B�������K�KM�Hj��H�(�.�5	f_������PX�֏����:⌕�l�gT�B?a��N��F���x�3#I�O8֧�.T;n;N�lo{��+Lk�oѬ�F�M1��C�]�\���I���}�+�3l�g�(�� �Zg�ʰb`���7������l*QU/sa��󻬃 !�$)⡖�>�if*Ӵ��\F56��m/m
��XІ�L����_��IQC��OW�D�0�E�>��������#�s�ђ-�qB!�V�4�0]�:�_�����ː@�x#�;�����������1����ɗ�-s��ǯ1�R�\����aD6��ݱ^x��βDcLt���O10ЀQ]?�۸J�A ���?���N.���j �ˆ��Sw�U3�c_9s]p���z�R!v4� 4�aD��H�og��:�NbJ�P�9t��>l{�P&�M��,� �&b�]
v� �	ۧ�4�|3|x�3�ܹB�p��oX���}�O.;�39�=��21C�pm��r榆�mڑO�5Ůa�.����d�Yo� n&�ڽ��G�+I�����Z�zgzi �;"�[���5<m#���ա�)��2;�*�)�ht��F&�>K���.�9j�Ǜ����Ib=��NF��Ŋ�spӭ�ja<U ��MS%��5k�Y��\�h3���8U]��M"���L�n^����t�-�Q��g�2��٥9p��q4�0���( �G"�mn�6�|��m���q<��b��c}z���#��5�la9&���zn��sQY�G�ۆ���1�n5Jn�5�=�1��&�y�
&u8����H*C�_����8ˉt����58����]c�!Hz�1�Oܩ�J	�~����'�����"�E�P+s��.0�vD��/��;+v���A9T����4tM*���_�R�ˀJ��@쥖�|��� 4';�j�	��\ŋN���B��BHK��o��t#��U>~�}����=��?��)���U��1�Ю�;@&*1!m�wx�6�W�2> �{�)�2X��0�-�܅�n��4��7����o�O!��W�#�{ʎ��$s��N�rJ{[��پ�f�Zvld����Z�>�T�W��:Nb���(�i���/H�Y'؀ 
i|����F9r��v�-�|�U6���TY��&�z)��i�W�9j ��wDTa��2��YB��ߑR�ii�S6�����Zߐ�.l���=BP���Px���Y�qci-���.���4?+hg/u�VOD�NM�[�a�	��Xd�5�Wlϻ����1~9�c��G4@�����GޡM��ja���X,O�YT��%����B��N)=����io��g���D�U?�y/�B��������L��2����0���W����b�6t\��6�[���̀��@�_X�
�q�zV��v��\W�o�ʀ��y��lja�W�K�&=ҁ�E�P�ѱ��-�䒂��P|O�Q�g�՚t��}�>YM��a��7K�$<`�A�/}�+;ֱ�<�ˑ�8��u��IOe��$�`:��e�N����&x�}����_B�2�+�X���csZ��%$�N3q�I 
�1�f�%��>����t����Fy(�Dh�����!I��m۔�y�IE3kP�Fd�<T��������2ZKr�໊~/�e��9����Ei�|F^N������W���<�,�߮&58�Xh&K�mG�(g�t�[�[�Q���U�6S�?-T{Ӊ�	��g���	�{ro�o4��'�
7a��y#�Vp(�xK�D������5�h�9���@�#~Q��{~_t�8q�7q=��3�Y&�˲���z��������i:�|�ⲱ	��,]4��_>*z��/&yd����믹v�_L�a��7�Z!�B36_Z��/�7���nւ��yM^��6��6�8%�B&H���Ҫ8ѡJ�J Ņ�l��E�h��5��&�~2�s�9_KlF�0G!L��F�|U�ᇑ6iFrգ�xt�fbs[��6=�?ҭ�w%z����RA@�Ϡ��e��z��!��W�Zf\�a��Ч�>_q
c W�Ɯh�֣~��V�ڊ3	�l�7-��1�FU�4)�%Wn�����C��jW6~�a�F�c�P)��h�Uza�F���ZY���#�n|θ7T�8#�L= Ў�s'�;%�A��p�����n�i�RAr	��,�)��hH�$�Rs�"�~˜��6�!�b� �(��G6	���n4_O#�p�%�?��f������yQ>:��cR�FyXW<3��	�1�IX�4Q�6�	�9��c;H~���!.	j�>G�O�&p>E������n��Z�]g�m����t��}�R���NF�Ν#4�٥21@�)� n�2�&2�U�h"�t���и[�u'�UL�1�/pj�H:�	�#*6��ػ�1u�����5��d � P�v;�6���뎈��'��Rf��̰G�sמ;�=��A}EPi�0Z���/u��i�\�:�F��t䃓����~�L�(�Ky-Iڅ'a�DĂZg�A�Pv�)>Z���D�[>h�I^Hx�����4_�U��~�7*a׃��0�V����,hF,��z��Wż�ohU�Gn�!q%�gU*�*F�����#���76��$1��[0���'HȰ��3*9=[����B͆dT �\v��������W�tm�����n�D�d��ސ��,��>W{K�_��Y�W�E�!��d5*��`|v�,��Mf�u�^�r�%�������~D�����&�G;<p �A#�7�(��Y"��hk��IRK��ig���Z(.� �'�?���A��f�h�h�7w�8`+����Ǟ����y����9�^�yN���ɭǐ{����(v�8����7�P�D���i��s;aj{�X"�w��%�縱~��,��J�8�F�S��� {|h�AhLY'
���N�/{R��]+`��5�dUa!?�%.V����:�s﮵
���$�N�J����z&�������Ll}bΤ`��p�L���Ј?MV���)�;L*1&���<�Tb2����LY����-|<겒M�PQ���Mii	H0���KigK�-]���P�FN��)�cR5MɎa/]������ZL�,%�7w�f�xk.�m�n��;l1DNƏ	�)�egA��ݣHB�U�VVk���)A�Q.���RRX�vk��W�#� ��u<�jl�/��p��O���jg}e���x�LC�Ѐf1eD,,�{��s�����N�n�Z�Jal��;	NRo�þ,-�8��0��l�ZePȸ�Ó\�gM���OU�>���"*5p��A <��:�S"�ƅy"k���#e3��>Q�� �q��_��灠�$�t���V3��h�s�B�y�pB�
�ɭ_��F�������tq��-�`k5Z�J֡�A�j�c�%��ژj0�"U�\F2�k�5�H���!���m��E�C����Cg�iO�CnM�F��A앳�7���t�;������>ga���.L�N[IŒ
�\��w��#ţ��?fa���䲋�G=a$b�cK�QL0�t����a�D <�]�Z;��9��"TXy_߻Υ�6x)�~B��=�x��:[=~�s}ϛ��]�ܸ*��ns(蘽v<5����YhD�sXSA>W3�H��V�$�?ߕ��N�S	�9��'ͮ&3��B�=�4;� �"Z�P|��D����Wד�.0y��~��{�R���B6糊�4��Yj6EH�<K��)x�M����6�2� ���Q��kC�
&-s*�߫��a�˹����2��ט������"�����:B�t?�!.�BԵy�x'O�1ןtɘ9k3L���|\V@�j-���Sk�^G��=�p{�-�y@�g�
x1�������<�3�%4�`q��ԏ�IF�')�x�F�B��s�K���+�����مO诠�Zhq8���iR��q\����["c�#�ce>|�#t2�"��!2�3�P;O=L�h��?!�Q����yzM��1 w��@ܥ�Oq70���c=��p)wO�碊 ���ھ��L�%zi��q��<r��鄇�U�3su�36Y�w����c�r~hvlc�(��P�׳��X[�a���з�s� 7G�-�7w�Jy���a*���-4q}p��g�:�`T�݃�yŁ�u"��q0�Y��X��V�q������]�{5�_�A�~e52�k2u��+�rz����C�hf�1��
dy�����`'m�ў��"��w�-:�P��� �L��;�ry�����vp��a�Q��p��;c�o��%h9�p[ԻAN��ղ46��Ԥ�=�"�U���^��r8��C���q��-��w����<��}>u�(����.��]�7yt2w���B�)x�n�s+l�K�����1v��a��h{��w��Z�����k*w�i��������*T���Z��vvH@�*,`�ޝ�ZC@�hmr�Q%�P,��/[,rl������5i�d�;�E�Y
y��b��;���V
�b��ƚlA*R�]��ds�qa~��!�5��>]x�c��,A���ny���.�{��v�FMv�h�:_eG���o	]��W �
�?��r\q�8P)���ȩ��������B��A�s1�A���+�rɠ�L�҅��xն�<�,�c���@�q^�#,�Ez��iP#��ZY�֗2N�*t�2�v6�U�>��ݬ�����i��V*��c�����[��x_3�ZkՒ}��<��U��`�)��e�%���)��Z�l���F'��A���g|rGX�۱��1��a3!$���v�Cy`O���ፂ����eD[g��F�:�t@3���#�����1]oЕ|h\,Ʌ	W�$RX�d*߻SFҀ�< �X]X�i�R�鬺0О_' ��p(m�L�K|��&�a��|L7�|��o�fq�8T��qA �������G�)������>�X$�[��Z��`;a�	����
&���[%Ng)
��Ug���>>���^��޴n;�B��9TP<(��~�Q�p�t��QO��q�FĿ�4U�n���\�Sz�xP�ԊfK�Kq��Z"��H�s4Z3�B�/=��'�?l*�*,=w���%D���BQ����<�M=-)�b�:qf�J,q�#�]$�����O�w�w���)rK$ݝ���]<�o1�SO���wl(_%'�-�J�V�$�֢_�]�����̡M<�ʁ�K4�|G+�\fɤ�2���B$=�Y�=��X̛�?׏��B����|�ѥ�D�7�"
BT=6ǎ=��lH<�9ӌll�K03}
���buE�����Ug~	Y��6�'�e��)b:��*\"��G��8��
p�nY(�sdV~&x�]m	O������o�ą��Er��[S1`B����)x���;�p����6�e���ä1iHy>�W�A�ݽ6���hH�v~�h��D�MGC�;Y�+��<�cQ�%m$�B�r.
&�L�MKt2g��{ �J��8=!���u ��Q�_�t]�7 �b֋V\by!�һS����dk9�:g�?�]����k��.�I� Tcc�ћ\�.��[�a�j��AgS��g�o�s �1f�Bi*&���(š,,%'��������/7C��2�U;�*�ʙ�oɬ�������f_���)��Z�)i;��F_�b�ƈ��c�u�C���g��?(����Ϻ��ߐ�ٯ�*��b��砊c#������[Q���FC�6��Vmk��⎦�	�!U�QT���'�{����@.���2��W�1o�rp9�.�b�p�Q:���!J��4��j��/�]�ԶO���v�A������T�@��q��:g��-߉�t8#���
N�.���ɯ��Iߨ����R���&����u{�qT7�Rt)�)�RIE(�^؋���Kb� l�_�"6�m�7�#�9�l�p",1�H����o�#��)�������U�Ġ��Z�� ��� �I�dB�����3�G�,�>������#�������K�B��/�]cw�<��}A�L]��.0�ِi��VD���^�D�D�xv���k�	���Fi�����2�����]�zP�z����u I�;����?��՟�`:;z��;׹|����]�:�Z�f�HhL߭i����0<+6`�c���� ;��� �l��ܵ��0���lqp�:����X ,��E���]Xk�.�΀�?@�'O�s���
<&��˸��b9!39{�P��.;����<N�~�?5\[�2�9����|�2��6�J�Q��@۳��W��Ƕ�ެB��O��avT���扦r�~s��i|F�����&�ܸˬ e4�����I+�a	�-�0H���=���>����ۗ�f�+7*oIz�hUܨ�ѱ�C\�ё�#�1,
�l7�K �)�h`��ԏ3p�&����҂na�޶彈����Ձp/��a��	�sb[�6���C�z�R���*�=��&rd���}n|�g��*����*��w�l}�q�U�@�.|���fQ���R6���0��e��w�Mm6�9�asڨ����{/�3u��}��W�R���T��ް�&�(�ߘU�?�}�
��F�N���OfX�K�~Z��"h�����cSQ�{��1ҭ'��dRG��.KS��i �a�t���Q(&��޵(�$�G�����Q�Y:Hu�E	�b��|���?�i���7�n��DM��z��[*+U�R��p��P7ˆ�����p�-����A�Z5s�����o#"zq�� \��
�bI�On�H��<��r*��R���ͨD����p���` W�%�e1A�#�����WJ$#4Ʃ��ֶ���b�����p�pK��L��7LUPVB�"s�Lܟ�-�曹��,N
��Y���O���/�h�o>?"��,��e7��Nz	n�o���X �v�W��nj�@i���~�=V�C�l��/_h�N寍b�=�m�څ���O�"Μ����E��*Oi`����E��N�^q5H�N.�ᘐ�_���(�ȼ�.��۟l�R�"1��w��=pWN�n��Υ�Lf������}���5j��*��l��M�d܋��X�	�a�j�<E�x4]�V/�b�yH�����܈���e�s�:���>Ҏ 0�Xɤ�Pp�Џc��
h�ɱS}�J�Zmȳgl����}X:f���S����@Mx��T�l ��`�w2����Y�{�+ٵ5���2g+N��n��� 5�"���9\2C��/wX���x �k��>�M�/#r�����>���>$��s����lx�����*U�c͖X���6�U�����a@����5��
�6�'r��T��(BдTs��w3E]��R�t�ϥU:Ѝz�����h'd�s;-|�����9��vH����b�Hak�&-3�N0-[��zǭج��[�=��'�,���
7�er)��o�%�[�o�#�A�
7�x���B:t��*�]���� ����"�A��Y@Zr����?��C��Z�t
�pc������;�PY�V`����/�:ҳ[)��R���Jq����~��� �(4�:�y��p.����0�8�Q_BL�k-���)Qv�S�k��!�)�C��_�h�dx �h5m������3pIG�&�^2�4�.��XX���B�ԡ����L�{��ÕRf!R���ѧip��i�ϽP��я���t����6�;�b���m/Vk�r{V�D�E��y� �����_��z�i�9��z��\W^ ʠ�Ё^����Zq�ЈH  �x�{�ǥ�r�rr�1�UC��i@�^�i�Iȃ&�0�����j:y j��x8^�;^X�R�ץ#���bY8� /D�"�+�V�5���}��γm��
���mc?�C�Q�j*�����r�	�y>:���4��c�AЌ%�h|�oL/���Z�X��t��w����y��T��u� ��ʔ��I��M��� �/$�I���� w���GU
��a������QK�Z��o�}u�/<]��_2��� �zvc���S�����a��.�ɧ�wt�4(T��0�ߩF����q����s�?�3C!jWǦ�ɣ���4�ٽ�Y#����%����&QCa�d0K�)�3�E����Ch��=ز��D��5\��r���U?^�U�����`2��o�%"�K�c�P�	>}^x�,ya����uY��$zb �'S��9�<+��<�{	g\� �:�z�,���Ԃՙ'�{���vC��i&�B�O��ӕ�	�,�����#�r!��βX�7�B|�#��n��K�"}��"���y��%:�)���\�s�[���֩Sq�]�u!Q�DR�Ԇ��lU�Ԣ��8/W��膗ҖZ#�V�h�܎g6ȉ�xc�IM֗����Ow2��i��^�LY��z:�g2�'ngu���
���|[+�խ6g��C��� K.�q~���	��C�k3d��f�kh�WDz�8�gD:$�xK�\�B��g����c,�(B�b�R!1j�0�����J�{�bFVv�sP���=:b��L�%v$�T��%"WB��b���'���c��3���|�?q��'2{~�4Z#~D��#��?j�e�N��`W�X3���|�D����dw�uz�}�	�+	%g%u��b8�!�Ƿ1�+��c(\�6��,�J�� �b�Uőy6��L�����yd���z~�����=�2�o�
a����'�/2��iW�*�˾O��f|��E�M�E�X��5�gA�
%���Z�`@,.c��5����YN=�{wI����M��(hzu�˻�+S}al������*+��Y�3�q`K{�P�ٗI<b@��5�g����.5����z���]>����G�<�V���C��1j���خ���MYK�^���f������q��1��U*,��[@_G�V�dYT'�ý�'�4IM�	�JTF�&�A]���@r�����W�1aq�F��J�|�x��0m�)�DmmsϠE?
q.K�L$U��~<Mӵ�Ι�'b&�h@�1\ٱƏ�>}B��&�|��P����*��5��s�+�:�p����+���Mm��c�s䇐w[a�T�{�!R���<<5�Vy)�co�YJ�֟ū�ҿ�0������J��%�Ц���� ��|9��h��A1�p�x��� ��m���yNS/�b���E�G�Dx��j�YK��<3��4m8	�C���?��G�hS���������酸�1�A]��[Z�_m��b���H�Ù�ϱ�WA�p��QQ;7i���L�>P���,,���&Z���+�t��}C����V����ez�{?�������C�ϭ�H)�X}��/S�}8��SO����%���, t�]Vn�z+Z����F�KP��G���Ay����2h�f�p<9q����՚v���(Gt!��(|Dg�����2�"2�/f��s�����\�L��K~ L���?첧j�Q����s���rH���qm�>Z��X��؇�4g��k��H~܁y\�%3g�7`���Ҽz��-�cX��.���u�p���ڦ�/��Cgu^�8�l�|��/�vx���J_Ķ�W�rݹ�Mv�(T|�(&}����~���+���]�L!k��5�·s
*4�S�JpEwp�v��иpx���M0��Tk��Z����~��D�~�Q��jr�f�K���N������S֝}��Cph�k�C�1� �L�V>z�����Mp4�{�Q;AL��WRL�j�W�����څ�����]'�9�'��4���9��H({�4��L�ȳ�J����#1�,��M@�eGlB;��<���=�$�J#&Ϧ��2&�//�����f�%�����?6�����û�����Uc������Ia�f;�
����=�����Ǽ��0x��'�wt��*eI-�Vʚ�R�v�k�<��#�o<��%QH�\�dj�ʍ���n��`���f�](�R;���떖c׆yt�l���yՅ��κ�m|Z��zR�Ң�!&�:^��=�`���#yG�֛OUg����ZΕ��b�<��6sK��+��Z���[u7!Q�"��	8�Q��D��
4n�C-�w�]��H�w���QK鴀�h!3D(^�fw~uL�4�4��Y�Ԃ�Q��1��;�,tm��t�_-k���t|ɽx5սn��`7^��6��(�(R���L,yZ�i���4F�ؘy �ף��rg���7�C�@���6�%o�.;��P��t��O,��Ϻ���޾HK�UL��Ɛ� :ʡͽ�O妌ی�Xac��T�"-��#�R^>�����\���B�k~;D�z|��K�e�/���h}SOF���u�o\x?��1{a�b�`�G�)���+J�����w_�m�C�K-���}Ef��`jo˓\ �SQ�����H"IOv�|j��^uCR\�A�l�Q�����'�?���)^*$����&@���KߣϹ��oA{z�Ӱ(��[c�9%�B9��,�B2�$��O9\�6l�oҺ�2�>Ɍ�({�G�YP�S�+��U�!���������WEN�����q �=�R�l�ES7F���-��(�x�+,�t���?H.HGa��7��٩-ǎVJ��\`8�=�S��Rد>�a��BB��f�^&�(��"C���6o�+�3��u#w[�b�Ɂϙ2F�?�s%Z���"{ U[a��W�'nֽ@na��N�P_���g��QL"]���g�u�T����^$@X2ڼ�P���	�k��)� S��/B���o\Ѱ��J���������pW�Þ^�΃�w�#.�3<��]��o���9�$���]2A~B�=珽 ]��"H���8H�b{����x�:�F��ɵJ�s)߆��'g��K��0�S@.�)���CU)�YV<D~v�f���s�`�}�9'��׭o������d�~B��2�Cꬢo�v%]�؛��̥�b�K�V?վ��a�P#{�@4�!��Sf��ɴ�:�h��OiP8��E,����\r�tP5���~�b��	�۾B����V�G+�q'c�Ǒ�c��W!���y�� N�D,˸:�%���{`�%D,��:3R���d���kD�:�#�d��4�������m��#�$(F?e+?���i0�4r5S�ޯꭗ-u��4=�H�Is7q�)(�" t}PB��[��']���:k��k풼g���ّ5�b熚�5�t/U�:���{_Z��˗UxDk5jU�p�3�~�^1Nx�`�$i��c���hY�>�ն8��:��H�f�S5@Ϝ���^�W�7��<��	|�X�`ꅟ�hM��~�� ��,۵%��W����8H	H8�h�~����T?�&�Qʆ�\�U��W|��x�����Q�6��Fl��*%/_�����v`�R�l:�����n�=��R��Jm��8�3�4��*{�w��O�[~�v!�K͆6�(1�,Vb��B�å�A���|W����Hը��X���SmYI85mY�l5u�^2�x��x��d9eQ��}��7II���x�NQ6'���v��7E��O�۠�N��ֲ����:�Y�U��x��iNm�v��T\7[�d�0ߕ�3��Nډr�E���W��tTT�M��G�^x�	8�u `��d�j�%�{��5�C�.���פ�)�N']�!�ƒ��l�3��+� \�A��Y��p^#NQ:x,�51��zTɿ�t��TJ��vW_���$3~�Z6;k�ruµE��K_#����q>=��d$�`W��XW���5���,=��Q�bs��d�6�Pʋ��~�j��T��3��Z���0���yv���o�P}������uHRw�^ՠ�Yf�s>3���Yl��.�Wt
����p��ŗ�.�~�b�����A';Ԧ�;=�����B���Ɯc�<��d ^)����0s������C��O��c�_�L�o����Zx�X�Ё�$&��X��|�ɱ�4No���o��m`��0˭SFk���Nٗ����PD��Y�=�0&ZOW�� ����B�!�9<�:w���E��j'����˲�gl>���ю?��� �-&�P*���k|� �{4��N��^.�������E���(w�E�x�ZV���[�A;��geJ#��*�c���I�Ab|�(��͑���G�Ԇ�/yz�d� M��V4�HlM������*�կ�v�h1�% 2pJsЂ(��\���q�K_���
��Q�����>;�ep�L��S>��6��5��t>�����O����A��	�e @x��� S��ᦢ�C?.L
���<� K]�v	��#{�kW#���Pi��#���°p���γ�5NJ�5������x�Ǎ.�NI}�H%
,J6`�V����t(�g$��)�ݙ���<x�҆�އ_��F��D쭛�ܽ�<⇴�9��fd)]����=6�!�8H��9��rPZ��d��оٸ��/~A<A �hÚ���9F���G���x=���	�K��d?��_>�V߳n�"�~��v��ƞ{���@;���y0���,ϒ�O�j O�1�41��}�W�Yg�>Y��b�㎄\\�̝����*�)�P%x�,}9WA����Ub|��F��n��:��.�a��S��c��mdr�_2�|Ѱ�b��~R���bd���i)ȉ(��j"���0��i����$�Cj}��r�]���O��4��G^��e#	��c��(4��F{�k���W����F�.�5�4V妀���Ȗ�q�@:��zAc����޵.���U#�C��'��%���r3�'L�9�WDf �k�����=ف0��uF�Ff~g��2��G��5��<�~�����.xt5_/�r�k'���A�|է�mOkSϗ1_��1���ܘ2;/k`蓁I� �)f'�P���^��ӡ��8M��;rZ��l��&諣�ޘX�Mn�h��`W���4��g�N���{����1�6��*X�A-W̲V�\�\�^mI�Ɨ{W2:��`]��3��	��[��@��;�z�ٛ���@�̳���S]�8��L���t#(F��{����*�G�6�U�+�uTjSl���%(嶢�G��Y��#׼~��z��{�H��H���+��&�R��[LX� ��6���;Â��w)�(��F���@F�Y��v�Ǹ���y�O����B��6逛�A*8�FD�K{��h��Am6��Y�$
!�$��V\��l�8��=�O�p��\oR z&(�ð�2� �?)I�;o0%	)t!���>� �Ց01TAOn�"|+����h�z�q��4�N�pG� �K�G;O�䬁���`b�H��������=��SQy���K���Ew�P��zV��$�=����n*0~',nֵ_t]�����13u���tO\����$QΎ�c��F�Y�f�H�g��1i���Ap0@�)��StS��gmz����콍}hj�T _��&Ş4sƳ.{R�>&2�s�����g�j{T��#���mFyt���r�L��%�����H���e�y,Z:d��՜��;��H����Z�էm����-3�~_�a@���l*|"�y�z�=�����7B9_�j�{fi�,]<�-����i�+�$c����Q���2L�D=v�n%Ƴ��������ͦ`�\/]_!@1^���ZGq�yݫ���2ߍ����� �|"CnQ`q�;�;G��
;2�gqP��]��,���L]<�*�+�{l����E��K�q����F�Q@�� "��r�)wr�p�\f�}e	�6���O�Y�s���D�X�K4r�?(��_B�G��pӟ��qg:v��^�I4Ү���g��`��	SH�~��?w& ��c��#Z|w�&(���*8%���-�2��nS�v�M�V7p���|���ɾ��K��E5j�M�Qd��WP��n���''�u���f��fIr�f��h}TK0���$0��mu_����s����w�m.�aU����T�ʌ$>B*	����/\���=EJ'.xI�Th�΀�]�ן��܅�D�6GS��Q�ꍾ�۔�YR�jjfw̚��k�1Qc�G&�vll������/#�r05'�t�ͥd��/��}�S��n`*�[���b�Ք��WA�I��8�L�D �f�c����� ��W�I^�l-8�zڈ��E��T���GE��L
����˗�����Η)��g�O�v�k)M]5��i�?M˖ob�k� E]Hc/�C�J~~�3��'1V�Su+�%���ϫ����q�2���3�Hܶ�����~{������W��֐�˫`w�5�ؾa��1�}�n��%�/a݅�ɵ����	̅$�>�%	����<�CH��W��gQ٫uM�q�����L�h�֨S�e.��E������z(h�������K
�lo�Bװݔ�]�o�ȝ1��{_�0d�I�����d�xN�H@z���Zԃ��� e�H��[�����/~~Ch|�!�<��\�ӝ�Ft����w�y�f$�X�u��@\�Ӹ3�AA��M��ۆ��@v;�0ƞ*��w��w �xv	�=�@8n�3�_#�w���<���D���I'�v`A�� s�B�B��Jb�?�.��;���T�LTV���X;"�(~'[J��Pm�LI�尮�U.���?� 
�`�LK�]���g���0C�b?���m�<���R�R:|�蠛{��Ct������6U�y��O��ͫp�wO1�_�8��\��`�R�0Y�f�6�D ���7<�2���/@����@���6{E�Qbh�MR"�E��]�>5�
A�0b �!�F�3L'[��̅�Pv	'�W)ohI>^�	
�ԅ�O�mC\@�]7y[%8�Bj�w�<�~�?���'O��I����lK��3v�2�IXs�Y�*q䱉�lA�����/=�P��d�v�����M�]� �É�0���ĺw��� �>̥�b���O{��@��9��-��+�I��3g��i�u-&�0o�ݵ�g)���"~�c�y6���_ ��#�m5Tj�U��7��/�ʭ7w��qۃ���k?�{�L�z��&$a�p(g�Sl
����a�Di����[!m�9��H�LT������I����@��\���q_S�P��z#����&��9ީ�?�	�,/���,��g���GK(�����TZ�݉u�{�?v����@[vȻ�-���KY�#6cP.��ZS���ȥ�{�BFUL��Fw��:$@F���Ԝ�'yQ;bq�ǘ�`���,m+K��Fbdlk����2c��)+|���MO)��t�S�}�͛l�k���!ܼ�l|��A\yın+�3��1����x�˧7�T� WN�(��uK�P�i�c`)<2����2+ ��"v��9��8���fDx��,inb��R�N�wH�K�Yu��AE�>?)�+4��!-��&��ir5²+xr�c>Ds���ɲ��-v�ȯm,���|�N��`��[��t��ʴ�\�j9+�l�q��_R�D?%ig��+���W�mU�^t���:܂��|h�	�0�%x6U�	wFp�Ze�>m�Nx:E�|+=��qXun��ʂg|�P�S�'8�5�
x�W�Eb�1(t������W��O]}�c��aϏ�Z"�'Z��j?��.�������qk��D$�KmG"��D����-�k5*�S���G*��wqy^���l�5�U��3�Q�!��m�,^�~5��L�/���(�Z�;Vch�l'2�َ���&�f���
�9C�7zdѾ��>˳�k$���o�9 ���S�2~�=-�ӷ�����
(���<[�[
��>f%p�I�Ꚍ�H��[d4�Gt��+E�)1�
�a����3ܐ�r�a�vdYI����"B|0#�����_�4�(t�����K�u#��چ2�oZ˵���0i�M�/9$���y�����������d�$	H��±�Rn�0��$���<��1���$�$�?��2��)�/{QՇekE����c��"}o�� �e���"��M����-�떚%������[�%��6����d�+����n�Fg��!�qѮ���>�C}�OY�� �����w1\"> �犀ߟoZ��,*���E�[�AP[��o������kC%ۜ�����Nӆێ%%�,����\�zF�̂�@d��m
�L+
x<��_���l�X���d�,Y����'��r���0���~z������d/�#w�x�U����b�
�+jb�D�
��;{y�H��<�H��6O����*��O*k5�C���IV>�ФZ�Q0f5A��H������
"����7h���i_ӰQr0��p������<h�X��.����9�6�x�!���UR}D�9 �ӽe�9�
l�ب�����v��4b$A�[� ��e����\a�;K�F�DX[	�^��iЧ���S�o����޴S�~��D�0#a�*0ݦ���\��ډ�hZ���ח ��?r�����P�%|�J}�}Y�Ϣ�<Xd��8#v�꛻W��3��ŭ�q�i:��J�T�x-��Y+�G�����Mţf�����a�Зh�b�6�:�j��8���	yB7��k��"�Ρ����������D�E��֘Y8�*��0��C���BmiNh�Iu
�����M��.���&�*K���K �&��^ۣzu��gw�uC9;��
Eq����+��~s��U�[�5l'�{~��n!����pg�����}pTk1����V!�G��Cb5/������yu&�u��w6�*���oU	0�e�nT�1@�k@`3RĥNF����n�1"l(ԉ�"q�H~?�>���/��Kq��� G���@�/�-�Ջ^�&+��ݪZ� ��Mx�M�W��h������$ؙ1��'yw�A���k6CԞ�� ��a��o����.�0����R��0�->;�e�"��ŽH<�rZ�0hIX�6�2�y|���������ʓ�o�#.{�Y_BEX��_��R�(�������Ģ+�u��\�p}V�ۦl:�R��Ҟ��.����!�����9`����1RH����D��*4��D���|�#j��������=|Vp�D�%����a��<�w$����ԩ"�ꋙ���X9SX�W�: u)���w��;�6k�H~�#X��iK���U��pr.rBPw�K�[��v�Rr��Os9�b�F��*�G�\����];b��#+]� ����
�X/��l��j��N&�nx�&�C)�㹴eP(N
�L]Us��:��5�Ш=���{������z�d�U�	;Ðv+���aڵ���A�.������[�;]���;��1��:�z�p��B�U��?x��	;��,�Rؕ,j�d|
>����C�=�bb��i�d<��6	˪��A9���=P�g����|�T�ĳ�����$���֟���+o9�B�l��ҡW�YE�0�U� �X7�����v� RʥM_�Q�ìi��?���o��#}�����!h,'��:.C�l���l��r������aX'��X�5]A<co�Ĳv�ڰ,G�e��U� �d��볛��=����������G����{SĢ��t���j�W<Ԣ�\�s��}��̙���7��0�?wlk6O�V�n�>Gvϯ�D]�qZ�+֙~��j*W7ʌ���
��X��5���5�1B����p�/���^�s�[Ok���~P����Qdl\i�N�� ���C�_%�Օ=�Pp�T\����������	2I��Dݡ��J����:])���#_���F&\���D	� ��F`���U�wFzIZ�4���_��O`F��h���J�߇ԛ��K�׎��U��(=�(���U�<��@%~
�s��3�L���j&�D��D Iۉ���Vw3��3�♳�v�x��KP��]����:c	��&�>���o1�K�t�>6���u�O�0��8�n.n���=(����	ư�Ft �4RZ�8ֵf�
��<N����ū����Op���7��N��i��E=�/��I����g|�]�^�y$���d9�u��I�m3��7���^3�'�8��-k���=��l��`.�g���ݎ����)({R��\���GZ��qNS��ECb�K�e�Kes����v}le�pD#��(���|��T�����g���$�2��q���8��
��SO)�E;c��I}��7Vq��J�n}!��1�%�U�P
+�1ZO�z{>A��D�(?H��tB����}�h%
b�,��$W
 �2J@V')����0�g��Xi	C�r:��U��{�zd�C	�u%E�����:�2���!�d��b��H�,�2��?*9����/<��x�F毧�c�3������xJ�" ��rwL٭^v�=>0�?�^v;����Eb|�6�4-�����%	�����vp�/	��y<�._�(�t���R�R�w�G����ƃo�^kN(-�N�]��I^�����9t����q1v#5a���rF9�|�j4���) �H���Y�($�*�Y�'�/�t�l�������R@�`UmDv�w%�g���0�m3��i����7�|�3�Z{
���f�l��?��H(7���Q+�q��оP��6�\h�1�R��T�\B=_0޴T�*�,�L�5[����C�����g��u
2��7��]W��p������M��I\��ўn���B5����R6�����'���G^����^�c|?����X�Nm���A���l�E0}�%޷/����*��R:��L㛙B��NS�FM#�㳄_z�q��`�}��!;�ɯ��?�����&�^�8p��;z+�5�󛇍{�H�kv�x�S��ԧp� wA�J�,�?�X��+���RZJ!^gs� �
��6�ɇ�����E��u�bc��L�P|E� 1Y
򓷂_��*�>�����Np���K�v,i��p��":iI�-�Y߆��L�	'�"fh�}�SQ��~��E-���#sm�Kṁ��|��=m����Dc !̤9�ާ�7�[gCq �6�G4��	&OyZ�Bb��}�
:�]�y^�5��E��g�����5�f�:^�h��`nZ[�Xh��	�G�p���\rq�>|@741�Q@�� �i��ׇ����?��6cҋꩾbςx�����_)�>�P�ڤ	ҧ��oS��~#NA[�4߂��3��$L07��a�}��=-G�.ct.x׳�qa�d�ƬZs���1O��T?@����-̝������/di�\3�6G7J�z�UF8UԚq��k-x�ȁ���TT$�漑;�z��3��S\��mO��?)��O'Ϟ
�H��Ʉ����2�l��$v2W��=Ϫ?������\j��sJB�	O�\��ܸQ*�����+��)N���rT� 0�Ą"� 62%�(r���&D�Tm�hs��E�:V�F�BW�9.�ev�L�v)w�b���~�>�7c̚�{�>1M�����=����xqZ�e
=X�}�>~v�0J�m���u�]:욣��-�Պ|�/M���m"�ʹ#B�v�� ��.B�x�R]S	����P
%�����|�MÚ)a$�It�I�έE ]��Ejʑ76����\��j>&���<���J>;�$-�
��9�\�˝o6Hz7t�U8i�bw��!�k�ģQ�Fa �qz�D��n|��l��q|���8��0��NG?�,Pg&Z�}}���!c�_o�!��t�f�땫S.Qq2���b�:r��3�Kbd��Q!Ry�9b��2ւ��9���\�7�.pw����LeN*�a�yDӄG�P\�.�}�_xVc�'� Զ��2=���o���lu*޹`������~;��=�՝�����d�9=�|�,ŋ�õG1k�&�Ԝe�>\hydsࠐ��J٢���y9\����s�o�?�뵲NkR��K�N��˽�j ^�;"�/B{�l�C<�S�-�Oh�֐/G\n�c#�Pu�a�	��5��DhD�!6�`�:'̡^!TѓM�=�MeD��I�x�Lc1�����i��+���̙����<U0�g�-��%�S������w�*�4q`X�!�綑K��N:�N�g�= �h��]I�O��a���q�����6��^� 2
[7�r��Υ��,���ƒub���ndc��2Z�L���x��H:�_Q����@m�����.�8T�џ��f+`�4�Y���(��5*���zU㊴�%	{}3Λ~���ԭr�0w}b����ޮF�y�-\qĴQz#-���t�ҁSd����a�t�2V.O��G�t������Z����E�ux?�K9� �+�	����)�|�{���9㴷��k@3��@�"|GP)���1��&��>|�!�����Q���-��,��ya&�N����~7��@�L5��d�)���G�"�HK���V�������A�gb/�$���[��ӿbdWz�Kί�u�
b�M��%= ���B�I��-@�b����_�4r��0�Aqh����zJ�NCG�]i��<`���ٕ3{"(xD�}�� l�l=�iWVAN�:Jb���9o�~9��m��٫{�2���c ya w����l!��5[�ϚF<;Q�%@@��R�^|��t�"�]�f��n��V���h.���؝lBI��������f�j�B�x��P�yWhq��b�^�(ه�j�"���Xy� �%�f"D����O�Y��j�渺�3#E�) ���ч�Y�VE�IIf�U�^q�J�fo�pɻ�����M�鑡%�b��I����(,��t]����N������i���#���$D�P:�X�5d�}��.���{��*��L#3��7Q�\p�i�Yӧ�'Qb�R�v �P0h��3(�of6���-�Ç��m�K��K礬���Z=0xIt%']�7�~G�>�]��/yJW��e'!��`����a��X��Ѱ^AI5�FX�%�;0�T�����z���G����P��;nce�9��|�hY���zeR�}��6�U�0|��ڭ��!�3#�W<��h	�B��ڀs��I���i�w��}��Ů�9��%�ىM��#9FkR����P���\u���i�B�h#�x�'[��������o� �3G������Q!>�}�tG˕�F���c�N��?۪��p��7�>�
���e�q���2��-�?K4mn=���u�^�{�lo��]�m�P`��R�%Ubr�R�/��s�O�6'Ok@�u7Ǥ�,h�!�d����߿�S�����{Fv�F��O��I�`��=;==O��[�>'��}��Og`)��5���k�JB%���b'����'��h�F?% ��qq}��of�Y\:_S�9H����C��p ) �QY��*g�r�"���?����:qY�N܌�=M�H+<��W��]�g���<t1^��v<O7�@/��>�c Ƀ��81iT/�9\��Hb��+<H���xT�s[ܯ1Td/��@�)���i>�3M�5݁*�|[��
�Ζ��^���O��m��;�T��#	�x���f+[
Y���&�ݽa�糭ڭ�&?�}Dܯ3��a�@@b��"�%g���,��	o�:�p��� �t�wky��D�f�l��m�᯾��`vt��j�Cz�q3�0�T�܃���K��ֲP��u�Ö3�І�Gjܰ��o(F�����w뿛ٶ���oT0{W9f8��
ϥ4�_�6p'��f��y#�-��}7F�x ����j`R���x������]�7-#NCD$� �m��/������~ic���|�8�|3���N�jUĉ��m~���p�1�fu�g�u7�8BE~�!\�荬=Y�}�f��P)�Nqo�RV��p���ʏ�k%� ��dF�M��T��ɔ��;6���>�
�;�:��dO���5J�0�ഷiБa��(�X0������]���3����@������"��G3�����C$LO��D�%K�����V�H�ﵪ?��~'���Z���P����r��툀�	�(DZ�r�5?�g��{�(Ɛ�A���^�^��eCq�Qp�]��&�����	X�߯:�v�RV%j��5�>�Š�,
��'{�����Ƈ:��Y �ٲ�L�f�(�-5�$�vR~��C��ߖ�D!ό�j�bY��>�&H�} �t�#�ړ �4���0]�EGx��ܽ?��ُ��4��[B?�W�zkq1|ಔJ������g257JOxGJյW9	&z
4粄����w��nd,v��4�9J�kS�T.� �ڰ�o$5|,c�Aϵb��ݩ]xr��ۆɸ�nL���U��-�G2��d��X��.}Z9�;lW�c�T1⻩<߫�*�!v퀰X�3�	�Z��ؒ���%g�%B�N�G�h#���&7j��@Dl_�鍯\��G���<ׁ�Fj_�����v�o퀘{Z��60��b����)l|	^�nl�~&\���:_��:�������~���~?k�����~����y �ej��vb�D�ƴu����G�qUp������&�5D?O!d�8)�)K�]�SC� Ҧ��_n��_��zn�@�A��t�7��_�j�ڸ'��hgr�b(y?6���f5pd�{<����-UW\��^B��s�j��Ĺ4f�Ep�>3��m�y�FR)�v��,�
o�����4!��Rۗ\��������"0+*=��Ǆ��ƌ�G���o�r2�}�R/�p62cW�%c�֗	�/*h<k�F�P<h��~�B1E1�6FL�6�l��ˡY���\n�I��g$���Ha�&G��vB|c��I��W��W�����7�g��,����9d�b¼p�@/xs
��vܗ$��,�^n��vm)�c鰺"�]xq��^���(K�(�>M��:m���)���\$�}	J���k,u��9�	y
���z����E%�۝
�E��vf@�28�ݦfZX����LZ22>��j�VY͍�
�h�Pʹ�H�90}'EA#B���J����I;���_|�i�?H����'pܢ��-����4:R�Y�'Z����?�/��!ѥ�>хY��󽟤�q�𒂮��B�q/�U�9h��8 �����y�ᷡ�������m#���9���U0q7;���t�~'9��L^L���a�����Qh��<$[}�$;R������cۗ��b�%��/��1�$�؋;]�yq�_�T��<]a�QV�Ŵ�`H�m	�����c�Ŕp2p/�a~�mܵ������}	� �ֽk�zޅ6������Q�扺���ނ����U>  ��HiG�A����Aۈ����x���t�Y�h <�� <��yԩ�?����Κ�R�Ň+&��Dvb!C���62�MȺ��z����r$$�^��.�[.��D2'������<Ox�k	�����V�C���`[8O��.�<��cj|�9����'M���=k� +�R<�byEGɒ�1�4]�<:ta/(�	�Y^P�%��Y�:�Z��ZQw��E��J�Pa�lX���G����VA�����+�6�fR����B��$��'ɟ�q�&kq��>S%�(v�Y��yT�+��D-����%��<�/���q2�u�ON��LR�s Ͱ%lI3���	|��n�p��E��߸z�ZB�?Ӵ֐[�����91���3�hEVS�jy�Ev�� �C��gf`���+�B��9Q?�	�/Y���3�9@���T	Ro �V��k�a(ڝ�3��P0��l�'�y?�_�T�:���q���$5���4�S���oI�#��5Ͳ9��H�M�l���p�,�� n�P��=��kS92�o�}M�@'����4u�C��A��=��{@��u1�a=r.��S�)#�5��0��?0+��7��b����]�G1�Z�x8���Drf�
�����@��
>���S����1�j�u� !Q*Jdn�7,ƚ �_㹃���|]�c�.��Wgr����鼟���%�rQEM�e����=�����Y���ϯ�*�?a�@D��O�?p\tq^�����Δ^:�?$,.�2g�Jl��A'���҉8-��C}�R��qD��m�bR�P*G�cǑ-F���J�%�;�����5M��/�����-�������N):�rj�V�s�nH)���Q̉���T��*T�^dN���_�&7��*��wWk[q�a��V�
���{�[gs�0�5^�	#z�����}MZ)S�]�V0[~��;z�O�x����Aqo�O���x�tg�u=x��酦��.Ҫܖ���Ձ������GN�=(��$j��_��(�e�'�p��j4S��vO���+���_��~���Y!��/_`Qt�+�(�]B�N��|�������U��lC�N=)�pj�T��iZt�}�v��F��CVX��U� ��w�w؋1
�������e}_�-w2���B����]�$�y�o	���kpU"�������5�G���I�)��a	^\4��}�R5D� >E;�aM�+1�f)W�D��� V(m�R�<�U���x��S�H�F���PP	vDa��2�a��G=�ڍ�	��仡���մa�̎e!RΔy%6��u(,�@_{�V�w$Ν�3b8��%R��j�w����G>����2z�fA��s���a7��GUY�(�cH����3B���a��S�˖&��@�c�7�y9{��2�^���rS��>�+�Hyv��z����\iy�3������m�T<�#a
�(�TF�C/h�i2��PŐCnp���g�{F/8"�HT���J�QA��	�v>O�����P�)[J�v��m�?��?'zL��:SL�$���E��'��_k�=SM���NoF��kk~��礙�gjw�� F����Q��.�oN&h8z��)�l��I�+Uv�%y�2��-�7��9	�?�#o�y#����N<�y�}e�?Hd�<�l�D���p�䨚��o�b9��_�<T�-+��6�8]���Z\[��Gw6G߬1��W�!-����R��)s��J/���K��clD��v�&I������������=�铮+hPE1���J ��wkA~�r���(��є�䠈��x�ƪP��ŕ�
�!|�{�M zBt��H
r^��?'�r�eQ�xFD'cwc�pКe�ӗy �خ�N٠	g�54��ݪ����W&�\aX�+Z��b����y�U��A~�Z�����ǑF=r���n��3�7q�ЙOE�q����_w^qD��%�l�8��w��ʬ��ѧ����T���P����ѐ.�h)����9��x���]��h������^B�|�$zӇƱ j�H/��F��.�@u���ssPq�*�4A�e{��x�{5��>�H�=�L�b�=�oF%���?�x�9�J�0f�QsC�i�J���B�u6#L T�%L)n
�~7��	w:fn ��?�� ���
&��Y�zL%]�zJ6��{�G|5�m̀0�XK6�6oh��m�z$�t��������	4�q��|��/E����u@�,Ac1Ql	�6:����Վoq
s�w9'zz!U �j14^�cT!�뭘�|_�~��~-�G4�?=�%2i8���db��@�6*�O�׵�d����ZH�=��j�wy �	������5�;T=��}�Ww!;�Qa�R�_1��V��8�dʍ= Md�]ldHS�4�[�D�uj(d�'��-^nx��I��*֍?����-�����]Gp<�w��ȩ���6�������-͢���<,g)�_hW�h�e�2h��pVU�A��O��}���\3���-3�9�u��j��Mn���Ϭ�a�Q!B$F�I*K�J��/�*�ebz"$yѡ�+N�	��P�8��`j�e@V�O�!~�n�@�b�!=�:��%���^&Nؠ�:�j�l�Ǽ9VԾ_[�s*��߁�Q�N� ���"	���7h	��3�Nkw���[!�8�/�����-}BGHҮ�&6]Vɤ�i�4f��E����&�@Ե*�d�k�h��9+�®d�~����*v�.���q��&`�����_���J�ىTp�l:c�����oY���-��UXYZv,h�E��ޢAG���A=��GY���{�d�2�?�4����.C�ܝ~�\�U3����	*�+&d�FNiW� �OS��^�L�z��t�B���}��W���31��mvX� c��X�M��Y����)f�օQ{�`yf���ܭ�|'��xy�j
�HE1"ࠎ۸��յY�u1@���Z��ehp�?�+��� ��H+����vf���G��D����e���	��m+@x�bNd��ڳJ]}ΊL��%�+�x�PVA�`��1�cf�N��&��B�1nZ��������R��������v7�Z��.SeR[�(��`)k�.)��"�1+���~�����D�E��ɝ>����(�D�"{�Vk�;�B��:����j�j��gb�����t�����#��PU#���l~(ԑ$��㵦!�y����X�"�O���َu=��� L���Uqn�9.2�
��pF�J��\ir��0�a���{��W��gR�_�v~�|[~7�g�G��줟���v�?Mr��f�9L^:)@��ٓ�J����@���l%�G���yp��z^�[��"ִ�~Fr}]<Ԣ_���� �T��'4՜�b���z�	�-J��2t�|�]z�d��o�QL������~�7�dR��(�:��&4�~���bt��6S��c"裘~�̢7��s�3�HVH:9��$O-���q�G�	y�W.M�G��F���WV�Y�֕�XX &ݠڊ��:��9٭���!ۏ���N�#���^v"���IF	�C�ӯ��z����N����?zȧ;��apQm���?[U0XI�E���6a���r�͚j��mo��}q�KY���)�#�*d��_�,��� y�������;��E��T%��[}���)����x�S����,��%,	t^3H@�Co��<�'L���~�(6sF&����=R�8P;��8��-�W�?��=�Ni��~��z`߼ၾ�H�L���#dR��˺H�<:��f�t��kt�gђ�8�S��;<P�9n���PV �����3s�s���ǚ�LC(�"a�/�L��j[������g�hf$@��T�dxg�<�c�0t��b�}_� 96�_�{��� �1�auw���O4��T�o���0O��	&��)0�����O;�o�L�V�B(E����W*��%7�.�^KNX?���*^�imjF�ʆ�!�r?��f	F	xL�}k�C���ӆ�1[���E65��la+ga���>��{�q��{��l�@����W}��kJ"�\�>`�N�)O2���e�_)-$��-?2Vj8��iGc�l9�3�i@E��A%W�U{�=���-���g�y�"o �r	vL �Y��?�؄r��,�}(��D�d�6w�N�,Sp?i�}ϊ,��Й:oA�Z�&�/#�
���m�HT[��ΐK�'E��͙G�/WD�+�2�+������[�~�0�tsB軅p�?��)��-�s����z���4'��3e7r��tu��ɱ�|���S�֓�f$@ަ��~S���B��TxX������.`l)C��n�o�&A�M,z@�K��۲J̫�J�yHW
��,�ɐ���)!4(��JP������'�;�)h ��7��#5�p���h�Cr�k0I�%���q��S�R�/0V��S��b�����'�/\�$�X1�@��^M��O��urK�'�N��5ռY5,�n���W-�Uþ±(]H�'YY��'h�h�gj�����s�=�FZ��1�܊�;h6!/��|ݿK�˱?��G�ﯫ��[LG֟�2���d�9�ѭg������Qi&�F��:PdO'�;0����U�Oh�o��k9��������	Dtd����h2`ղ���)h4s`GEcc��Y�J�No��?�Al/�h���ҰsȺ/
�)e�{�H=��@1��a�L�o-���&1쐱���H!%�0Qf5��#����K�p3GɘsME�@��]2�J0�M,�"R��џ���9�œ�+�s�1�����qh��g�D��d#��@\Q�;$�5H���7RMq&�ZTH�n;��lx���3�q��i��LD���Vh��G�>��g��u	�Z8�+	�C���B|b>���8Td�(Y�N�X�B�rFC�@�6�t�ʥ�@�St���#�S
&�����a;������l�g��.T�ͧ���1n_��[�@_�Kq`�0tP:f��5�#nb	f�
,l�j*��}�A_o:`��(k�6��Yk�0����k�!y�;d���o�PdS���ġ���l~Q�O7�sF;�e���� �'��n�h3�G{�֊�sD�3�>��[�ge�0�Y��O�t}���{��Ѐ�稿�\ C��<��-���	ʦ��mW==3TɃ�8�y�"�{�#[j�E�R��>�w�v�6���Y2~>�H��ϮnB�%U�Y�d�p�RwAT�� ҝ�i�����n]0�<�p9�;A-�R����|�+\���)����d�t�k̻*�[zo�a�u;������rYm�05˵���/Qn��������V�C��oV`_�͖�6tN��"�m����ʌ��*3W6�x#��`I ڜ0�;4mP�_*@,������Qo(u+����*���M�@B3pg��K��Hӊ6�Ut]�Nn�(��l}G�F^[,� S���uyh�E�hJ��=t�����K�s�dYo�!Cb2�ܨo�G���yO�Z��?=M�3�R�W_d76>
�]��\�pq��KL�W��ɐ�m !�)���fq;�`/�v�i�E9�˟ua�|�-]W�S��p0��������&�����{e=�Z�-k�H���.s���?����'����U��&|�"�W�݀!b\�u�a����'�@�
�eC%_�0C���1C3���ɬ#�rQw�څa�Z�>�3��mn�l')����D�������=�#�ԑ�z_΁B��w��T�w%{y��,��ײ�
I�~����� ���5�|�ۏ���Hk5��bd�$�'�X~�%������ؼ�II�E�����N�<�JO~�"tg��R&���P�(oY-@��$�o��c_LB-d��4��H��T�X�?�q�?^C]��p`�"P,��#&�%M�8�ǷῂjhtE�;Sp:4��;���L*�F(�����XsJ">r7�%���94����@ ����V�ν�S�g�`�g(�%c2��k��;;bSH�eE�svA���]��ӵ���Z��|�=�۴��b����m�8�)�FA�YB��կq��9Rc�Xt"[gzS�����2d ��0I�V�D���hWԴ|�*��W2��?��<������Nw�r(n%��6�8�u~��~�m�5����It��CS��(!�֮;mi�V��ZL���"�bH�u����)�X�n߫D�&�&�m��8l9@6MZ��C*��-�Zu(S������P/��wb?���P
�ܽEhwIF���@x�/�Fr��|qg��?uI{%�qMsK���E��i��S'�O���9˴�(K5z�+��g��]ðz��Թ��I5�7_�����7��䏳T��r���Ҩܥ�����w|�C'�W*�����x�dg��9�9�R
��+x=�H���l V|w��2|M�a�ב8�#Y��֠����I���t�%�����o��>@�/�t�5p�m̈q;�7���۾�0?/�£�&Ցş����=�=�����x*�x#IdЉw�	�'7V����xY��t�f~f��>�t�o90�
'y�03Acp/��c�Z|� 6	[L[e�m)OXx&	
�52�#��N�`?�;�ěh=�m��>�X2�ҫ�3�LU�j�dɫha��j�d=�|@�MpvR#S�*D�v�E������e`_����~��^hΧ�[(�hz�m���~ L<��i�q?E�}��:4l@
6�"���o<�%�E �D����&:f��$��7�gKr���<»�Hl�K/d{���>y�'���Z&2�Rjc���`��� �h�?�z��}U�o��#V5���>Z��  Q:�U��J����j�[�I����4��5�pc��)ǘ<tY�"3z�m���˪h��8G1X�iC%����*���Xv�6��`�6p�L1i|�g�o"+(X�!ؾ	L?��0b�C]TRpn!�zK�����	�����h�êս�S�̺�F�����<y�9Z�b���m��>�n��R
�K �����>�B�H��ڢ�h�} Nm>>�Q��R�Y��}�2�'3M�.S��R���f��b��<���X0�RI�Y�Hs8R���I�Ƴ�c�e�^�.��.�.�~��� �R��3t�h�c?����v�8e��q���v<���Y�Q�
�/	/���L9�}X0�vM�J���U\���y	��o�"�g"�#`Ju#(p��K�o\X�u���3m���D��;j��Y���=�6"�ɢ�ug���n'�,�h�t�&�n�}H:�o�ڟ�!����[�o�@��c�y�B��V�J�oK9(��%a��꼫0B�6�����sl�%?�����6	��rf�V}�|�F޿�`|!n�����IS���h����"��q?[�3�Z=�����)�����L�' c��zƵ�� N3Ldk g)��sW�M��a,����잳�cI���j�`�>��~u<�6�:L�Zh�8\�w�/Fq-����b�W�ݕ�����:��E��ӌ��
�BbhO���FV�d��σ��\�J����ݕ�u��+���%�/�m�~N��[2���/�)�����4\3X�S(g�(�X�ai�5�^�|��Y��N�.�~t^F��z���ڹx�(n/�dN�Z�XI�����On��֮(�_�JlP&����&�|F�� �݅ 6y�޾����va�Z���&^��9��o�%����dm�%0K�C���d�t؛���Fg�����c�pn�u#�����B�b��I��HE\4������ȏ���U&�.����G���
��G�����bbf���8����ϰ��ǝ�o������ƈK����N��n%�h�bo��Ǹ��|�"��L$S�+��cB�&�"�I<�/�
��zeb�5�9�I����#�[e<����u�����vd�|���ߒc�J�W��� 5�Cﲋ$y�;��8�n��Č��ϗ�0P��x�����5.���Xۦ�R4{�жF ����X��~
�5�(���G�F�Cr�)�^���a4t��E��q_������+ӥ� K.�ː���E�iE�O�*"�Im0'Ҝ�z�Ep����2�Ϝ`Z�AgA[�p ��GA8-��-.�)(x�9��,o��"���|'
�1��v�����v��?��VE�Mx�d�z������L��}��!�".lp� %p�=�g��Lv3o���ϡm͹`�Dt�1	Xg�9'[7����pF��L	�ۧ*E� ���ߥl�|qӚ/:���^��q~�{��k�iS~�ٺʰ\#�'f{�H!����N���*�sp���s#h�\���8�����+1	�vC����T>L�"���,q�t|���g:�����d��kh��.����8M�q[�����q&�T���Hj�;�7��U���w��(�ޝ�4���$d)΋�O:l�_΍��<�f-�`�.��5�#NH3ҁ�.pM�3���l!���Ky޼��h��\'KL9��b��/XP��!<�%E����!�U�E`|��o�1�@��5�Sm��m���G���N�i!c�e�|[�3�ʚg�������޶���r1��燩xc���X?5�·"����g�
ޓ�����ˊ�oU��	����QB2��8��T�P���pf�����Ȳ�aZ:�c���sA��z �]^���0��\>�۴�t :�#����ն'Ѣ%������%-�D���"d-��y��srvn��8%�0��Rg�7�����m�'�B ���oT�aɂ��������Zՙ{��]>�w���A��{ZU��N�	�,�k���Ҡ�C��\�s���x1�5ё���*�|�|'��F�B[�S�i�i�Md�2ԍ?�gv+§�	��U	�r!;H�u%�L��ǀF���VfQǫ~��l��~�|E��n������'ېN��G�j+W����鲚0�_\�F��,jXN�*¢���O�쪛��ڸ�bb;șǻ��*����ھ��,9P�pk�s���m���X��#��N��(<m5
�����{J5H�V�¡f�Y�z�-3�|�tҮ˷#�k�u���l��_�mCݦn0.x�����4�[I���̃�H۩��ǡʺ<#L��p��N�b�JiW��+E��|��C�ܨȢ/+�f#bOQE`�7yP*� �L(G���G�5�<&{��l�{�: M�(�!s8�$��V={$iR-��^��jH�����3h��ư�.��{Ǆ�j��=���6�rF�CYhK��́B3�7X;m��w�Aq���_B����\�nM��ě����oG��D�;^[!����y�rG��lKc�m��`�����t�K!�	����N�/���52��p�h��	?F.Z�YJ���9"b9o;�*oh>0RQ�?�NChp���N����K.!��X+i����b��u��Q���dV�ȋa��=P'���;S��4�D>]�|�*l|P��;��qzQ b��=�["�|�`�*E�D<լ}z�^#x��/3

��P�F��`ω!�Nb���2q��}�~骗9Y�8�V�v�b�)M �J��B�>;�#V��af�떱z�`p
7h�6b�s�Z�}?u�����8��.=�\�L��� �D��Ǡ�ɨ݃P�͋�'����b=J(G ۫$k�T�R>��#腫����q�s�i-�3�,}z>���i�L�'y�{��& ��<��,|ES_UzWQso��G��zL��+�8�����R�8ٻ� ���_���fȢ��ق���n�x�	[枢\��	�D���c��N�F�%���y���:���}�b����Y�%���K���?UC�t
�@��-��n9���� ��N*��C- ��N�dF9^L��Zk8��$�+�h���I���2���Y�����4�F��7[���3��gA�'+`H[޼� ����R�:S�_6e)���;����\gX��Ii}�KU �(�����.�֦���?�­h�����YӐ���� &E��7����de�TQ����󸒫�W���  �Q�}�ކ�
D�k	lƈ��G�����8�=b��X�õj����J%�B�i��9�M���N��'{_ђï��wz�]����Qs�v_Z^z�� }�#Dٺp��'ĞƁ<2!�bI#$
�=M�fM٢K�`��US:��7P)�u����?�W�"pOZyuZ����j>v8���u ga�ݣ�D3�T⪪��k�cRM���dp}��@eBʶ
U�,d�P8߳��Y!dlz ���Q#A/�g7�Qlh�	͗;g���iC������Vb5�n�$1I&~�
Cƅ��fq␠��rS�J�C�G��h�y6�:�9W�;���,���|�������:�|6���0h���4퍑57G�*�Tl�M&������ʏ�tUz�QQ�H�
蟻�#�^N�XH�%����S^>�Xs�'R4!a �97f���ҟ�&�K
#�h�XHs��Lj����(~� �S]���c
չ������AzL�}_�d�O��3+ae>�{����ƹR�{�pP�sƏ�Qܹ��=}�X�]��@�����nT��_�}�H7_��3�H,r8�t�v.�k�vԲ�qܒ_�3Nq��əO9�@��휤��l����.����],LK��}�nZB��a�CS�GZcaz6�_oI9c4�-n���ڱ�1�B����&�R$�߬*��5aէ�� ��xu���8�^ϭ��k��贇&7�)Xnt��a	Y�Ӱ6QA�QBEoK�{��ȧa٫|�i+�c|��d:�4��� x���1�
,�V��벏F��Q$I�A�[b|����Q�#���JR���C�/އ�O�z>gK�~L���<	���׉�� #�e��;~�u�Ř�Z�UF��}p]�Z;���2�ܐS4��9�Z!t E��ۚW9&�PS*�A˙����õb�Y'���ߒ������O\.� ��7�*��j*��&p��a�4�;���yb &�����HT�J�H|��S& �kF`�s��R8�[�T:G� ��(�Y�'D�4�h���r6qF�WMB�|�{\��d����ϭ~�>��Gs1(TlQ;�͌�G�%����)ȑO��8hm���<���Y��N%8�R�m-%sK���_"�e�be0�R:���!�W� �Ue/�d>�%�P�ư�#����v��6�6��@r$;s���U��89�yA���$��M�N���w�[�kXB��X�@Y��`x|�w���8��R�s�>�}O0�'�������  b��4M.嘏������������w�O��t\}'šI��B99^���OtӜ�_Қ�?��MxÏ�ڤs�S���uM��;\���/�W)�cѬ b"��.��y_b6�|�6�J�":�A��l��,��*�+�W��z�/-�W�:�w�A��W0P"2�R3g)T�\�v1￞D�C�Q�Ί��-O��.�%�op�(��-��o_s�����ݕ38��yjZ0���L����C��q\�wz(��Wӂ���:uAe5��LMyҧ���Nh42����0~)
�Ӡ����8��8�[�<��W��п�4�lK��� �Ⱥ�f%A�^|>�@꽅�v7k��
�0�-K���0"i�f(�(#�R/ؘ�苁nM�1�` 8��AZ�y�M�2р�[�%?[�o�{��_���A��DiU ��m�_�m�Z�g�Z��Da��ʽ$�P%\�,ʙ�/kՖ(��
�����D὎:g ��*���9�<J*��� �e�M2'��h,�EY���!4"���P`7U��1�����؊���9�k��!;��I\�C8 �.;+M�������uFT��1�EA-ıfدȟ�s�(TK�P�¸��ϖ��
РZ8�����㲈Aw�캣�d�ga�3�'K	��Z�ʜn����F�V�I�������-��������5�����3/�b���.���r@��8U�e���B�D�&�M�F�h���EX��KEV'�.�a���9ԦMO}Ǒv�i�ou��fqI�b�[6�!�/Bǲ6^��@Qz����]����SA���'\e��a��@��г؁�G�N�������12a�8�<��͊8�c%�z�0�Erk'��YcaH`�mL�Ϳ2��Y�
MC혣8���棑r�Ur�M>yv�04��U�����VrK,������Xٮ�����b夆��R
F/��A�O�N��g��y�l�E�*���Vj�F�b.���5������&:�Q���Nb�bg��.�GK_����z�R2�6E�}��I�y��D�������q�p�{�v��]�,��gCe�>M� �QToĲ��G��?r�)�Kݙ[�������?_/lM,�İ�>�j�Wʖ��׭ �\ا7�%�S�g��ȟ�i�5o]���ޅ���
� l0O�ŗ��
��ve�Q�c��H-��r ?}J�&�(v{gW�@��!�������<�����~����$�ts�K�Էc�G<6�[|��&^u��%��������/ mXV,Rs��D"�r�>%��G��8K��3����Zݜ�9D0����fn)�I^�y����x*�&�2�$l�O*<Mb��Dg�e\[�)G���GC��1^s������� ��)R�����b ��� =3��a���:��ӄ{A�����_�����>�g=p%ѡr�� �K���4��� J��\{;eQ`;��>��?�Þ2�|ǃ*̆�uV���^��PaQ��t��U���>`�.gfUq�*q��;dz���9OeU_���EK�����^�X��y������S�S�t��Ҽ�SIvC4v\��"V����h����=���eࣵD���Nz�Ϫ����� �b�p��J�f$��*���N=�u�=�VH]ǡ�cI�:���}�P�O�>��%
!������$�ؒ���<݁�l�p۲����F�l�	d�Yt_` ��R�8��Ë���Z'ߑ9��q�.��4�*.Y�C��M��c���2���aM)n2�=K���+�7Ģ/s�k�X����o�Nµ�������2�)Wd2%��Cc��8<_�a�@��_���gd�i�^�Κ��;�a�y5Aѫ%�g.=,x����}&��̺����	����v��dpFv���S��H��_�.�zV�|C�MG��\��yk�##�"��57G;��t�_چ�O��'ܛ���*�w� z6Bna&�aX-�IBfNY++|��fkT�[KoS�n�>Α8\������Gk�A�/���j�g۸�:�t�yiOc|b�`2A�N��m���C�Θ���ޓ��8�_p�=7M��>;��
pG�����b���3��#phkM��/�UJ|��٨�f���HH	5�����!W�,�L\`�ڨY ���F�+8ڙ�wI��)����Tx/FĖ\���S~�섳�8(��Vu����V���-��~q�b>�8�L�Wۉ�I���.\���g
�{Z+@x+�y~:�x�߲�Q4M��h�r���<ay�vB`Y>Q�C��i�/��,�r�h�8n��tg��N`7�~�:Jw���,�{ϴ<�
�I��.�^�w�cq��G6�p	�^ӌ���f�L~�r�����nG����V���Y�Fa
���TL��i{z�>��:�	;�VXW�r86�@~��H���fප|�h�I�q��sGi�xϴ�H%��	7����s�愌l�]}��Ob��Ҹ���w��]�c���Ճ�zZPԡ������!���=,Ci�>�NO��.7����aYu`02~��֤������=��Q�)���(��*�8?���D�Љ��E�Q�k��3�t���r�s���l�ܟ��c��?v� �HQ��e؃I(cu�	�.L~+����7���Y<����i!���D�{��ɲsI����$��T�-kR6I���e�|��VW/���M[JX�3F>�-�*�Mهd��`bBe>e?��V���T3J��B��(M�⏌���OGk={��\LÆ�<�v$<�'�c J��%D��a� �j��W�;�>[��Q J��mk�.gK�zy%T�;�o�N0�	��z��4�U��(Ԅ�~����о���1`���9�z�+0�6�E����~�2(���c<��/��G�J�}+�x�)�<��.�����:	�Z�!,bz_d,�	��*�
o�+�o~A~i�Ut��x����x��'�`�qhNm@�ہZ6$xz�"#fB�\�����2����w���A+�])�eHn�o�i����sPZ:;犄�y�6I߈����+iۖ�b'Z�j����f���ks��T �+�ɫ��Mdm��>,�֞���
�*<O���)po1Fy/N�3��Wf$u��r�_��P��8C�$;�8�K���ySS+�����`1�xðY'�����oy�:����H
o��]�ʝ���N��sV�X��鈢��s�iLuXN�u[V+Q)o��A�hs�?�/W3c'�@�֠買F-�x����j�Y3�����KZ&�� �6VX]���C���ˆ�q���]�E��1��}'���&2
cb熜��B;��%d6��x��?W��4ػ!�ѣz]�1F�g�_�j;��!\W�?�|NrȚ!�*��Y�ɝP��s��s��*ݤm�/rj^JJ�4!6k CXu����Zr؋��3BP�lS�AyӟSZ���b@�?ʥPx���m��0�$�Ȱ~�j�;�i�^�҃N���{lkzk �o�
H��R�F����m׍���}���1Ѓ4E�ViwgOs$��,��H��Q�Z9������o%'��2�d��L(i�֝69 �L��)5O3�V~ذ{�Ukx��m���DA�����	����Pvv�!G+��۹Mfnϣ�v�6���Fb	��D��#���	�DF��q|�$?|M�f�C��Ʒ1���ܧ����(�n���w�Oc�w��o��ӟ�l؛P����h�0 �5�#Þ<g��1M(c� p�"^2�N)9g�RٵO@���\���+TX�&�؛Z�'�q��0� �a�^3g��"��;z���1o�b�B%��i��B.�߉����{�d��U*m1�-�C	��=I(����UD������=3�*{��J�Z%��ל��:�����X,{WK�)�T����E��nG���_��Òuxi*���u�f&!��F��x�Ū;��W�T��2׃�Y�v?w��>��W|~��/��Ƭ������E�%���
��r�Y,I��C���s��h}�`�T,h3$��XJ��r��xo�`��!D�ѳ��Wb��l�t����W�r�"Y:Kqc6e��EL�2��1-%�}�&	����K)P���qB�	�|̴�W���k��^�-�@}�9���!d�E��	 ��^��_�M��+fX����������2:2�t4����|a"=������'Gm���V��k���J����Jo]�Ն��®S�h�u��S���*�׼���4�嬁$�Ao5�=���®���=}_���ݝ�2�.V� [KG������c
�Y���p ����������n���w8��~B?!�|��#��9J�{�ې��\T��,��.���Up�)���t�x_Xs�
D��e������#�P���������+όى�^I!�G��۬��zEUXuZ���`��!)�*�������f����i��j���Äs��>���ՠ.���bA�7���AS�� �/2�y�BT��[ �&V��0MQh�xsݲ3o�l��7r�5���N�����+���#����Q,�ieg/ރ�0�3rQ�����w��&�c|�F���J�-�� ���dqY�8H��mhZ�,#����c����I��F/��9 o��ϲ#-jR=�#�-V�г���Ay�m+D���ӟ�
T��0��+�'�A���e	Ǻ|�`9�hӡ�eΏS�Ab�����b P���B|ۏ��m�ǩ�ݘ|J�qH|�Oi̵M�d�&@�JԦ	
����[m�j:KGwo�Vb"���iܙoH<P�%+|��4��2�����#Uq��q�@as_Mk���:u�P����m�r��J϶n���mg���p}���i-����yՙ<ኑ��$��zyד%O�i�;��(+6,J���E9��W��a��@Њ�6�fG<:�߂EaT��EU��.��b�k���M�VVEY��Ĕ�Ԣ3��l���wDd+�d��?��Lju��	�xCu:�Dpl�Rf_�7O0�,?B)�D !�u5�n��tG�Gs����u�,�;>�x�9V�^�_��/$�o4�@���}�x���q�v̒��A��\yLp��"W��(�_O+�
J�D2�@��5�A��ѠQ�l[��/����i3��}��S#������ǘ.I;��]�I��۷��l-�B�`�k놝
O��#���Κ%���8���p]�m� �I��T�>��ȩ�&}S�-�=:�5}s��(I)��f��� ��- Q���;h׆����~J*P��!���4��O"4�qEn�Wd��*�&�I[
&�G��5}���ɨ����Q`2���2�=��5�ީI<1���ُm(f���+�4���-N���I#1Őn٬���zo�c+�(�V�N#m�lv���!�@�Th{�1P��M"�_��	rM��/PQ	�g��(9��'�B�b���48T	��sf�F�=mfr�k hC���q������`����j��A}���:���_��i����pM��X��9%c�ݟ[�3�n�qd|)E~>�7�dK���s=��>�\W#&2��I�lVt�$��2�ؤI��5Q��`�x����L� �O���(������#��qoZ�Dz�	Fi����]ԝ�һ$Z#�Ak�����zjV9)�bC�H?w�N�<(.��#CNʶ|�۵��j��߃����/�?�,BtN&�a�.��$�vik�����4�Ҷh��_8��~�����@G�P��e����FR~�5Ca�X�������>��[�Eg�y����B\�F�P���}k3�Nm�}*}>�W��xps<�m��D��v-(K� t0�h�H@����W���Z���d�l�2���b10� �c�#ؿ�Rc7U���Y�Z���jf`�q�R�{k8x׌(hK���
�#�p�x�5_m3��,X�bF?O�� ��O�i|�+->�RO��s1��(�C�k����,�2->�]��U�Z1��w�|�St���Q�J$�%���>�U��X�(��s��. "�����S�M9�M�h�k����'p@��²i�|�-�7�H�@����ٔ�j�2�}He��ۼ�r�=�7�����}x@�Pp�����ݙ���rbˈїl��0��,�1�W/�Q��)��qA�]7��;y�./���pB��%�6d��<������-h��1\���d*�^���׳�V$<L�h�94��E^�n��a7Y����fH!Pv��/4��W��"X?��8A^�QN>��f���w2��'B�\�V��yFz�D�n}�9Z������`4��p��od�Ia�lq3�OD��Ӿ����>bY����|�1�_ʞޏ�S�*��+�2lm��IU�"Tn�,���2��D���;��0#���[%ڑ
� �� ���wi�Lڍ�
��Jz<�( m�	���
Ĥ\7�L�����}��+!�N�50�ƞۨ��h]���`��QF1�4��t���!��	�HZ�d#�w!���#���f�CxZ��6�9+VuQz���w//'1��H�A�H�=�Y$�O�� Dn	n�����߾���ol�ܫ��ڢ��H�#�+Ph0�N�dN՜��0⭛V�嗲JXHh��ڃ��?�p��k4J������>�7}��'7�����I����]����O2cܢo������`�����[[-F��r�%��S��4�4���W�wP���<�Ӣ�ʛ��4��H�6[�c��+�5�i6�64C6�J�O�h�c�QA�"�TC�{����&S��?	�)׋q�{g��a`�RE��7�	-O[��`O���9ȱk�� �����'�������^b٬�Ŀ���Yl[���֍��L��%��!�fqNRL�1��TE��K3����J�7B����z�Kɯ�^�E�[��Ё�_C>U��a቉�f],$M�Ì��I�D�g��C�z�	�`�P�]u�ұ�; _�j;� �/e���T�W�Rom�^�eK:ח�[s�|�H���e�����u�%�P�j�w�0�7��m}�v�#�d��YHT�#�K���x^��<���`���wIo�ݏ�^%�̬�LM�2�j��F�'P�RŬ�#��*���D�d,uE]� �\Bú[��{TC��L�U�S�\K�=��??���~i��Lh=l�i)q{�R%.���rO@"���w�=zG�*̓/-[�O��>8W�9/��/!�$IA�w�[C�K�@��0�f.�����|y�6觡3oY��y4u���(���]m�e�b�� ��q��B"����Z<��`!=\g�y�uK2���@��8 ASU� ��0�C}e�A�E�I���!`kX}�E�9 qF|�q�}>^K��O�K#�]�'����
O�Nz�[���[s��8Yw@Pl	�eL�G3ܷJ]!M<m�tl,=�A8�Y�ʘ:�v)^lMV;8���e�1�|KW���01��~ Z����֠���qJm�	�O�V�؆�@���}Tk�
�Kb_�#U؇���	��,/�H�1N����=_Օ;��X���Q�c�r$7��ߴ'}[0x�]��/�B�������S��I�o�Q��D����o)�k�q���a���v��?�un]��sr�d���w����>p��u����Q�m�&:���{1)�pd�ӹ�~Fȕ�)��MP�<m��bޏ?�� =ՒImmYI���L^ES��!y��A��'��w�ib�v�V_"- �D�K�/�?�y�J'�{&:���z�YU�������>�.�`�I����:/͐#͝-�_��e��L�Êح�����4�������I11�.���ܯ�U찇E,�ÐV��עU$��}�����sa-$��8���.������h�:��e�5AW�]i��@��V��O̵�^��+3�"A�:�|�<i��kIQ7�e#��p�1�4����|��Z1���p�S
KE=��q� 2�U �irW�s4�R�z�>m&�6fbG$�]��,��&<-m�Ά�0Ia�mp+���%4�uS�v�e�
ҏ	�IPN�:[�}T�����E�7����iY)B.�N)Ϗ@{��9m�j��0�=bWqm�i�y�xy�[>��֏B8(����ij$�; ֦�yiƴ�jñ�@{p0���~�%x0���Ք8+d�S �N��RP����_���=�Lj��^�i�CD�l�<}hf	S����a�u�8G����c�2]]8L RҘ��rt�+����7"�Ӹ���v�7A��*H�4Xڛ3psV %��˔�tf��"U2�ɈC�Q�~j�g �A�`����!�Z�~��YM(�(Nk�[[�nӴ��f"�����=�X��بS�������J��p��RZ@��X0��M2�n���Q]���,�L��i��.vG��e�@�[�,�W�d�3j��-�w�8������@iE>����Qp�/��f�8xI-�9�b��K����K�_ �یʹk�a��
f�'��~�zv�3��<�NG�u���4��O	��X��
�]�f�z�V�c� ���)D���djD t�6��P�U�%�;����g�c��y��3|U�Ii�k�%혬��'��xy��!j���R�����?���j�wohd�m����"�̑��V�ў���t�:-s�22��=y$[��8mf�u�΋'(�p~�_�es�U����&+c���i�3k!��VI��9"��) Ű�S@�1�>��FC���V�:I9_J~P����Sme~jրp��%xZ��������Q
��b��k�"4�:�J�s[Q#�s�2(��ګ�rg7��
�ɢ]Ud2@����i@���&�6z�r:	x��R�?�M��憠�K�
-��+|��!�f��/�n�lB26�/ ���l�� ֛�e�?�V�:�Ͳ���d)E9��ب��t§8�F�/�� ��G�N ����1�}N��+y$�1���Ƽ���vط��&�����n���ڤ|�}�󓶺��C��A��V���v׸9�nAhN��mñ�+�r�W �^���{~(�[ˆ�+�������0FN��i^�m4qA;)��6t� 5d�}��{v_�̏?Z='&53e��3ݮ�-91l]-}NHd1�+Z�=,�g#���!FĚ��/Ȧ��Ls�	�G�|*��>�8 �-�^Ǻ� l������[+������ԛx�a��4���kF�b�	�݊ٳ�z-�����9�7K�Yq2dB�iu�V&rޭ:�߀w��G�1�R d���W�b�=���o�主�6�c��A'B>Q��@�u|7�U��Pf�A�؜J��P�~</*Gh�{$�E~�l�B�������]����j8VI�G�����/��S�R�ﳡ��z�5Uy���XCm�Z9,�&2U���L���Ƃ������w���Q�Q$7p��[|Ihx�̠��:x�J�Ұ�	�����l�
�:R9j�?�ƉZ����W ��z�CZ�NzH3PZ��'T��$r�g�����bU
�eϺmݎ���{�`~)��,�lRv�:3��-�O)p�]���һ`� �W���͚C{꽬8������Zw-I�$��m_����<Z�>�6�[ц��ʜ��L�$ja��VgFXtmx�ȷ"+� ��=��>�K��j�B�gx��+o�"G#vԪ��)��N)�})��v*_��2�ҭ���T	��-�ń��
 �m{)0���]|9u��@<�o�Rh#ɾ_�����J��H	�CkȬ�)�(��-~4�y�%n?�n�R7K!ڑz7���m��5'�0�D?��Ƒ�?�AW�m�.���.��u�����V��S,=�P-C��Y�
I��mId�X�*�t�ڥ �ܰ�=Ҷ4V�w�u��'���DkPW0�->��;�K+e�sM>N����m�"c�Z$��� wtI,sI��N43�s�8��%;B���i�̡Y(4��]��9d̱!S�Y��^,�AWS:kIG�9f�"U�a�}{�(##�6{YL�X�����Myf�N�`<�&�O�!bħ�cl��Z���N�<�>�H:Ǧ��32����%����x��mCS^'�ɮ㘶2��>��E''v����Q��+����� o��{_�B�+��k{ZD�Me#�;����#t�b4�Y��Q�x�R�f�^�Ѣ��"�E{�m�&�j~�5���G��A��`�|�\A
$��� ��;�K���c�����+����Lq�Ck�.,���e��K��H���w�B����t�8�u+LGK����7�&�,*.��݁�Ȩ�'|b��=�a=Q�\)�H����ԝ�ǂ��� ��n3k 6.R�<���� �of�?�|�<	���c�N"��c6�4$/v�k�:s�A���#r��7� 3�ض��
52���q��(W�y/܏�@a-(�j�:�蔣X<-	ǳ��܄�O���s�>��;��eV&�i���C ])���g&��h��6�]bS�e�	^��T"0�ip�*y;m���@��h7�2���U�Ѯ�`��k!,[��ʕ*|PO�i�<�\D���g�m{r��av���ݰ��GcBl����k�'�ɯM@X��۰ u�N��W]�A�f��|8�&]��R���ǹ�8Sf�V��~��KO�)?���ôf ����d]�JG+�9#��4FR�����6����4��U�-�#��+�>��Ƌ��Ս)!�\"??0�9��%�+�(ڬ��V�^kvy��"#��BE6ό���� ����Y�g[F��,r��Z���: ��g=�+Nfhp؝���ϳ�Mۛ�v8�x'�57� v�/)4�M�f5�5G&�L��q�}4`��;�h��(�Sv�j6�qٙ�'�]]f:C���.�Ӟ=�ʻ�;|H�'�b�
y#K,����lT��-�G��B�{zy�"�^ƽ���4��'�o��OWO���`�iÎA-��+k6uեz��\#�qϳ2��W��䈔)z�; �i���]d�����;�;o��t͢�x��Kp�ޒv
�����W�a�r�!=6Z���!����*"!�}D6y��4v���bd�8�o��"��d��3�`/Z���A�
\?�|o���u����X�K�7��[<�=���:G쒳W�}@.u�]��_S(��У	[�a����w5��:�w��9)z����?�=�����l�f;$��;8�e#��B�4�"%
�|����"'�u�ի��.��T�������}��TZ�+`H�JM�n5\zpQF3�'`j-���(� ��&��Q��i�I��U�#�T������k陳����\!@��C6�>x�@G��^X�K�Tz9�jJ�:�}��l�*<Ι��6Uar�]��'��4����@����Є�#�gw7��j��0�]�Z���(�c:��ݨT��	ƹ���H��9�-fS,��1r��o�F2��d���Rn/�����SqK���@81T{�q9���B������fo�#�VR�����/�s���/��]�W��D�gE�~�yC8'Qy�>�n��`9�4�Ԩ��r)�gN��r��n{���}[/��3e�\�����E7���V�e�e�@����Jim�E}��6m�����:��5��7켾b��ua�7�,(��E����B�9��m٘� �>�H����gp�p
����~,�z�j����"���<*<#�f"P��YH�V��/��2��5�OXY�C�ߚ�!��V�iL)?�C~z�����+�>���-�(�u��1������<�(��Ȧo�D����Ӳ�%�n�yRC�3z�H�5f(�?)KF�?+*�J@;�LFk	�Ʈ$r�_��y`���`�+��!#g�L2����Y��;�
Ʌ�÷�
r�R��'�mB���.��`R�H�eu+km0�Ɛ8�W�k@H�x�x�k�w�.��C�KG��퉏��{�3#-��!�|tÈ`��6���"i3o���@kˬ�hy�7��	��\�qb"��rL�;�D b?�	��W~�/ �X���ڋ� �R��'��ƭ0���ڗn�F�
*H@���ĲM/u�\T%��\d�^�aB����T��Q���
.v:�-�&��,�����*��ϤV�7^O,��,�SJo���F�^�wϐH$���cK'75񝾡b$f��9v��[&%�*.F��B�H�fnb�Ǐ?��6x�Wȹ3���~������ѽ����?Pz����|����U5M)h��Q�wJ�����9�,�ZԛW��S����:"�W��?[��?O�����zS0�H-'�!�B)ηx؍� �S�أx�6��xy�~��	�!�������	yxt�*{��湭<�V·a���6�����?� X'��k���=
�XXf{��~G��i{�t|<W����,�;��ܐl@~HT������څ�(�^ϕ�(�JTӷ�p��������E�ze��cS�?�7_�u[�ˊ,�˰� �i�mF�Z��N���Y��tՠ�O4�]a�M9���R
��ʉ�K�f�n��<�:�n� ��Jf
?_�,c�	�r�G�v8ńz�%���p�O�ٚ'TW]�b={'��,���J��Le�<њ��;�hp�M���]2�!.[��)���h������AΰM9��]��A�����Ȑ)�6*B���}��ڋN��=��o�K���8M��.�F�Ӷ��G���Rvk���i��f%h����sE�!P���(A�MdôZ*�r	"s}ǖ�T��d���Ij鄛L5���\�Fwvn��c>V�ݔT[�ȡ��=�m�=��f5ƥ�L�J4x�5CSϑ�S~UJ`i����n`���
�	�?;T�"o�O�ҏ��EP�׼.p�=�&_�ܹ�����-g�G�e�J�
�^U�"Ԋ:l1k�>bSǧ�9o�~�e��;�����{��bnpQP�u9Y� ��TI��$1]+���9&␒��z�aՋkU����ד�*��<�a�G�Ǌ�]�]�y��-qƃ砐X
<Cnm�2Dd�m�G=n%�zP}�I}F PkB����sI��}�����b�N�k�����)gp�L���u|1��������r(�"_J�h����(��ӲU��`�oOGt��TC����x�2L˝��b?����W���3Zj�jUQ�O�ZvR�f�=p�w�p�#�F�Cݣ�))�m~��V`
�H���f��Ide��ܿ]�����TP��k��M�O��9��j"yeǩ[���G��v?� ��̅>���鳇;���
��a����C"5(a��oN{֬���[r;���ծXz4бZZ��?JX���I�u�J�������!���@�(U+�O~7��(!K:�#Uh#x����ڪ=����6������[��4bA�ர��v��7��p��jZ��%���q�m
�_�Qg��2������ꀴ����p�l�%�P3�9%̫(3�H���uaՓ�϶���Q'�������y.�(
���n�]��z9£t,	k��/�y#���Cx��j@2(h%?�u���˘��Gs�R��M[-Ԣ
��n��V��b�+�����L�\�΋�wSr ����˒����*;�.g���mA�!��+�<B��4׾o�z�.�g�V޻����Q~���l��Zp�8������
#�����$��?����S9���c2��`�K��g�|)�d"JW���; �K�piB	ǮO�|Yvp��;:�f
�b_(\��G}�����/��\�%@�U���T���V����5�݄V�t�6�'����]{���_����;���e��G���Ŏ����gPX�fh��S�4v��N�&	|U�y�0�{��oH&f��}wg�����D,�����K|3}#��Nw�y_#��2�G0��}�( �1���q�H0�GsR2m�Ft%�(�,O���6���y&���:@�Ð���f)���F'��!�����2u��	_Ж�Ir���I�u=���/�q���.�"�|'�JP�ٷ�%DV\T�TZ\�6%)�I6k��1j	��O��q_�U�hs�ŅU���+������0�#q�R���G�&5�{^���0;=B�N��f���َ|�/�!Q�
��X<��=�[��ŵg�9G�J������&Y�YS��k�03E�,��t)���W|��GAԞ�@�9���F�.(�w��P�dD�� U���!+&�D��L�\��t�Y�a6�m�5�D�fw��d��	*��l����A�OߎഀՃ����Z��a��i����NŰI՞2i���S�
q�QAe+~E)�X�-`��o�u|��M@`�@��Ӌ1��K~i��۝c�M���QݸOP���{�����ӹ{l������dS�����'�(��#ÇI�m�$��p.b�|��u.�۴9S��{�N����p�Δ(W۬�_�i�=]���`ގ6c��+Cx����1"sc�*̍�订y�d��<�Z[�֛s:�[&�~?�v�>�w��?Ei[Фor��`����i�W'�uiJ��b8�E��IM�ĵ�S�-�wvy���g����.ǉ�x��%U4E^��ʶ�MY? �����2qY�;�����?�u�~(V�A�m[i�︛���:Ty�@$ݎ�Q�.�s!LL��e��k���)��v��3!�3Ą˚�7%�8�ٓv��H�� �Q!��gڄ9��?Q~q��͝Z���NJ�U���eH�W ��M>k+�
3.".�&⺪P�8���YF��Q�X}�%oSXr�j ���D����f����j'��cjH6��@����R�Aؓ�m�����8��0���B�W��n'udr���l� �c�f�\ɽvс��:�uT�ѧ�PAj�Rڻ�1M[O��2��E;�U�4i�X�e_�3WX@�9
�.�2�в��E^k��!���J+��x�"g����7#Y�9�?�K-�WHe��f��-�m��,�R箅�i��.˙e�5\��
�:۷	?��5�.g�����m�4Vo���X.���f�chQVN��p�o���& ���${�ㄦ�UrhɽF�<�k�X����k�y��4�0�^�}x�2��"�-I��Fgo O�P0�JvC2S�b �
O4\�j��wa��.=ͻ��u�Ø��VS�.��WF�#���A�<�]f�0s�'��"�	�Xc��E�����j��c�_���7{=r���t>/F@�y+t�>�P���tU�##�T4^��:�s�cV⥿Q�Ǒ�GfľH�^��\� ax�k���0�c(�"6 �ȘW��ٔ|�v|X��6a�RVB�6ҡ��x_��W �Pŗ��Rq��~�̵���{�,M����6:���χW�&=��-�jT/��i��������o�xMmqk/��tqF��0�)��{��,5:V�x��ؿ�T�����Ў�X�G�q�#����q%�NCz(#Tz+�xAյ3>9mb�8j�F�6>�����U�N���
=1^cX�i��v�n���E2�B��j;0d�t�bڏE�`�@�I[u9Rr��7e��Ekh?o(ׁ�m
�b|�������p1��W�C�;�8���|�<�*�6d�o����>����:^���{�z�j�ϏLim+���醌�Vꝯ{/��BQr����[���.���-���kz'���҆�Tzp�iss9�Pq��^2Y�7ǎ_LS&����Fm�3���/���ؼ���t1!���C��G�Ҍ����>'�,sV]�Z�c!?^�$ ��-I^Y*�i.y'!��T�y���I��+���z�J�@��T��%o��B�/=z�S�FNY܄4���vºޅ>��dXg:q}#�1끂C_���r�R�5~=�鎠��|��v��ᨥ����o#'�'��l�~��j��@�'��&�w a@ڈ�"��D�����fߕ��w�-/b/YV=sޤxP9�Y_5RJ�";�o����N��r?ڇc�8�V'^���R�Wϓ�hZ!+S�v�%��{��Jh��\��S|�P�-�� ګoR�pF�_q���U��M���������
�/ef�[wX�� W��"�?X�4S�������^��l����a(e��F�����5�����TO�<���vQ"HmqRSU=�*�W�xq�x`�s+]��FQq����'�CV�9��WI���iǗZ����>�<��W�y8��40%�;K|�?<��wm�C�S�O��M��jM0�El��U.U|�� P̰��
���j��vt�<E!k� �2���Fհ�MI@q?�m?�H/`D�~�4_i��(�x��'��n����#(�`��r���'n��3\����X�b�G��f7E�x��� v���C�ڸޯؗüO(/�}{D�iɗ�!�eȸ�p�����U1\�� c�H�Y�C?��]U�&���!g�J���(v��qU�2��8�@�Q?��GUV j�:�j�5IǁĘs7���8Y��ֹ��.dG�eĢ�[��)�t<����<�K�to��'��qd2��ntHl�ǌ{�&�����u�S뺹�ci����d���f�^���G��g�T��,.ˊeG�\] �(u����9�4�κ�����v��N_�b3��~b�aXwk�oa?��);��V��`v�ag�� ��sR]T���m�P:Y��.�o XI1j�����K��kq0�Q�<�v_�öxa>v���T죵�'���}�?������	$���TJ����1�/?F�I	g�mN���=�.q��ֈ~��{ݠ,hs|���_Rv�耪�0��)�}��,ˉ�UF-�4��1{�Q1����`q�,���z��X�
��s�O��{	E����:>:�xˣ1JR��l��
�;n8��g���B8�s)r��$�#L��l@�ޓ�&��������8yt�a�fQ��.&1 �Z�n���c|>���;s�%�#W8�g��I�ԍc����|�[��)'��@ 9�1��d3rA�H����\�04<["U�ƒ8Қ~�$�Y�����G�gʢ	h;�[Z	QVM�qr�,�
����E�I]+*D9h@9w��_\'����Y����WV�V���^�$}Q����^���շ�>��wy��0���Y�[�����K�I��NI��\��K8u����)}i��~�L��n���N�cԆR���6��p�x��s�|�ɒמ��X�fRm�\xڝ�Xk�[��#L��5����	>{����;"C�:^�_��(���6s���؃ ߾<fi@(xa|��N-i�Hيp:,r,�)���:���Ca�m63�KLٴ�MՉq���Sx�Z�R�Nہ c-����@D�<���Ey�pL:L��Go��A-��]��Xh����2��4Z�B%�yٝǐ	���Wqz�b�A{���?�j�
j��Β H�����Wəe��O��.�ҷ���X\o>T)ܝ8x���e�P�G��0��̼;�i��.VMpЩ��r�z���E�z�d��I&�J�`
+�@_���AĄP�XvM�m�ʈ���>*���r0�ْ)��]�~1�?����N�D���p9���(+�a���.5%6^��du�w�	��4�>�	UuV���?�r��KR��,1�5zjA���$Q�*C��x���@z݄�ͦ﷬8p'�5*��*K�H��!l�2N@13*{p�:��f�RǮ�\���d��U1bw�ujq�R�ʜT���@hV��X�(p�g�}��襒<���:
نB�]�������=�eE��ڔ@16��M�xH��OO�津\���π��4��fg%e�=���@^���I����o��	�D�%o��X�4p���#ty%?-uoM��i��[��Gv�p(#�TC<��S؄�%A�u�����n��G*�5e�K���DH��(��-շݚ;
D��2Ky�^�[�2����Z����&#��{N�a҅)ށO!Wʱ)��Io��sR�W�i:�aȪ'O#�j���o44Jn<`���F�:�9��YP�d�m��f��cl�M�����_��:3�Y��L��*Y�7fP�x� S\�`,E�6�M>��� � !(�5!��Tr#n���W�f0���"~yM#� ��ȵ+��^�?�}��^{��g���6���S^����K�(��&�^^ex�]�A2|�
-� @:�/��a9s?�����_�q^�.�6�H	�+ﰸ!�����2(c,�
����xx�2q4�'e���W��,�}����`rCP=K��E��O*cf}����R_�?�WH��i�#�,uU�����T���-C��Y��<�N�:ʅ���u��h��CZ>��*�����V�;D)LI��3	O�)x�,Y�|� Q$�RY=�̰�2$�=�Z�Y�أ���n�7*g"�����������"u�ݘW��ѓ�\�6�U��c�_M]D�	�˺�򽘞~���ڍ���3V�̊�pu^m2i�t
yRd�
��S�4����?�ו����h��9J; v 7EF� �NeR�E+IL	�d^37��?$M<�큂t�BY���@���[��V��L���ec;n��lE���5�W rE�c�ӍF�z���<x�@&$��(��\�����S=ڱ�����O9�w�(�D;��e�$�Ne�ʎL�v��3T��Z��)�~���cs�4�E��)g�����-s��j�mb��pt.�zlQӷ � � ��������پﾨ�s[@���vFb�}��e�s�"d�UJ���S��F0@�����&���g����P}"|�C}O�(��ϗ�n8O��x^@Z�{c�� 4a4-S��[v�Wa}�x�4y�ix����-rhr)��;��y3e���1�0p������/��� 9F�oVfm�S�u�*��3��m��Zz<���y�t������lzy�� 	nlY��y�t�˨`��'��O�K�㦱EM����??չ��y�"��/L��q�=�_$E�Ɠ�!�%������r©}�ϛZ���H�-8˹�abc�\YKx���
�8�G�,�n=ix�F��	zV�g.g�/�7oyb�b^����$m	t`Sa���&M.��[�a�;�"|;W%j��!>�q*���K�cYV�+]]���d"X�<�S罌۷��l\|�#��mx9���tA�iI�xS�@������l,�I�7y�P�#8����\�Ŀ��l��7�p5�I�V��Gh�NO�ѧlAE��+t� ���;��zF<p�
G ,���J#~�^����M�7��/wŀu�
EI�a��k�˞��?{`�#�q>I�?�*�4�}�[m�p@6����i��8Cu�E��,W���ԫV�Xl�lM5�g�'z&�Ω@�t�"=sQg�:��gg%��2N�,��}b��b&T*w�8,Ǜp�=8�\q����Q��c���{�r��p��̤eH���L�RȏN���z-����@Fr��,��_�7����-���K�m��[�'�ȗ����&g(S����`왷�%Y�!Z�W��N-����ŧ&�Q��ɬӴ��B�n��4���#��"0�F�*�m9d����r7�ʸ����#cΐ_0j���q�mZl�ߒ�#.O����`��l��o1�SS���S%�=6	/���l�9?�2� ������
+�MW��67�)y�M����Ȗ'.����Cw��I�,�(���P�.�ڮ����I��U��y�2�iQ�D*��9KL2Ti�jY�x�ą�x�6�	�o���~r�'	S2"n)w�t4��܇�fTD#~��rPC|GQ�cѿF瘹1܋ʼ��z��/�F�.�n�Eu�)Kݪ*�%�9�P�G�|U�3W�0� 1��x1�cm���bb�%d��,��$a=	�bz�cT�pWh�J0Ӄ<���l,D�·��Jg���a��d��������(�p��eAx�<p���{�ា����[g�`5nTF�Nv/�H
U`�o<�p�TI�NX�a�p1�D�����l]�ɕC���q梴]�MA\ƏB �G�U�*��������j�VĞ)��f+�D(F a~�*z_�8D>Cj9{���C�c���zc�j��7x��r_�!2�8C�vO!�n����O���z
ѵ&�J��y�x��7�=,Z�+�zU��bߡ��q���B�ͧXC:�
T˭)�-�L��ڀ��e��!#�@U_{o�RUG���?}>S/Y֔�xщ��`!�zի�|g(����m!�*W����mH��rʲ��]��#ve��ay��.ڈ��*��E�8d4ZY8e�������jD����ڌ"�Rz���F
�a�¡9V��Oc
�}�Bl�Aݦ1�a<h�������/Q�qU(���)wi ���ל"$����i�Q4�6j��lG�X�!�>L� ��Q��{��ZnB����DY-jŲ��!�"Y��	��ry�j�t-�t��IF�	w�Y� �ۄZM���d��yZW��	�٦����Lxkj��c	B���hpJ���-����t��		+~�3�S�e��#�k��+��J��V����é�ݼ���% mK���.؃�����Gdǝ�
;�8܇�����ԙ�PC�P� 2�����$��U�f����f[U 3�(
���!C	����y+��[?7�Tш4n2~h�RJ'�Y_����jⵊpr�}];��HGT�݁.M�hd�n�U+�#F���!��	�l���z@�9��b�7Z4����6������-1K���r���P{iG��L|�xw��>��$���v�6���Tz��b���zc�m	���40:�����*���tĆ���$�z�e;�S�u���\��ڌL��t�el�۳Nf��d�y2k����e)����i5J��Z.���|4��^M�7�p�۲��-b0��>�$���Jqj�ˡ,ϔ�*� ���,�O�`c����ո7�}f5�WXo�Z� �N�X�u�d��a̧���B��]��{��Q��m��I�3/2JN�s�n�'�!����E��<u�r��)9�0Nx�+jM�p�{���;�|?*2N� ����������Ӝ5���OmW���n�n��������B$EF�g�5�)��^}%�����)z���m��d]�dRMĥ�b��2Ea��k��Bf�^�X�z�k��r�����;&��Yӌ��#�D9o�M4���hֳ��җPR6ݡ ,�j,r*��pÙ�^E��p���s�j�W,�k�z,4fS�]��)�U�N4���&l
8�Po�0��]��QP�Η<!N*�k�����W�{�,�vC#4�p��N̀D�U��c�)�4b<��X�1�s��M:H7�28&��<�2Ć_����K�t:��@J��^{3A��Ѱ��m<����eś�A��t/�P
:��Y�l��/��yPB�6)�4"FX+R�����\8��cY(�@������o��y��^P�M�eHY��¼� �!�."qu���-Oכ6�/������V��F��>8�<Z;yE�xަ�(�xS����"�=�Y6:%]���7}/JJk.�@���S�� u��`+�y��|S�3mZǡ��|��NA�� ���Q����6�Nv�S�@.o��F���F4�[�o4��Z�O4\���uH��pr���n�����h�M �0�+^)��8��'��M�2N6
c�#��8l��Mw$��l+d�Z�x��+q�4�;�o��CN�����ؾpV8��9�\����:z�X��i��ua4Ә^[?H?��y\���P�_kЉ���-�8w���U�"z���A}�@����[�f-����p����lԃ�wB�,ݙ,N�h��:�"{p|D��+�Z	sF�Z�]��_���<��2lQ��ai9�Je�f&�d���;e1׊��&,����*v1q����V�Y0<&������v�,]?b^���ʁ��t�_�D@�7����8m��7	d;�5ėo�(�X>���v�Yշj����EV�j?|| �W�Y,芵JT/Hx��|N�6�f}+�6^�?��Bqr�?N����l�7j����e"���%��7�Y��< �I6�A��Hh�l��ȵ׸�|�4�}���xߧ)� �����,(l^���x�oTL��|����j�n
�g[?H�5��'�����<��_��Һ`p����0zO�V�� ߪs*AS(@�.&�ú�&GK�8e�F�h�j��ގ���tG/7-x�%�D=���3"-�Ƭ?�����3����)�V�1$(/1j=D)�ю�}V�^�9r�8��lQ�U�x��Z�d%�
֘���~Vi��m@ ���PcE	�9&H}��=D�j�S�U4�]�5���&��-G��"�"b��-�E�5��z�\"[�=� ����/P������c�ja�*�=Y���C��h	�x\�H'L�摢_�UV]��J�����0��4V�	�w��[|v@éU7�.����փv�U�ӭ��\����7!S����T��y='���Ļ�F���O�*G�ʠ���S�Y�\(\�c�+b�z5]�d��us`�lVWҬR2�6w����&�I��V�[J����z9!��Ⱥ�\�bbks��%��c�����ϔǷ��X*����+��y}�B`{�rP�o�Y*��b�}\ 0�	�����/d{�����o��cG�Q^�K�NFu1۞���N�D%��Z�:��C-�t�.u-"����|�{c6��RdT2#y��k��9f�jg0��V7��Q���G��4�o���Xr$�_OY!�3g9p��qsL���k�/:���agi�I��yz �"����D�t�~�8L��F)}r�Pl<ǅ�q���&c���X�	S�~��@b}s��r�P���Ù��j9��n"�Ug�ۺD\XĤ�T�B}/@[،��]r�������NZB�x�O�0�m��|����-E�*=��q|R�	�b���v���bG�:��S(�_)���*�d���Q�ދb����x����*1V��{_��:�<ђ'I�>�b0�[���@���� �Q��O�;�k�ϭ�8��6�B�-'�L��>o�����E�'L�������&_y3U�V�*2���X`� +�>m`eraWк�������لY}�j�K���B�%xv&�!��5�Q�y�o��KAw�Ε����e���N�� *�4�������rm�����gl����6?��Bf"�V�����?��JLD�Rvv?��I��8�T��W�L�|ھ^y0sH�*�Z����-����mI�jgq�i���T�4.�G�>��(�`���*�
�D�\��rЖA��O�v�M$4/�v��8�Nf��x���k]�}����� ���r^D_��Ғ�ʋ��5(��?���<=�4� ��<̘D]��Bg�)C�L, ~�� �<$J��1y����au ��J����R��:i��R�����!��5�6K�mH��!�8�S��_H!X�'���DÎX�|H�hJ���Gͫ��-��h���%8�M�w
V)�u�_����5���NW';���ia�ZɃ��V��֞ί[�n5��H���?����[���\��Q�ͽj��҅��һG|��������F�'�U��f����⒧��n/�c�[�ۦ@Ƀjγ0F�
�&��;4����5Y}p$@�xΞ�_Ϙ��w��N����ICr�(&1�����,�L��S��@{zFP�۳�ĵ
ԫٸ��d�m���#�0�ť��?]�vS�s�@����Q��`*�g��6�L=�q�����	� �j�f`�b��ʂ�S�14��9��9�X{���ϼ��j�+�4в�$Zł~�0I�E�����;��φXm����]�a�K�rm[��R�)oC��Pw�t�ך=��,�=6��}���~��(�&�v� �/�3μ���`�[���c�j�ykyWs�S�Au��|�#Z��P���J�u��<\�]�� ��B����-���Lre��խ���0�p��JN��l�5�h��u�- b7��֤������I���d����:o�-��:�mO�!���:�Et�䶖�Ѩm�G`�4W�VE>�t�����,���*�&�#Xk;U��M��N?���|��RIlQ:��x��l�d�kҐ"0���?�� e�i��z(�]n�EQ���5��)�񽩫��T_�W^k���{ޥ��9��3����6�v�4����i�E+����W��FO��p�_�4���=u9�
�S��i�m,I�Ba|C+>�i�t�i,��Q��	�ŨR)�)�!ؔ*�Q��\�޸�73p�G)��]!�&[�@�D���L�L�a��$-W��f�Y1!���Ii0{MɂR}�ra<B��
wU��6��Ur�`�֐/������j���Yt�8���^>	��W�7�i�qjI&�����m�S�V��Ê��W��Ȓ:�_U;����z\�w�^u��	Z}��o�Z�KoX��E��+��a�nx�-6 �	0h
�@� R6[t�ʐ��}Ӡ����.�<���1���>z�O���Iޖ�{�� ��T'y��E^��V1�[�'��;"tl�xg��[����)�W�>�?�2�<f���ƕW��[�x�΢3WCNZ���g=��~����;��q��jG��nڶ����ip���Z�̧c���,��<��3�Z;�,��*����(�0�]�'sDTϫ�d `��^Io���:��s*ђ�6����=�e�Q���:/�?°��{��[�#E`q�I�@x���N�b��ʦ/��(S"G���T�@3��r�P�6���w���I$�e�0�#��jԫr8�n���U�y�K�Ҁj�����M����Č�����������iAg#�as�+®>^�,nk��@}���P�b.e�U%I(\=�^�"�+��"�����0��3a�� /�X�	zC	 �x�᠓��.K\aJ�덅Vn�N~���Y�}��i3�����!�Ӓ��˲��`8��)pPn��P�d����h������~`= ������uok�ᐶX@��*��NhcW����5w�57V>�C�Q�bR�B��.�JA������sލ�خ��% ~�6\nJ��7��/q��� �.S��U������rrr�wj�p�F�жOI��N��s�XxW�
-yU�Zw�pO��R9�Ĩf����&��{�3)��"\��ԢG<�m&���8K~����M��j�n��螤΅��w)���&��������0-�yt'[���|DHc��_�`a��K��b_q����]�E�	�EdY�u�w(u"�{�����[dc�������G���X�(R*Ҝ�{Hs�g^'΋2�~v�*I�͜����W��iO�E93\A�N�q e�W~�������¸�,H2l3z�]"��+��bK���?h43���V����<=W+�|Hpe�)B�sR����g�@嚎|;؊��������~]|�ņ�9�|"CSu��Rh�2��h��o�hű�����B�G�f=מ�6Q���}�n.����C�X���R�a)"%/�9Z5����Ox1[	6�2y�2O�kbQ�A�Z���I��xiv�#V�>�^���jJ�C�Hx�8}��K�Sh��|"��.�>J@�s�*�`�0F�[@m��V*�s����T�Y�4aQ*V�-��5����u��
Lhr
	��f1��ú�w��~�J¢�����%�<մY2����醸���}���{1eV¨�����t�_�o-uś���2�Bj<�a���sA��r�B�aNd�ʷǏ����}'Μ���<��s�7��A�<�ʽ�<�0�l#�����A&���峉�Ly�)�lHPV.�P���U[0��8�f��.�]_N��̠��
'����ܢ�*m�qx�0_v�sk�֛��^��ە��ֳs�S<i�z�AG����*p�!����j�5/���6�C+�*|x��a�7'����F5d���2Un�wفi����+Ǳ�w)��j�p�;A���qY`�:��;��EZ(��
;R�DS5��;�|��!�Y.;-�g��0�^�3���7�{���M����C�L��L��y�C?�0EE%~g�~K��]��f�"����Ἲ�!S�ڙP��0�[P&g��1��ڈߵ�Q>J_��m��FK�#��1��H�ۃ6�9'�O��`�4p��z�1�%3�����K�����3�G�	�!�pa&�}�'�^��:��?��+]Q�bUeF�w�'(!�x��d[��Ʌ1�Cld)��發��;�)�ǯG��P\�⾜�V�z�����mJ��}�][�y�A�Dτ�jouI2
(��,P�2��АBcF�^:b
x��Ӡ�ՒhѾ����
n�37L�@!���~z[� ��W�6DK[i.$ǖ�n�1rr-�= ��{�P�N~��V=WNt�{\F�
���q�ǒ�ci��^%�)��1���&#�<�G�8��/*`�m<�U����N ��oȳ����ۢ��df�T�	�6�$cMvL�' �nɭ2�/��� �ĥ���"gLa�>Rz�̒r/���>���s�ol"���������>G�S��hQ_�Ť�kNl��Ʉ�=���n�9�c yl��g��u����rXI��l�x��K�l����\)�# �N$���/zwc�_�_���6Q�I�u����#ak��GCj�*��z�Yɥ[��Ј)j@��� �Z~�Ya��l�SwL$n@x~��DU�ȄNu<��\��8���$�ŕ��"i7?��;�턲�&OV�'��`g(���@��7:+E��#�8c���E��Q��
_��'v�Et�c���g3em��h���?֌�D���f�k�3�(q<��ޞ���S�����hP��\�dQ�L�^Rǯ9� ��7��Yd��̀F�t�o����`�m�t���a��C_d�4���]����k�F�N��1u��,H��h�F�x��@eo���~9e�, �l	h�uD���8�]��i�-�;5\�IȺ������<�m R����٧2��цo�]�}J�Gr'gB�d��Px�hL��Y�Tm1��h�f���K�� �.K��խ�Tkw��X[I�j�5#/��F_�*�g���ƽ(�\; |&.2��iV@���}+�T`7wʇ���(��"�dݗ�W��
G��+��������հ9S��D���;����-�����2�7t������F��SȳD��*��Y�B*� B.��d��G
��W��@�8 �Ӥ9��NK�6��<�+#��>�3�ͮQ��RF����0�Q�L��.����{_�G_B�s�[Zz\������q�U�%�9���=.�E���C��V�(�^7�b3���I'ԝt��+�� "�,	�z � �:i�囐>ۜ""���TZȡ&�C^Km9���q�
]|��o���c��k�mQ��w#b5�̨��p�5m���W�t������S���E��M_��#�T��Ⱦ��x[x�{fc{�Xplӕ],�%p�TC�񷬿<����$�4��`��d4�$�iI�l��x���tz���dw.k��T��ۙ����j����Z� �h�����(n/=��D����)�/��& �4Gf�l�U{q��2-��ǎ��O��#����"
�#u��(z������(EKUkU�5_@�h�+Ǧۦ������z��]#=���u�Խ��ı�愳4l ����E?����ߜn �Aejݜ`��9���o��{m�]T�Y��l��F��N�����Ģ��
Rk8ֳ^�O?��qH���� Zc�<8�i��<����q���<�}ۂ*���塛�1[�Hhv�:�L��]�6����o��c�F9�}6-I'��h9���M*�V�{��xB���.�M�R����t��"��yU�x��7=|,�#�>���JT���0̐�sr� D�B��=��{1���^FwRt�n}e��iAE�]�[�M�+�U�1(�f�,S3��]� O���u��O�ϸ7� �E��+0�Ԍ�߾�B�����N�,�,)�~sw,�ߣOS%�N*��7&lL��\�׼�A�h��L�1J�����:�/SE��AD˶����ޜ�G�WWnX�k�(n��o�\2[a����E�ẅU^í�:���zpM����[n��QCXD֢|sb�k�oC��&���,���?W2�ͱ���=�y��D-�9�_%I:��\K��F�4=�K"c&�n�9L�z�=oD_���Q 3�׶�Lr(�;Q\�`�j��2�F�3�5Vg��xeړ+iفׄ�ӈ�q�-�-�ޫ�\���韤�)�:S|�{��PE9�O��fNĖN���;�\�V���^���/�����Z��E�D��|�MPo+Ѳ����p��RT'����ő௔�����!�m~���r���D��:h��m��$�K��6]ҥ`���m�愹���c��T���lf�$ψΟ2_K�Ăe����x���pȈ��=ԡ�+��j:|�-%J��F��d����s���ݾV�ϟ������B°Q��x�,WC��Z>�����O��W��J���<sY:���۩�?=�/����Mv"O�����fpw333e�Oŉ}��`Zi�"�����/��mE�{	#��:����k�*o�htc,��gZ����r�NކtL!�O�ϰrlWV6Q��"�T1`�W�,��`B5a�sc�o~Tm�O15�{P;�u���:����l�pǹ5C��e�K+\]4�{j��w+���K�K�k�гx�|��OiؔE��o�m}��/9ۍ��ف��Ϝ���5����hdkJ� Q.-�b$�BHN��g�y��/:�����{I������;��B�B3&c���)0�tЖ"��|1<l�8a��΋�Z���0�Y8��Sx��1�LtĒ�h�_f�3�:2Q4]����?N�vc�ʊq�0�C/DH�m�]Lkn2��4���A^B�C: ~vȻ5��$�U^�@�ı��:5�6��>/t���Z0�c�Ǉi</������j��Og�$z��t��Oc��}_r��a��oM�.�3J�L�~�:Μj;%I�W~i���6-ZADt��\`G=�/n[����k��*"��~��e�0'x$:w��6A7�q'y6g�u9������"q��m�o�F�
}�Y`3���l;ਘ�fՔ��c��a�2�J�p��.����j��>r�����	J��B?J�質@M|%�Č4��o�=�W�?g�Apu��ZV�Vu�QW�B�M2ϪVA�_���^d<�=;��>�B%������?k����pܰծ�ߐ��R��'x2Ö�z�q�@Gq-�V�my�w;��Z)2_fN�oK���B2��g�_y�E�:��ug쩚��	�`�m�0"��Z���wrq���n���#��I0���})��ش����5~h�T����	�gM�|�;���;�}��S�,^����N�%צ�^ă����i����@�a��:W�PMO�LAm��^�r�a��خ���⧤�G5 }LB_`�^�1f�-���� A��pp�SQ$ǘ���R^����{��m�V��.���������*w9b�S!&r����6;}/�<F�N�X=K�O|w����#.9�&�݊J������w�d=B@�knLW"P�0��7���J�k�8��t
_�
�/m�/�����/��УMy�ut�k�D �*�F��U3��5��X��hN�j�u������#K@�sOP�q�|6��+��z�x�;M��m�o�?�N�Rz�����ߏ�8<�=n��ly���h�.�nU=L���=�Lf��a+_9�=������ܾ���5�5�j�I��aY�Z�3Oi�-�'����rXէ���p;
^���3����?�yX�i=y������iL���Dhs��8����Ҵ�o����뺁��H��	s��i`���d��zR�o]z�t�~FȔ�*�W-��{�����R�OW"Q��}��8�Y�α�����ύ���0�c�+)r��[�6Z#{d4��k�U�N�ѥ_]�m=Bda>�u�z�UH `n"kB�,��pDl*m�U���|�q]���}�5,Z))�6c�=|^���jI�{@Or�2���#�;��3�Z��rb�
��
8�ü��Н0p�#�*�A�ǉ�:�a�a{}O��%je�� s���ߧ�"P�Zn�_�b�������!��-���b��������]��
k�g�+����6�hTm	c�A��j�1�&�kn9W��]
?���X�:x����	�ڎ�^�|醟c�[D!訪>OX���F�@��좞��;G�`��
�Ś3�F�\�N�'�~�N�.����Z̽襒��cbؖ�j񬫠�Kc�U�G[��^'��C(m� �~s���b�篞!+��|[��kI�ڒ.Q:�$r��oL�����S�<��$�y0]~QL-既�7'�I4S���U�=�K=W���?���Qg��x�J�7�v��]$t�		v� f�{'?Qz\��{�ܛQ�`�G����H��Z�Z�FX��
B�in��� Տ��	:xG��s�L�3*̬Qs��)�f��_� �$�O�B�BښVpӿG�/ ��5���-� ���
hO��(��R��3��9p��bӴ]nl>-�f����뻧N�RD�,R���|k�
��7M���߫�� �%�S9��m4��/�xp�����酓�ktM�A&�|�~�;D�'u���uZԑ	���#�f|���jw�BZ,�Q��� ��D�3�@��9�"�k�$��� T�w�#:��X� B�|%Ud@�(�	��UZ�ҩn������t�Hno�
Z���+�ш��́�^ųҰ�<'ҝDG�z!fC������B�U=����jFN����Q��k�׀��Ƿ�L���,��� ��tc�Z�v�=J��\�䵂B�&⏕!M�c�����Ɯ��F�֯;��VX'ȿ��f�>�ʴڠ$ ��J��d�%w40&�����J��=@�}�&C���d��eܮ������Ǿ����|�2��[������O�6 ���=膌��NS(�mA V�a$�⯃�f4N�,�H t�wŦ5��#s���/��q�қ^���$
��f�b]2!*O���Ї�FJOt;pȦ��}��O-O��7}����-W�� �-l�D*;�c��WL��$�Q_���*q?��y� ����j�l��4)5�CK��
 �B]���I052��� �=�jc�f�]���ZHD�(�����@C4�^�t��*�)��9x�4����>x0/fOX;��x0�YY*6V��>����U�8��Z9���~��ߺv
�z�,,!�t��M���6F����G �
�v��+�|;L�N ,Aύ'�	��,��/��E��������\_��0�J���:�1[ලI�����wx��u�S���,�8�E��.t����D���~�C^^Y��b����L��p���0ˇ/a�5��at>��uxs`c�����5Ö�ZeKa~����:\���"O-�V�p�����_���_F:�/�`�]��_*;)�����;]���7�:�7�<���3]���F(��X�-�f^�ץ�}�� 謰�����p��٧Ͼ�#��� FV�Ǯ#��C����]Y$�&�9,ǹ�QAѻ��[��"����1ZO0���/Np  ��Ց�Xb�	�I�t��nʹ��y>����O	l8C�!�lo��4wT]���5�M�0�A���4�<��9'������(�Iri�����1Z�W�潽NhD}D{���2�H�pc���8k�3��3
��4G�qJ��gK��1~�iS��mێ�{�)Va����@��0�)T�X�� J`��I@��i�����l�q�[�|�:��u���=c��1�Y(_�D��2��O¸��P�ri!��M?�n�+��V	w���b�G�[W�ð�ׁzvW9�@['�K�C� ?	Q,�����YNC�,��7s[W��oUH1v:mdcZ۳!T
�pi����$�����@��c�s(�W�^ �i�eU�����N]X/F�$��z����g�l@H�$]���;H�O F6vI�%���X챆�-0`���gִ�{A���(��Z᮵��G�Z�ٺ��7� �j�Z�N�D�-ņxY�"+�q�m+�Fq���y��"`��DK=t*d�z��d[΂�bIE�p�~Һ�3�R�I���I�I@U~|���)�N W�#c8�5Y.Ԗ�S����|��ұ��R���SA4�L�r8�ѮT��W�5�̻OɁ!TQHak$8�9� �y�ܕ�Ar���$[���-������zNd���ӵN��m��L�����dӇd����t���,y@�b����#4O�~��c�
uv0/I��d����H�Gi4̛dʤ~#(g�B�ٴ���N�/�����lɇ���UT�!0:} ��	fW0|�.���4��u����7ygO��K�%���N�e�g���4f}��?]U<I$��ʻ����G�p�*�A����w���c�);t�`d[fͪH�i�q�T#�i�H�L���ވo�h�4��R�Of%�yR�أb�Pi?�l_��7�s�h�Z�.���԰�T=�)�-�k�]M`X��ʶ]::<l�z2^�Y^�2�m�p��&��B�*�����v�Კ����ڧJg�<R&��>q]�p�B3;n�Q�%&Gq���B�_RH����Hƨ`_OV�)ͳѶ���*fc�����y��O�wN���(n5�n�4�~5g�H�4�ۨ�G�'�R�Vً}�[_��e{�n�o�se�	sK�7�\�)ǭ@��D+�k���W��	�zS����II�hy�t���{Q�IO��v����2x}3Ɔ������ٕٗ��ɪ�m�B_�ׁJ��<3o����c$��.ΝB�,��^�B�OS'�^W��D�+�M$������vQ������O�֡��H�UL.5�����c��B��^��٩?O��݌ֆ�vqH���2�c,��["�œk�m7��/��E��	]�h�ϊk�#�bg���My��e�] o�{�oB�1�.�;�gs��ݔ$�nCc�Tj+�`.���S�p)�lI^�ӽ�R�3Y^�&�/�5��F2<%E��~�����E6� Eb{4�0ȷ���Y�/�d���0�0a�~tF���[��P��F�0���ޤ�
���t���R��G�wOn#j,@�rs����V]f�ws8�,��6��ud�gv���t�f��f�"}�&�uÂ��a�K�W�(��yfT�����,/q�⭤���?]���(,��S2m�TO�׵�m�h-+)\�0ݽ0�/J�$����V��K��}�,VFx�]�~�o끰�Su�8��q��UQ��0��Ġn�s��p��,/;�2��SBމ%}�u�����?�NA�m,�^����:�z��O
�~���ד�x�����eRpci�U�W�8̇��L1���Y�<�p�λ���A�p"{X�w�@� 	���*(�NW'V��/�~�`a�������~�����8��W���^�Ԩ�@��V�
���F���aP�4S�V�1ψ�:�B��!2���ED����9�̸з��)�z���q�V �F�J]#By���*e�F���JK�#�̠�-��6�z�~q/�����/_ޭ���	�����J�K�d3�ΫZ��=3��k�գt��0���($�#"B�̡��	����a�4�I'eY0	eR�K��A�9�>4�l.��_'�7������9.��u�U�����B@�3ԗ�m� �2�~{_�;[�7�������ou��?��>_)]����G��,������Ou�@��0[ ��AK���z�9�O^T+X"�E;�V�-Ú�Z/9�I�/�u��>���,j����U����8%��;���*m�A� G#���oeT���𖞩��^�*:��|HO9�*4,����b=��b�?�K����f��{I4\�>�~>G�G;D����z�\J�Q/�
`ا�����J��j�tV�-�W���-��Y��-^�u3O9{zk�b|.H�8[�Vy���]s�S�U�rķ9oj�&Td|���cJ�%���K���Q��1Z����c]�!n|%Q�X7M�V�6X�7��:�G�K&y�ri� �"h8�J��|�2�7��A��[���S$Eֲɐ�έꝥQ4
�|YL���-�ƆJ��C�{�Z�BA�ɪ��
��_�4��a�h����D_e�06�|M�a�W�Gs�"VȘ3/�fЊ����J<�W��R��Zm̘��y�l͠#UE5�+p�~�t΋��<;�ªhK� S!(u�K)�R�WC��޸�R�6(�"ܳ�#s�>�z�E`�l.����eV���,��yS�R�������*���˛�?}�� �-2H�ᳮL˝�Y��=�<��4��e�K���jV��94�Z����4c�~�uvKݹm���?8p���XW��!�$`$t	��Q��-O?���W�����O�%���DT�qm�����&e!&�:ĉa�Q�{!�����]J>�L#u����t��R����E���G����V���L�.}����ĵyⵋ�[��t倭��h�D�q��MFIqya�
Qך$z�Yq�#o��78�M�z&��[�S+��GJq�f��g������J��Bs�N�Oه"���͒�o�:N4�i�*u�3v��,>C!�4�G}�h/qw��h�Մ%9eu�s:�c�t�p��+�� ���
�y0-K�������7����i��bK�qRnO����.�jS�W	m�_���0��x��#d�q��8�i|�Ew�퀠���PVX����2�j���3 �����ثs��Yk�*�Zm�`��ԋwj0F�d����(����貀´����k���5٨�)&�;��r6#�|�j*W��(�ٺO��h�ŹFS����1k�%a�'ѢC
��NR�z�9�.c6@S�U��c���yUqT����9������Uµ��L��+{�<<���˟��^5>	���w�H�_��Ǔ޼F�X�a�/$�ֻ���4xv�+8f�j��E�Se��C�4�WJ���Kwͧ���l67���Sxj��oѰ	c�\뻽�:"N�.V��G7z�:h�4 �Q��xs|؟{���s(m���9����Fv�"} Q�WÅ�÷���w�<��li���#z���C�3p1����~��c�{x�1�/��$8�x���X��Y���op�벦���j��Ki���"�Aq_#IFa�;�{v�A�h�dr0����Q��|��=$��bvF��#��G���()��C�z��E/< G2�`����H�E<�������nO��_E{\�aHS{��@���,k���1�]���A���Bg�dB�u	b| A��5�ŉgp'��)�S�f0e�b�������+�B5-�4Ħ8pm�]����E�5*��Ӭa��T��q��6��I�b.ʶ���\$��'J�ar�~Y��bT�+/��&���Yġ�I�n,�of5(�`3%�h�������-�MLR�0u�$v9.ʹ�n<���M�A)Y?BuX�,��c�HOH�w�Fs��$¦yK��6!����qU���%~7¤�Ȁ\��B�@E���n�a1yڠq.��g��Ā ����,������k�F@�Ҵ��z+�9�pM����>GI
K����{2����ַ{p��H�o���Y�{����F��2͙�D��^�q����J(�ٌ�({�	��i��H;~�wۃΙ�,ߟ�t1�*R�B�m��(���dK&��>�"9-�Fҽ^k��T�OT����H}�!���0`�sff��8L���p��Dz�&ĘY�2>%ŕVx�[ݩ�#����=�
���$f�t�]z�@�YB\W��R}���<� ���U~ЁtO7`p�Ƒi�#���9���~P�D��Z,%��@�M��t���;x~�DC��-{ć�lM̛�z�М����J4R*�ؕ�����p|�Rܩ�r1�������bs�{lr�Rz���BR�=�����W�}-=��%XYB�l ��ɲ���\��������+��$hg��4�E)W�m1���q�S�2C�����a�Gs.�@��`���׬L��⽸��^���!�Kx=������Y�5���g׀KM�y��\)�����M��^#W�M�4�/gNq�h���O`�/Ԅo�T��%ڄ�k�2���������6��泔[B�;�����y��$���n���p�S툫�p��-zP'ݫ&�0!�6� ��%����l-F���E�Y�PJ�`�@]�9���@0�U@Ǻ����(���HP�i���%�to���%o�D�n���¥&�'�N��a25�E}�U�j\#����A3F���sr��l�����{�_r�Lr�`}Y�/ұ�rdɦ�D4\�|e�Kj���҈�����p�W��+���t$hE���@�pz���BcR���(8� �
��o��N_�҂C�
��m������T���24�i<����᧜Y��T!�|~�����Ƥ�*�L�ƮԞ���˸%G��?����oϜ���@r����YT���S@�b�!����Q1V�Q4��SXN%�ޡ�0�X%B1��Kv��[��6t�F��|< I��8�K�����f����J)G��v]�WK|�
K�e͢� �U��EO���R˖����X���߷ Y�m��Pޘo���E��>�#�6�G=�����!S���R��0����9�	�&�Q��N'&��Z�Yj��ۊ�q��v���o�5Tɛ"#3zd���1�C��M����Aj�#=����Qs*�K˲�bU�wb� A�2��Iw�zA��T=�Q�H����Cn���=�Ŝ���n☾(��;�- �G9�[�����l�	�^7Pm!�G��_��4�`�5�����@W���l���y�f��^T���K��Gv��ԩ�&r�p�#p+��5��1�Nu�8�yܽ�F4�Z��!�p6�Hkw[���b�3��{k#e�Wvg$q�B��yw�>
����eG�2�n� ��l��� ����3� ȓx����-hr��<i.֊��\ :"ĥ����KQb��j�Q���4��R��u������o/�|�\��k|^�P`�m̙kz���:��L����ri���_*9<rN,��%����*�<�پgʣ^�k\&��;2����v5�-%;;u1�։."���������䆬v9*�l��"^̕\VCٍ΃�	zfQ5@9�Pe�)�ݟ
�5��Zm.B�v����=��+C�r�?��K{���tT�R�N�?ъBR���p#�UԼ;�ml���R�
�(	(�B%�-���'�R+�}(gCɉy��b!����{�ovDZ�G�l=�"L��#�H��j���:�p$`I�16��՜P?~{���"���=,}�2����Ʌ��2�aVae�n�����a�q�\3��F�0����l`l�8��=G7��Jk]�>1��X�[}�i�R���S�V�;�4)�|���Ԉe-J+�����:)��W0���-�f����V�8�����,�眕�@���X��NP�^�L�R�8�)>�Y�����tm��3��#3U���>Y�������ɞU�'-\p��.�@9����fC�w�˃���_͎͗2h��'�#v^|V� �9�*�ȪK�x�;u�T}X�tCs[\z������s�KT)f�Y�e[V�xp���#�퀃>��C�����m��Ey����n��\�4̜IV��햾b�I�t���	ss
^ �7�:�=`����20&�]C�N��y�I�	�<�29	�����Y��7�%.
���JW��4]��,w �M_s�d��#h���'�e:1�"L�A�Ӣ���ҹ�>R�Cs���g�Z�w#���F���q��.�����a`/�5|\(}��-Ox�`H��31����w�B
ntp�c��y�G�4�.��)�+��`]w���ÈT:��:��`��4��#�*�B�4��AѼ�0}`v�*�}���N�?���M��s��np4�TJ��Fa�A� ��)�T�"��0�m;��J��ˍ8���2�o��	�� �GДa���Y�vX��O����?��֨�'����e�^w�t���
�2TCG�r���)M��Je�cg�H=i������&��!��V*��6��,a�%ӭ�M�3��� ����E�+X=Yb_N��A�_.2����Ok�e֑8YH{Ehnq�L|@s��DŗR�Vp������8��,P����a�%R�PTT�Ǹd.'U��lْ�ow~��c����O��c�o�\N��K��h���4w,���Y�f�<��Dq�LSm�)���Bp ��Py�M�ۿ+xM�M�6cb �e[@��BU�p�g��R1t��8vq�������r2�܂	%�:-O0��4,P`�,�P4����d&@��v89i��1I�a.�P�%/u2��)L��&RE(����rgBK̮�PP�(��6R�_l����~����-�L�g�gs�~dX���S�"_�nW:��&��F[�양:P	���hd<G��Q���3���*$���j��թoi}��m�NAP�3���v3#���5��"m�v����vM:��f���X����?����2ߢ�d�0�-T������������2�.� ?{?�� *��������:7X����
�l����A������ze��z�@����~?L��o'1"��7�����#�Dq��c�פa��ؒt����NR��Ӿ�K��@�:�� !�5�*!�6�/2��IElp\z�{?�?�g�M_�"�Xb����a�9�y"�%=�����t�2U
�ۓ�����zye��lm����-[=�����D�?��C�	�v�WP�TҼ:I$�ؼ��"���J:�<{��]��V��������6���>�L�J�N�WlR��G��Ѥ���[TIp��Tv��B�U�)��1�	z�bIDv:	9�ʅ+US6w3z9^��K�1��6G�,�%l���xY���T?�*It�z�I֎o'�/ ��1)�E՘��a�G�n�䊟�7i���(�� d�aF��9]�4F����0�}U��uT�9^�����ȷ���_�T1/o8>36'�a4E�p�TG򛨤�v7OI�j#r(��X�8����2foS����u���ܥ�"�tW%rg�ejJ���	7)����a�k�;S�,�?�ɘ�>�+���>�]��2��}��ݳ_'���ug_9:j��I�3]�F��;8���kG�mDRQ�˯[�8���E�ݼi�ѷ�p�)��oq?밼�
���� ��h���vB��X�VQ�3�ŉ�}�s>���C���a���a���}G���<��ē�cbV����r3�A\�J1��Z.c�fJ��@`��<�Y%�wѠ�tށ������xy��+��X�
�`�i�N
�`;�g0{[�A��"�W��U��#r�v�a�����Y]�V����K����31��i��66��%N��[^{_��y�E��9���f�mF-l��I�q��(1"��3�U2���k�[�ث���-�&[L]_�z��
m@���n��W		2�gLIi{&�|2���HeU�Li3���t�3� ���Ss�9cҥt �Hꐚ��~�*�*��q\��)"���g�FY������Jzˡ�'�J�\/�۠:�F,�B_���(�=�c���=�ҋSk/���` L����^�evk�Q/^�i��a揕�5�oR�qfG��?S\uq��E��} �߅<����QaK�ڭ}eWJd���eX�W�7<5�b�������V/A����V�Z��w�n��E���T&C�Q�ک?{�v�|��A�q?`�Q�҂ �ܿO����ԺM�K�>��3L�67U-���@+��iJ�~��%�C����GBcq� �,̵s�����ψ�v�F��81K!��qom��f�멁���ՕPe��N7}|�0~"�A�1�~L��C�:���'7ƫ�a�zo"Q7�Jɶ�(%c�����i���'�I̔�t��&v���?A;/!D��&�H嫣Ddu(׋nj��VI��#,(�^V�=r��Ԁs��������\�G�ٸ�ZW�֦z'&���;�5�`8���.���j~�x4 
�����NE��H����ޤ~�Z	�/�"$�>���7T�m�t��N�%��r��G���<��iA�"nde~�N�C2���<��C�+�X��2�4��C�h&tQ)��h��"^�� <c�;9,b�|P0	��a�1���@d2�GN��J�X[Z�EȰf2L e�P@C���4m���g�Cz5�D�ܵ\�r
���^���B��q�"[���������zu�O�BY����Q?M��u�Zhv�a���/e�j�/�	�����ɲ�B���R ��O\�C�i�t�8�R{��FMwy��V�%�T�����Q-�͞�)���O�H�S3d;�|Y�mA.�3e��-��n����믄WZ�Ny�������w(]m��a��x��j�"$m�&�H�]������ɦ""i�j��UK�g��.�3`�T頃��4閡<rOF;� b�s�����|e�)��b5@Z�c&2� <)�akS�1�д��a��&l��	"��w��`�$���o�<x���Þͅ[��	�Li�d�AT)6A��3��}ܽ'�C��i>�}�epì�@v���,�x�Rs��WI�ܻ�<5):�D*��G��nE�L	ʍ�����S��:&�Ҙ�Tn���0�/zݝF�c>����_������Ӱ����!��i �kL7``�W=�Y����ƣC�"*%��5Pѣ#E�S��ղԈ�qU4����A��}�j��l�!��ɚ ~��d�����B�9����ctU�޳z{�"���6��T҈�1�&�q5E�Gd�7��{u�@��2���[��6�+;}�6��+<�d�����ݷ��š��b�ֻ)�\?�K��z�����w灡��\�)j���tiS���
R�l���S�����7����1�iq�hi`�s\�Ҡ�����n�[C
�oT�n�2G#�֘U�,E��ޜ1B��N��+�Ս{T�L�0P!�R�5���4����=@+~�&3�Bf��+v��eK��"�����rA56�O�Al��Z4'F�B�#@�;[� =�51�֦�p�JV��,�/\��n	���ͥ�J��k��Ȋ-W���#o�`ٖ S3K�0�/��Tc��)�E�>��a��GT���2-��a�"�ƋP#����&S]c�$'��{hS)LZXjL-xXB�a�D*%@V��(s
;�S�$7���a�6���O�w����T{0��oO2�Ow��P2���u!�)NP�d�4O:�C�M��j�b���RC�b'dӹ|����0u�������b�>)ظ�q�_����य�Z�s�M��(�w�|���w��n 2@��#ȆY���V�02qI(L]^�U#�k�c4Sd��.�E�f��h?>��;�uD'di��w@�/��̿Ƥ�V�侜�;�t���|�m��doZ�1��f*|���@)�g�k/��ha�=i���j� ����-_��
�ľH��lj��I��@W¢LkK�@W������2��L9�]��8T�?GQ�L�3Pg����d�'�&"�ب����QˈV-Q ^�w��>���tmv�g�d�bΘ�an�mHs�aÌ��(��,�R�x���-U�us���� ��y?��h=0��0�ּ�j�ԩy�b��j��i��EȔ��Wzf��3�K������I��������/Y��^��bq5;]�m���UB���Ӫ��U!C�W@���H��^�Ct���`T/��H�N�U1�U�����*w	���F����SMQp��A�Ȝx�J8���.\j(��?�_���5�T�@�~�j�;�$��]eMכ��"������qT^�׉ӧ�U1(�g�5�e<'q�b�I#�']f��-g�K/=��@x�F"�:f0r�uC�܋woH�87���o��y�K��nr7������ɍ^q �Dw���d3�x�JB��1&�#�����>�d0�iv�v<*Id���
)|���;�y5�&�� $oyAzi��B	�$\$�*��Q�����d���<���|���ʼ-�o�F>%���_z|�Z��9�����)֭� l�������Mj�:�h����X9%8LXj{)����<2��<��<�ȓ��u�o�ϐ�D��ߞS����!��)��^D��P�7���''��zl�,Ra�!-��n�gN�(l�M�����jOb��#��&��ha��wZX-���0�P�f��\�>�*�: �k7�_���S�dqد0��|g�<��(��,�'��%�tG���5�:�G`�3D�9V�/�m�À���WU[U�#�Өec�H���������3���Ҟ���^�/�j�Mrk.~n��>5���%���ri���D���ʗ}1M�
q�OM��d �1�m��ӏ��$d�߸��/�*b�T����|�xN�~�l͚#��p��ry��r23@��߻����WB�x� �ipxE���ɫ������&:������&
ͦC����f��P�˚�5<pE}��G eqK�ۆl�2Q��d���#:'�⏓�Y98S�0}b1��c�ʶt�@����x�T��XS��<���4�l0��+�&��5Nr�2 �Y��a<�F����d:�\3��,zXn�F�C,2v�0���%��&��6���9ș�9�^x��X4�s��Oe�
n��<��/����Z	�Z�����lv�f�3�9_� ���e�H�7	��u������������Ƥ�K�G�W&)��x9�����ŭ�|X�X�S4>eaT�K������i�so�2H���y�_�*�y�R=���t�7�)c��: �iu�h��_q#��K-Q���lr,��]�[�S[�����XR=B�Cy1��5S���y��k!��й��V���/=���a����؛@��\��G����4es��2"@G��Мh�t"N���qW��˥��^��$?B�s�/�J�m�����n��´;�]i��j5�H9[�h-�톣8���a��b�}�W?�B/�*u� ���r�k���V����)�r0y!��F�򅴸�����B��G�~!բ(�F�P���>**��x�D��,W�.S1,�����gD�y�ZJ�����M4f#������*ߋ�*0����z}�c��J��4�����d��PnX��m��G���2����F�T�3��/��)���!w�!b�ܟ��>M�זe�eP�XV��ZR������s;p>�u���Ng,��%���"��'�|�����r�g�m�\CO~����|��Enk +�BˤsJ{[�RS�z��\�#�5�Y�R\���	����-���Qj%���(iApe����f5�0 �yU��3t,o�y;mٰǇ��d�����9��{ψh�᝚o�k���;:��G;p�KV��;��gZ�Y��J����/U��c�Hɭ\�Aȓ&��e0���� �EZ�z�L��!�K�i�R�#�_s��v�����D��~�>]��b��a&���v�W+���!@���@��Q(!�u��t(�{�Xĸ��1�������3 t8����f�����V�|�U��pO2��N�����FQ����{@ڔ�����ϰy���$�}@��DI�=��} ?v*��j��q����F�z���l/+�w��k�?�Z�ph^N��?���\��ŕ�Ak�y #�M@�4�{��u6L�Ȇ��I"z�1#:<���/���:BcM��4�Щs�	�}j��H��^�0Ŗ�:ݙO�6H�ǹOh�B��?�N�jw)�rR��V&D��ts&�q,�r��pR�?X�O�x�q<>�� UcuY�D�5�-*��v	Ź���x�1�W��Y����Q� Me��sG����)q�-wi��E���ߗ��3|��U�)N�N��������R�q�bp�>^��:��@�i��Sy/�B���e��[d_Y�t�h��`<���/�@>� &����Ѝ�_��id�:�y���x�4�G��縫���V����o�m�$�R������H��bʖ:�l�����T~���Ү聩[�=B��6XU\�)�R7�>��S$'!Y����ɪ�a�B헖[��́��I4���RX����\x�����{xE=d� 'E�(C6�����p ���Xn��"��T�'x�~�#|`��"\�wd�޿��4���s`q����bNx���G��vW�Q�.I`��m����EsT��6qG�h*���5�����F�܊���vS�?�$c�0�&.n����xiB'��|�f�����o/L�;q�s�R��w1>����)�	�'��b�TpwȨ"`Rww�_r���}�D���PJ�m'�G00��-@�X�t2g�챭S�5��b3\��C�	��oe!��,N9L���u�!�ԅ�����Z�ĥ���M.4-�~�%��<���0 D�IʺK/U�o�K:�^�o���N��[�*�(�'�?%����Ѯ�Ȁ@��8��Pʃn�O*ܽ唝\-^����p��j���b�)���?�5Q��WP��&���  ��}Α�C��~�ƕq��6�`��]�*B���s�=���?%OLt������4�4MC[0����2�Cˆ캸�\�Ɣ5�U� ��a�n�13x��]Y��Y[d�ʗ[r���\��	^I����ÿ�R=Y��Lhe�}t����D��Z�Q�Q���Ҟ!Nd�f��GD��;���>�`�mW[P�b~�%+�.wo2l���R�h�υ���6+���&��E�c?�/��{�S��ҩN9�/�5J��7}f�+�@è#��U�S޼V�Nc�23����L3C���J��n;�tYk���oEd��Wi���p����	������<�sUxro�O��b�8O'$cׅ��<*vB���0�roCC�sl@�S:X�'���+1�^9N����g�%�4H/H��.�_ڲ w���\^˕Z�H=��[ث.7.���),Ǟs��#�br�!�����,���. e�w⸌m��xLnV��x���L[?���ԍ��� ���g0�	���@5�*��w��� _��n692�zlIr��c�S�P���d�O��_���oI�.�����Z�y(�X�q5�z�ԴQ}���(O�kB@����	��u���n&�8���m�Ö�	U�S�w�05J�@�k�t3�Ԗ'�N�V����n�Ӎ���_�|��c7ܬh!�K?:a�~Ìb.��<)eϪ`ds�y ������z�;�|m�WZ[e<�)�^ٹ�]�se�A�2UeSfq��3�a�Ba�+@#|�G�U~���~m��2�<ļa 0��'U[k��jF.%�а��6$�g3ۺ���h�ĄX:B�	���z �@]5�QX+�J�mS�F�o;�N�����b�YN~��1�X(��t�u ���j3��A�a�[��:��'�el��Gse��,O�n���/�?�/���E�Lg��3��A,0( ����XC�?難�Q�ђm��<'��l�v\�h���\��6�?؎��	��V��sqV}3��?:�<��|IfԼ%��mܺ��;��?,�U1I� �W�E#3��5�t��Mt �'	L8��~�3v3��7�\�W$+>Ұe�o5~�\j?���,��h����+�H�V6�b3��T�3�ig3��v���_6ԓPTtk��ݸ!�_X�ʄV?����(�se������QQ�,MM�4We{�2qrG`���Fc��Tt؇WJ��0f2���;d�/�9�5X:� �T�m���-a�|��������?;s}�V�W��LY��gưnD���5��W������J�Pj�s�1�9t��b�= #V�%��ܜ��bY���i�?��gP��k���(p�Lȡ��:pE���ʞ���j���q��\8��Gu~�7)��X�XE2�s��Gۜ*���s��3�N��^��D��������94i;DZ�v����Qw����Z������Kf^���Ֆ�Di"+��ە��
��������6��B���t�����mЋ�Z��m|���n@�:0�B@L�[�F?�Q1�͢@�?�y�f��<��Uʁ �BI��b�����y�Y�ii�m��PA}�:·u^x��1���d�&c�d��4���̄�'�H,�2,���eD,,;����t�b+��0�X��%_>z������� yXh�t
X���ו%3�1�$��ܽKvڶ^�x���l�v*_�lI0r�n{��>6�Աs�}WɃ).�y�t����
ߣV
��t}S?ߡGS�-ny�e����͍��j�EP�<��U�"���*㥅�7fZ�ކ�H�u�Lq^��0!7o�ow��m��oono���	�
6��]3kD $�a,	^pE�J�qi(1�Q�0-,u�uq@h|�k4T ���+��e��u�d�3�:���-�p��ba(��BtpA�@�c�a�L/�Ӑ��,l��Y��ɡv ���T�@�0���BL_'�Ʌ+�p�S�J�(9Gghe*���ij�u�L��v��`=4��i��&��R�7�>�Z�z2JTxh���g���?^Լ�\���(�"Ok�j^U�صZ��o�WI8.=֊.I�W'�U$�'R��c��@`�
X����ħ�K���,�kL���Ϩ$�|E�ǆQtE��#i,�a�K~�R�9�Z[���'�q�-پ���d���
�}|+�0��\9�|jI��"��rbR]�괅���5�)]ځ�7Y�#���kJ���ݜ�_��)�	�
 �uYRK!��-�A�����>C?2���%�J���4XV�$�+B�;�,f��2�P���~�I�6T,�K�jv��F���x�j��G���6ӿg�[����ܽo�}���%�ZG�M�E��RF�uj�OJ&U4^QH�5�^o�ɋ55���a��f��|����=N^�I��8���Y�QpF�o)��[�q|�CI+���Itz�I�<"��U����s0�g�8����%��[̩ۉH��������^����蕈�E6�F7A�k�;[ۑv/���&�_���q���F؁68���Yl���6���8٘���i�M}�#��m�u���P��)ʓ��cɣ/(��ޝi�{����]6f=N�c%4���,a�'g0�uMM�P�_���}-�`d�6N�-�lv�@j\Ĕ:r"dI��������E=�8�����CY�$v���_u�a[�Z�01~,���F��I�>�ǎec
"�ƄB$ܳf%�N���g���yG��_����}:��]�& ~�O�GR�[��V�D-+)$.me�3��U������%��M4À���ZM�Ou�)ML(�;�j�x-�`,h���L3�9n�Y�Yz� n���������8���8�i �ԁ*�tJ��P�f�bi��;��C0I�@���*gB1�n�q�ԣ�wb��!D,��(K,���;�"A�@2��MH:��Y��RNipd�R+�}Ct/���HA�PAv����I�$�N�t�xȒKڿ��+��~L���d�5��-�x��xAW�cx�K(���=�)����e��&ʱ�@�\��9����%��EF�Q)�A�O���4��LB�l\�ZD���p�W�$քV�L��������zo89��;��`#���XZ��ߊ� �1U��@�Y5:�f4�'J�g
Gz��o`�Z�0v�k��R>'�|�X�
^����q| �Ga	1G����(���q��n�i@�$5����+4�pz�b���fcjc���p�CW�>�='͓_OEy��`U��
�E���JU4Si��j{+[�}9:mɃ3r���Ȱ�������#�m���k�V!4y��n�ɓn٨rS�ۘf7��`��t%���!J+��$�������i��w����r�TZ���AB�	[��'q�'�}�;m�__�/b�|]aO��!Z��cV�O?s��b��=ׁ�ȌMȩ>���3���0єdG�f��?�'�"�pǻl��F�>K�v���m�S�Ma�тPQts:���h!��a��o#��=��˄�/K}�b�&�W ;�b��o�%i4���%'1X�5/�>\I�X:�u`oҋ�lVeu��8T��7�Ƌ��Z(�P'R�%%�Ax՚��K��� �yȁ-�(���;,��A���'ǟ���?��TP��z���e�LF@����~;=E!7�)��H��o�_�d���w�I�+��]Rc0:�};מ{Pg�rpoō���m7�C������M�v5)��'F��TEڱg�G��G��ͪ�V��tH�f�� I��U�M2S�]��I�雭>�=�w����sߍ��@��P݇@t���	�S�uS�� �m���)nX�)�9q�5�M���p�B&PK��Oo��v�P���V��6�bQ���,�Ĺ�+�u7^�2 �3���_8]��"�܁��~�p�ݍ��5��fe�����,;��J��e��s�ARw��4�&����wd�Ą`�w�]�I@�ou�������qn�zu�K�*�F��iu��2�:S-*),�_$��$ʹ-�FNdSS�^a�;���[��c�	oQR/)��(g%��[wRO��1XAM\���熈��`Һ$T��(�@�.�_�y��ܚ]��1<1���3IS����:�\�u�Y�}.���V��|�4X(�K�a����%Mo�ɜ����\AL��e��z����6�(u�x���^��[�*)d��Q#rdEB���D��>0Uf�d����؍3ɾ+'��;�ʴ��v��<�@����š
>0�Y�!���B�0?�G�9_^0��Sh��+��ʍ�Ni�1�=���{B���`� ��$��mJ�n��@��8�9oq�O^�rɹ}ֈ��2M'	��)L ՘T.������gx����R�/9�4Kz��!lfiğ@9�{�P���z��KK`�H�FzRL�K��b����ݞ���7��)��ѢIIxѵ�<�R��]����EN���'(�������р&�%��4<'�~�sW?k�y9c�O�a=7x��B�#�
c=���=��fO'�����m�������9D��ӈ���gDޟ�+#��p�:���B�J%4�����'�a�u�׼ͺi뀓I��0�ߑY�Q�2�_���s��'�L���2� %۳9e���ڝ9���:j����dK�;�N�k�<#�d;$s�P8B����*�(o$�I�+.pZ7���9��s�ۦP0J��D���ԏ�ds�},!�;�������J�w��`�ڹFӃ��F�1l$��5:�����su�f��C2�;�$�B���[.�pZ;�>5Q��/�G��&��*U�.(�~c���|W�P�"-�fFp����MLЌΣ`3Kx��R�kh�7"�T�l�r���eҔ�飛|'P#�ͻ�љ�4J�8�ev&���_�=Kj#SόQi|>�͠����U�:�k\N�Z�:
6+}@�5eT�����K�mFXb����^�&r^���ǡw��d0!����\8�o�+�~c�Ǉ�o�g�q`�򹃄��˫k���	p���|�/|B��c̤F�-H���u�����"��Lm����3�%�I���;Mf�Z`��l��u�~�*;���
�-��d�x��öj{D��C�+#j��%�^2�^o�(jSY�J<�p�'6�v�&�UXr5Z�d�;Ib%zYZ�x̓'%��&.7l��8o��M�E�⒄���R2Rq�O �$o�Ӏ����b�JJ���a�%��|��ը�, �(�B�����ܤ	�tq�������n)��엱*�:�"���W�$(z��񌾠�R�K���է�*�_b��o�Š�5~$���v-i�L�*��o�%t��ծ/)MD"3G��蠁�6t�F�wl1u���
Ix�*x��='��Ǳn�e�е��<Ј	�������yB��Q|.$]�5^@L�"�y^7�0�c����F �Թ:�lE[��R�;Rj'���q��c%#�I��Ȥ��̰���#���@�c_nc�}ú����nJZ�K�זg��Y� �;��t�*��eWP����Or�W��J��&���p����aZ?�����^6�9=�)$���d'z�*W���a1�)������h�Q�M�-U�/O	�y �u�mm5�z��a��oQ��9i��;��R&������D]����ʝ �v���1�C(5�e��X��0��	�B��q�:j@��Wly��V�	���n���m���jm�o��)�M_�I�}GY� ϳ�O�����软�Z+�W�FyX�/۪_��l�U� ���~�+��V�%߈���ބ���'zO��O��n�5��D��� ��D@�i��燎ke9�B1�w����j����^�*%NHvhI���bݔTI(��^�|9S�#�8M{gDz0>
 =� �3(�@�<XڤRM��AE�^��`f��8�_�ַ�1"�ݾ4Ϗ��ϲW�>s�[����p��x�}���@���O{�V=A���@�$�$5��4�L�p���?�#��MW�`T7O�V˫��V:�	J�o�����jZ׿�u�y�`rV�� *�߅Re�cF+qذ��� ���GE	Gr�1���rT�2��w�Љb[�LY�lO��%-:ơ������b������h;���\2�+���u)GM�M��Gx�#����l��t��B8�](9�C�G����QQL]�����w?޽�uɂ��쬁�t�)���Ȉ�x^E��3Y���lp3�k�7�~��y���.	�Y�&|o�"��f��Z�%Y~��!4�i�1�3��p�ii9E�Q�	��o~E�_� ��X��kͽT;�K����T[��Dq�Պ�3Z\�$ 4b�6gl4����AK|S,pU�<i%6@��~r5��Yc��k����{>�����eFf�~�Y~Vf� "�
�^���}=k�(e�V�$@�x剁,fQ��&�[{Ee�!�dG���{�훵}U.%��\@��5jW$�sN�"k�|���� #?�}�>��U���?��Ho󖬍�[a�h�Le��W��؊�N)�t���]؛>��8y~)ޞ��Fצ8�0��|Aφ�l7�Xg�u,�8��}�b�_�ߕ G�t6=�v!ԃg���Ҧ�iJ��j�P!kp����&�ͅT�\zX����TY����]���s��	.W6�'�yq�X�"|��^mk�?�r�f�r[��ǿ
��|��2s��Jlev�8��sU�����rR�N�N�z���W&(�q���t��ڐ��x<Ysd�);������v��� ĥ&���On_��ԕ%�i�YlC����4s;%i����o�d�v�Ż�b(9��Rn���[�hvT��T���)��'Q�ە>Ầ΁��{���o����&G 0u��C0f�L�ڦ�TZ^���=��� -B�^fe��*9��0e���?21��l��ք���rp�&�E���vŰ� vߧ^���<|�,�u����F�w����]3����]�"P�#�ڬU�F<���4�sI9"�V��R�tt��� ��Ե�g9��E��2_�N���jO=���������I���F-����Yv��Dty?��ɓ4�c^F|��Y 	�-M�N�ͥ�ج~x�<�x��5ê�M�
|�0HXe���>,>����E��k��󵤥�#e���5���o\T�@�_,��V.ܭϨ%���k���$Xz��xmh�?���N��X2&vs{����ib"�nG�X{�Yu�6��3��4�d�%	"-��%��6�/Ŀ���֬���/Z����EmT��5�JUB���Ln�&Wҗ�M8 �H��RC��&��+�R1�}G<u9�ʸn��S�nWΕ�h�|^��?n���ܶ�ӵ�>a��)��\'a;q�!��d��V�A�u�-��cB��Q~���I���%���&ڇ��?���)O�}�J�}�D���+?hn�x�"W�����R��Dss�	���|W��/��ҽu��c�������|�,xO¸i���зԾd��g��*^ K\��y�>rUlS����t���<�����S�{Ũ�4J�ȣ)�]Ԝ�~�����*��{!��W�6�\�Azp��G�I��Ò��ea{�Y�-46s��������1��+��/���Q�N��Ib��돥w>�:�@��%��o�nϴ;o	 ѥ^�I��bU�qy`,;�dv�û�Bu�2v��6��o
g"I\���/�x�M�Wд؉!B�5��K����ĹA��Z����~���)rҢ���˷���|��g�|v7��}/���[��j�����;���h���1�Ϭ�@�Et�ηޡ+��09.����"�k��:�F}���zf�¾#2�tj�i@�/98$��M�'}�_��'C��0|�l��fr͕2���@5�ޕc��Yc��Ƭ9%��05t���+��Z�V�A�	]�ߔ�� �C���7
CD�����-�+�1]���ƾA�3�����I.�Mm������.ߏO�C�I��#�_�ƏDE�nۜM���˫j�;73%�*N?����j���!�ّx��+��>���=��Q���������R�I3�N^x��d�%r��h���,��s9!f1�"���(O�V��G������g��#�LY�׋j<9��KtO$nN;[�S�'$�~g�v�q�B!$ʈ�)t�~#F$�K�L3��n��i���B�ޚ��%���{M+;9��Ƶ�h*"9��	�P>��K�����1�;6�X�IN@{?;��� 8bc��>��15zD� \���M�aj"��H�~�Rǁ�ߏ!:�]�F�U�X�Z6-Z�$eO۫\#�O˝��3������s��E��ebD����K#t�ptiF�O� �W�4n�V�۽���?�ʛ�V�0'q?������t�[H� 4��I��D{]V��,��x�vʺ��H�� |/��t_��}l/p�-�/X�WQ_PN~��-i���6F5���e<��4�J��Y�1k�3���3iƯm��D5���Ԟd��������u����c�ֲ�$Qm�<�ir!SQlɒ��2�A��]RI�d1F�d��l���Kab��(XX6GZ�[Q�[n�Q�膿)�)��qqw#Q�h�v},�/ٚr�Gi�هVZ8OPz�&K�!��g`u%��x������{�0:2c����LL,�#B�H&r��	(�RD�&cEUX�5������m7�t�ZSx G<b��.��Í�*����/�Շ���蠯�����G]�y{n��ٵs۱�MM��e�o.�7�ēw���R6W���0���3��Q��y�2�a@���e&�xd:z�衴B��@:?i1x�D�mː�"��J���/�*��fpH@��D�g��0#I�=yoH���SN��e���e�*K�*.����Y��+�>t��EF� ��ݺ��ܿ���#M�!�#���x�-2N�G��pw��iΉ�B𘙗���V��wztL�QdF�f�P��U_./8t�PG���mIk6��`�T��f#]�h3o�I3#�Ñ�|��e��o��7��D`|u��Biz�N�?֬Wmqǵ�"�>��H�&���in�s�	O��<'��wC�w�"�?���D��g|�g�ط��j�LAwc8�#BY�ó!ٵP)���X�ݛ�	��P4�X|H��;v>��=��j/�Р-s��z$�g�$����:�,�6���8�DcP��N(یC��v���݈n��sҎ���'J� ������*�d"v�k��`��c)�n^�F��ƴ�NRt�+�~��B���o�!��U�]C���sQ=,��m��ܷ����Ԕ;���'c���>ʋ!��<��������� �f@���Ưe����pS�?���s�����*��~�O�Jٷ20�[Y�D�*P��`a	���d�h��z#��[2��%&���#��?�_f�@k K�_�{]o*޹s������E�=�ݍ~�@H'�4-�Rq���.b��F��1a�bS�GX���Ӯ�4) ���k&�/����_H�H]�Rv-��5����:�SN7�������e>c@g�����9�A��0h*���7�R�"��(Kx`-�h�~���I�S��5��v,��ykKjR��P��t]���<�}%�Ȓh��T�L�<�R&j��J�L��s�N�w�U�Ϸ�Sl"�FT�ʕJ�upH\��'��2v�y�y}�3Hv�A>6�d�U@�Ӝ��	f�))������x��9h�g����鏾��#���:�a�l(ԙ��3y
�i���:7�u�=H��u4�Wm��T��OS��އ���H���uzJ��on���P��^��hʸD"r*N#�)�݁�M;�<
��	ڋ����̂�rb;AG�S���傱�������f�0�`�����IA$e��M�S*2"��|#���g[6� �AUS'��,xP��F�Om�	�]���U���a��67�,�0f���D 29���>x����춥k4�P�Wf t�)���c�stܭ�! ��ǒ�����82�a3�'��rUxl�F��*��7��c:b
g��]�\�w���ɨCQz��4h��ij��1��&��g ]��~k����:�d���X3Wb�R�����
L�7����*�q����r���K:1�G���w�l���m���bKf�(ʸ�T�X�=Mc�C9����-���gk�J@��~k�4�ι���&�i���xx&^�Z_���}f�1a���Rl��~�<�����=��<� �ԕ]�:OHh���x�CM���������*���%����=�C]sm0a:�.J�0�lf���;�C�w/n����nl�=g��~/�=�T/�!��W߃)��1/��˝���R�P�=SI�5����Uϒ����(��=���im#��)�DF�O� �'������Fn�ۂ��_�*�2���<����?e_��~� _hN>�~�u�D�~@)�����?�n.�?�/olk΃�Yw��k�7���� R��=�K��jrxŸj8�D�uI�;���w̹މ�ѫ�EV6�B�8>�/��'�!E
b�G�5��'6����:_}rE��]Vd��B'{b�Mܙz�	
�����vŸy75��d��5UO�$�	*�[[Hu6�W�Hȶn5�3d@a>\�`�Q���Q�����߰L��<�7�Qd5D�����KUc/�7Ds����^��������m��b^��0�;��)��F�\3`s��e4��!���#!�mV3�~��M|lx,�����O��z7��&"�b�a ����E��C�t�_�e����C>��5�|��vo���!��c����1�
w�e�J��f�Q�]	�+�ք�M���wwh��1��"W���w��9)� �h�˟���HdO���dV��_�um)V�9D����-�+�On�up����$�"���O/J� ����B�)�шTI��@yC��ZcL۬D�~9,�T���'���F1�����R�E�jR/X�ϖ7�M�0z7�M�L�|��l짪X'1��뛦%�&a��&��8���~RtP���u4R��m��皫�f�ي����Z ���S��?uFa86֛�>�3������=�dTL�kqI���u,��+��P]}/�@y���
$*�xduq#o�Ipx�C�qW�����`q�K�wU2�QՄ&��*�s��Pa!;��F���v�N�	�,�z�>-Fe����n�T��Zm�U3�hP(d�M����/���D�M�����[JūZ��u�m��4������AC͑/�	�ԯ�Y�z�GIR����p��
:�BI\�p	a������s�Qxac)����S��v�J��mԳ�`vL=@�!?P�F1���IR�\0�3o�S��+��9+���Qu��-��u� !	i<Q^+�t玖ыcI����!�����;��P=�i�Sѷ�ͳvֺ1�̃�7_��]J�>w�M]��c	�z�YS��`K�o�#�|�C�,!L���Vrr� u���k�	=J�u/�,��49�"]�	��R ��dW����s�ߏ2�9���cn��b�!�=4��.�,�K��z,�m �K�T�LU6�����j|�ڑ��t���{�����ja��Xyf!+�m�f�Q�y�v�W��gn.���p��+����o[����c{D6Vm��Z�R����N�k	Ëup�囈�i���%*�[����8t������uC�L����%�;Rm��7/��d�X�9L�.F�rM�Y:`{���슥��u=K_��5w!��=�ω�<��O��V�G�]�<6smؔ��癉�� ����6Rx��T6B��p���OȺFl��`���Kma #Έj��	7�r���O ��+m��+i�Ks��Cin���M�ߊ�~ Pd�3�o�fVr���tVe�P�{p�����4o�pҎ�� T>Gے�"�G	�t�߹�B�륐ۡ�]�+;���\��m@�"�<o�dk���Q�uK�Z ~�� PT_N��a��p�-��$�ɶy���	���_H3HH#ƛ����vդ�m� ��^�6W<I���N�D�h��y[c����eݯܕ�6��sN��)Bϑ�<�x�E�T褦���N�*�y@��09ĉ7D�/�mJ1"y�i|�1B�W��B��}Z�����H���1� �����;�\����XnDr��L7�W��*��r��E����������I���bx�!h�@Pl��!����`��7EP��r�,KmzL�+H޴�ȫ3�b�z��_��Jj�Lv���;�c�[�n��<���v�o����'SqT>�D$�'���D����@��B�(�=��\^ŋ_(*'��RIm2����@vEj9���k O�!�"f:���G���$����h]����N;�8�o��.����Fڅ��ʖZ��>8ڞN���?�ld�kkH��`�76�u��x��Nx[y��P`�;ѧ�s���fc�<;�,��[($.�=vʲt15\��,��~ �yHō� ��噪�����Ohڇ3�,�*�0�L36���X>59Z�*]^�G���.�Œ��ނ\�uf��m�s��1]�1��hG���5 ��8�p{��\�Z3]8V��JDh;tpD_y��J4ǣ>�44���V�C��$=[?�'�0;>[�U�v?�2l�p�|���k��	��|�-
�l�{F>��V���.AC�����]�j�3ϑDq�"�u�#��%u"<44�c A��f�j���$�O�u�7��?�+E��^z��{,S�8fr�X����|�P�N�C�����I�=�d��߁l�~���آ��d� &���|p/�[e��lwhS?E��޼z2�����bL� #���R�9zLg�����`�9Z��Ǔ�y��̓9����~{��Rǭ��kL�Q9<��;f���J9��O!mnF�,|�!5v����L:��q��W�ʵ-x�ٌ���G#�a��9u�-y����������&3+!��Ӳ�d�Ő�M�(�O;�&�����1G� ܵO[m�ϭ����o��?ݐl�Y�@�4��%.zPf���6��b��/�� ���²�9����2� �5��b���{�,l	ni�*C�������]ϡjb�k�c�������i2C]�,MCk�$��%ֲ��v	ǋRTY秈;�^A���ëK��Sf�:AH��c�U��D��
�SSQ�/�-F"�inPM+R���#m�T|C��k�?b��:n���`�,����A�⸍o�u�o���w
XRX�p�����vV~�b����i�J;P�Q�����,J!G]?��~Q0<�.���j���v�9���^��̕���I�n1�(�7����M�\|Ct��r�%w�&�:C`$��0IT�'3~y�ۊ�ّ�ֺ�I�)W��B�
uV�J��ƞ�F�h��� ��ae칅��f�Zn���ԙ��%:a�Ӌ�Ԝ>�S�5Ɣa�I���7|��|�+��Q(�`4H/:�L��y�D	u���3�����H k��s�[[=��U*�$���<�O&Ǔp����**x����'�ˬ0B���>&��|�dueLW��jaЅ�l`>b����#7XX� �����Z �4�7Ҫ�����Q>�wڐ���F)��1�u(e�{��?�S���ɐ��ugĜ�N�����e�єlh�-�$��l7���YԳ;vƚ���w!k���؁��.)0�~9(l][ZA/Έ��5�a�.?B�����4혊���K��*�F��F[aZ�V�Wz�����
�W-D2~Y��3}�޴�{�w8��xb=�,ϖ>�&����W؅L��%�E~�S����p�@S��[�`4t1�No�L%^KM��ܺ٥���;��C���.�1�>����a�A�z��:���(��Ά��c���b4�����2��,���˟����.m�4׺�!8�:N�+v�,D�8N]=�EK�q�d��%F�B"������{7������K���~�k�Hsfs������)��ck��ƞ�)��#I�E!up7W�`��|K1@��j�����z]�m1�4�-����BZ1�E�����䓶�����e%�}; �=�,�h��{��#��E��e�.!�(�Z���>�|�I�l�I����ࣟ3bp�gϷ�a1�F��m��Q1|�<%k��C��m}T2jKkh.��>-�'\�DA(g�(��6�3��u��R���p/[m*�"�e[��2��8���ˡ���_#ގ��Q��A�Q��J�=��&�`F/�V�w�<�G���2ٯ2���rj�>�I�g����3k���1��-�u8a���^ZEo¬�;R�e���������=�I�Mp2��*� vH���ҳ+�#�_+���9��<�;�C{ �{:r��mf7!ⷈλ���n�c��T񒒆���}�Q��h��_���g�\�Ϯ��O��
�Ew�f�.�ً:�0��0�"y�n y3��|Ql���Py�V���[�m1��j
�`Q�׃��Ǯ�<��xg�$H�lDq�+��u��D��	.���A�'�o�����{`����HBH���$]eH!+'�7#(��;�����ȨL*o��2(��V��i���D�n	zfNT�;f1?-!,°�
l_ % ۯ$D:��8�:=~���r���t ���qY5�2)	����\G��e�*���
b�>Px�Ĉ��-U��/�Z[ס�\'�I�wZ0�akbx6
KN����|�Q���hi��
�c����(�U�����l�+Lq9y2�����e�5>���J���Z{�'�5�Έ�C�e#^�}��"j�k����Hj%��ˢ�|]I��یjn�;fS���x8O�!��=���ٖ��Q���1=��)r�7����ي� ?���Umh�E�j������+�b^�1(��u���es�v}�	CV�@�Ũ�Kb�����4���BA�V'� 
Cy��8�FRB_�
6����"D�\��m.��/�Vy��x7 �p� ��W3^�fj��� ��G(*�D�Qmqa����Q��軪�t���ixٶ-��38�[�2g���m��:5T\�d�-I²\���s q2����P6��y)Ȳ�F�|Ek=f�=&: T	� i��Ρ@��[3>CHlU����:����/N��e�:(��N� ��D��3�ՍߤF^�*Ɯ8h�?3_��2zɖ��v�V!S6���1��5�E�ə����i��1U0�S��P�y�	�����*��Mf#�=����ef�W�_wD��3H�&+�a.��"t�S	a՞pQ�;n�L�e[4�x�'����_�s�L���$�<�t?��%�x҈���[i����KDxepT*�c��n�آw���-������{�/�]�%�IJ��P�l3��Ųw� ﻷ�P�r�$���z[�Cp�:�w�6D�U��A�p �yӿ�}b1��g�+I*�e�!��f�ؿ��\�@AB���ga�$��_���/":�'���]D6�tR49 }}�N�� ���*ea�'��'*�?�> ��^�@n��Z������7>O�����W�8�k0�#I׋�8�3Dt�����ӻ�IQ�]��+��p��w��ZY�@E	Rb�W�?f�r���s��s3s�W˂z]��a���L�*]�BB���_�\iPQ�Ϟ����� �^ܙ<�ֽ]��������A��N�рo
����ֵ���«���Æ����v
��*@=�a��Y5X���:�le�.�0�U�2k�p#�p�n����H@�
�h�Y&�N��Z��b�`f%d1=���)ÔN��E���"*�R�Mӯ�#��s��*���B*���ɦ�Kn�S�����)M|�����)�&c�Y���1�@H�Cs?�T\�0C�H<-�,_e��2H�H�)k����^��7ΩV���P�4��J �#rj�ny���IbQw���{Gv�q�=�J�z���X<�_�����L����?���ׂOv/8��A��$>�G3�1�T����\Sm�xOf������+#�t�B�H���l*�	L�pi��HI�Q��N�nDG�2�������(���J�|���Y��z�����X[��$�Q&RQO��oC�N���V��|�.�[�v�n���b�Ǧy�^G�����ipz���vY��3̽��ʨ��.K��z�z�x�>�*���o��b��:.L�ë{ � 1.0���[9*y��b������x�
 ���u�W�F��٤q�c��.��ֿ[;��8e 7S��0�7gp�
���O��c�}�t�����J��.�̖ˢO��8�B	�.��z���k��י]�=�a̸�%ޭ$=#Bssr�>��5�2C�uJ*A?<��Z�=���EH����=�+��������R��<�sh���'��j�3��0m����{
���Cm�����t��Irs��Aa�@������!����$v��&l���O[��Шdb(te��׭3�X�u-!G0�m�A(�oΕd
9����W!��f�|��dxY��CI��S�\F���E��[c�%ـ�o�M۰����CYE=��ƴY������,|����n��ݣ�R�C��s�	9ƒx�D	r�x)��*em:�Q'=�)�1�g4?tMjaf�̐����g�c�ڰ@?I�:�GWЦ����$LI��~+xd�_nr�G�8��	E��u�WN�5�g���G{;����Q�����Ir��WN1Q�����v5�{�3b��V��2#&���+y3�Ƒ9��9P�5��{���d"ܙGzVteJp���5��'�(N�&̼{�90H�x�
��m$�Mד����e|ܨ�.��h��Z�b��o��v�N&W��_���D�ge�|ŝrL�>A��5w�oAx��$�|�AL1�٥U�a��t@���IG���]�W�\V�H�osF��n��eB<	���9œ�����4B���A�-�=�j�vWFa�Ğ �q�v�,��Џ�uڐ��?D��#0ɍ�"�:l%�u��bX�(P!�n瞳�`ԻD�� ���H�8�n4ӻ>��֖���A�9b�e�R��]j�Tkk{��)} kp�p���u�5#�\��sH�xS����\\�W^��-����9yH�Ek[vQh��&�K�����["���<�\�������r+E韺���$�NO�g�����'n�a�qt�U�xK"+|���v��A�;���nd��
�*WLi|׎LV���а"��M|AC�J�Q�	���M>w�>M����
+D����^�u��u/ϙ1xO�nֽ��PO�i�[J���Ł}���!�����X&G��KU�i�M����e�F���E׉���7�Ժ�ݫ�=\cS[�JwX94�?�8�̙M|vr�U��㓏��48�Rl�f{as��a=���6!`��,��E�x���k�q����9�_˞_��r�g��h�*?�&���0����Z��m�G�&A����P�'B%����JM{�N�F�.��'A�-��F �{�@�gr�n���,�A�鹟���8Ѿ�4�[���񍜫�4�X��w�z�)E�4�1@�>^ͧ
+ݹ�_E��a�u��߿��+��c�f�WK�#�"�{h!�~�RK�8o�+�^Z��ϣ^�s��x#�=��}�M����x7�1E!��8�I[l`͎z@ҿ{_HjOPq��
���R�5�n&3�<l�p�v&���U������J�jtG@��9��_��U�mGr���Ύo*d[�Q�E��|�OK<��昣6���&Aڰbh�K���#羜ީī�4x��~���ٗ;��Ǐ�5�ZS/�[��]f�D���tr��ۏ��{S�l��S���Z���vkg#�OP�Sm��%�
�0�'J��=���-%�*J�˽��|��/�M��=B�(1��O���0�ae�*' �)�iHS�%ׄ"j� +?~b ���vز&v��f�O�����W�D��R���z�ƻ4@ ���t��`@q+Ee�gӔ l�d��sJ�1�ӵ��i�ߟk��+�B&���}��c�Z�Mp]^�o'>��,�d�<�^���)�r%pq��|�5�h9޾��'�̂�}�Tr������(�@)!�mP@��l����J�O���V�q�O�8��l	���z��	2�_�w'��^�����?:�T�<mzY�l�%���ⷳ}�ƻ��O��7H���M�Ə��4B����:ḰFS��� ����k��mj�fV{���efP�pDF�1�;S���֐k��Ċ�_��Q�Ȏ�6��=���rIY:���r0�udm�������LU�7�B�Z�)Cǌ�-�\���ć����-��{�LA8�m�/B�A�t�	x�Q�&�w����:���э���������c<�+	kȵJ�Mn�����)�P�ˀ �9����H[��}�\�Ce���I�qW�t;v�5���R�LY�*��7%A�cm�ZX lj\wJi0i'͗�5M҄��=f�]>Q
;��]D�l��E�gA��AM�<:%#]��3/�_e����.����^��?}�f���R-
ߴ`
�����F��h�+݄-�P����;�ˣ�R���B5�K@F#[S��'��Y-��pl���P�Hf�9����E�ì/z�I@����%��H㱸�F&
��*��N�>����v�KA��k���{)��� d���A���j9u����ч���V�|�M$����3{2�Xye��.� =1��2�js�?$���IG�U:�覴3���<kwٲ�"��\�����^&�+Sa3gמ�0��f���0����D���)����Q�;p?J���<t<�@��/v���8;4A�x�y��!����$؞x4�<�����N��*]�2�4\�����@h(�?�h�2?B",��u�����Zd�+���d���;�K	�5R�ד��+a��dwP*\	�l���mEر�s�>���t�����|�3p��L��0e��:��ג��Jl����ޟ����g���)-���Ȗ?�:k��/�.�I�UM�3W�����
��f��!�e-7P鋁lW��#\�t�z{ ��H7\����������&�dFva/!-�v����4��ǲ��c��p���ʩ���/�N�rf�H@Mz�bk�J��C[���"}Z-0C0;�12`�^����PH�&�`��,mh_C<CE.x��G
<w�!��*�v~�Ӭ�?����;z�tz^��\�
>a�(�A7dx��wݨP���eX���ˈ��R&˼�1js����]��!�2M �#:���g�8@��-�}��8�~�>�ё���h.r��!";צm'�����qB V'���K7���\;�'�g�M�����ԡ�d��%�4IKy$>�=�Y����>z����d�C+y �8�v�n�C����REU"���&��2��'��/����%����{F�/_ۄ�=z���0�z�	M�s��D���K�Z�99�ͩL!�l�m�ڲj��TT�w}s%� �s��觉G��8[ O^�Mw�J!�^�l�PF"�홄�ɽ9��%�)i��Vج�=�@`D�������uYw����� _�!g+��q��� �R�6�X��d�w�MD�%��V������ej	�����S�?���O�e� 9��
�N�N=��ز��}|;�T�6R��)R�-=�g�
��.#7�(a�xo�-�8+���b1n|��@UN�J;�WU�V7	�~��OoF��_�e*l!�7�7�s�q�m�PЃX�(��W����-�7Z�2���iF�y�ۚ"\��Z�K�� ��۝\tQ����'�P̼I��p��� J:p$�o��`�󁸻������_�(zl��O0 ���EJ�>�P	F)�E��2��_�\��3�E��No��v^:��30�{{����j���Z^y�l�<�(]���&O]�b���D��J��ӣ��Z��Q��u��gQ�H{R��z��lt��:Z�����hV�&���@��˔.��c7)B��
��d��=ܻ��iK���q��9v	��,Q��O�\���?C�C�o���g�����;4s{��)*�~���Ab�.����=$�kx�^���2� ()��kƣf�ko���f�����'65�p�F�����Y��Es5ϬQW�� ���
v�9�<��t-Q�-"2%�A��{��xh�!s�p��}Ki����FsO��z3/*��,ˑ� �B�v�I�C��:e�����y�Z�*�j��s����G�b�e�(u��t�d��q���^G>�������94~���LT	���슘s�;.�=n��y�~�7��{M��3?�
KcMhL��21,	�Ri�7�:�����k��cs�=\(LڍcD�й)o���v�(��X=�@�V)F�<�Im�ě9k@{~{�B�o�wqC�L,e?��z̈��P������m��B^�����]8`O��2=Q8�Q��p�?��`������ݩ�$�ۄ�Ə�H/��+~�X�}���s*��Z�~7��������Qk�'�7��q�i` u�$V~�Xu����J.,�����r�y�{���<�a���i 0��:�4/^��l}���T)�'_�A��L��r&�Ơ}8p��-��~����u��)�9-HR�X�ߩ�k )���_}�(ޕ!�������ig:�}�;W��T�kqأ؛Rs�qR��Z5�Cd �;N?넚L��n�#J�tg�+
}��i-K�T�hLr����%2����l�`@��� \�㸥�$��c.���lj�ʗsbi��F�Mg�0��hW�J�H��% ���^��+�{�>\�[�_t����ʞ�?��+1���dC�Kd�k0�3�"��i\��[E�u^�0K}�[��Jߗ�w܉����Y�J#��O#ʉ�\aY���{��e�NY��P�J���P�W~�C��z��}�g�7	瓓�.�5_c�^&['�ֽ)Nژ�
z_b)���\-���6E�h�(��(�}�MS��g�2�<=��Jg�@��)��u+����Dr
��Щ4t�1��^a}�9y�O���)�u�����#�"�<C�g��/C�^e��xTb,��>�{FЙ'����H���4�����Z����X\��w�^A������A�* �vo/��@b�E(4$L����Q�:��l��ޏ2y�0po#.��)]T���.ⶶ��(�n���܅���\��KڥO6S���=(�0��/����X�Y�7.�lCU��zeA�� ��������5�`���_�xr��yZ�a��m�bU���WC`F�����xsg��Y�b��k9 �K������Z�m2���[���/�Au�kj��ɑv7��3�������w!%���ћ��&�!�v��� Ow[�/0Ƹ�1�|��y!\��������5+�0���lkkz��|�{�BG�s�Gw��>�l�jgʵ���ߴyLS5���	�'�1�D��a�k�9L���C��U�/�J7AX�b=����M�e�Z�U�}G�'+�qk�թ�E�7yTK6k:�����ɝ�]aN��bgݿ�J��q�P�;��&��
��2��k=5^
4�a�l�n�`*�L��焕�&l
�	a�JدOVV��2�
qQ��=��bv,1' ��j%���_�X�G6�l�e�)�ѫ�ĉ�� J�mdvN��{``R�Z����dw��l�h [�v��z�.���$��G�����&w眞eIE
�RU��|f�	8yݘP2%��r��-��Rđ����v�<|��rD�xo�ѐ����z���`�t�3� ��IL���ꐘ�ŋ�q���-$��(4�P$x�4�wv����Ƙ�\��i&�����?����oU?}�/�����W��)&�4�&����(0�1���c�8�����t{M�ֆ\^���VM/�D͢�����+؎����N<�׮*6�6c�,�����PO����c�-:�kK�#~�v�"{pdW��;8��Wym��2�u-�x��s&��dk;N�of@�U>*_]Ԗ��46�I<9R�aԼ��7�ƬA��\Ts�:��Ǹɩ
	����޽�l
X�4D���]��</iv��hK�IR��&9���N��܁9�_��0��c*l��"9�Y��r��wj�O���Y>�
�e�D��C+|F_&��W{��l��G��ux���L��/8ζu>�0�X����/#�fF��摘9��%"��d�9Q"�ŵ˞����X���`����Z�|73��A�f�	ÿ+��~Z���+�$��ș��M�T0պa�SymjBhȩ��m�������5*��]o��3�����<��œ�zA�5Á�_0$�ҤȢ���?�at�(N�8��ʈ��](�V%?.�@������nce7dˢ'��>ڎ��m����pc�'�U2'��<�5�~�k�z���%����~�^�f�xfh��X@J�̓��,Rs]�B͝��<s�P�<r
���x2��gE��[���o�)��F��W)2��B ����\�#$��A(�^W�sq�]9���p���&p�)�K� ��b�u��v��'�}�]�I�{�󏬣x���a��4?���d|P��ƌp_3\�lF35��6�r�������xv�,��}���Ģj���/���~�@�+y_��7K��W�3k����,91F#�Ȁ��%P5�}6�u}E��_CRԖGjg�(�[[b�b$d�v�y3�89#����r���
��r�n7�և�()���T��X �n<��6��
*�G��W ���`ɾ�Zk�i��0��%�̒=:K_6+x�U��hkN��T6L�2j�m1"�B���=S������T_Mq����Cvj��P=y �ՆL�|�[�FS�X��ø\6����Ws��Y�T�yv]Ԏ�5-S7ct#K�ϵ#�� ��G��sBz���#�	 �p	�����g�NZ�h�����te3ᒛQ^�❧0&�a�ttKQ*8BIY�;���-��T���n���/�W ��'�D�������P����^g$�/��4����=��_����O���y��WM�{�OL�ts��7�×LU���<�#����)������`��/b46# �� �����[O��k���@��L���^��K^�3�@�B��I�{)_�Wa��v�"�D� �g~e�:3Wsw��T����%���>ie<��uw��`]��Ā>5��WDn!zi��D�B�Ҩ�Wsc�1��<��܎���#�I� ��!ش���"�:����9b��ή����2謢D�������뤃\���XD݉-���2x�HcS�+C+Q�Aw	�[�,�+�*�G�$�ML�~R�� =p����!O�C�w��Qm%�#�8��#$��J/�����3��[�tݓ�|�M�vb!�L����D+�`<
���x�3P�O���&�V-�5� !*��)ng�%�eaiG��bDU�I��@kφ�8V`1���f��M
��fV��0\X��]��-���4�,+m_]ꬢf9i�C5T4,�>3+dY%����z��>7澉4�j_�Z�UN�C�붎��r��r�x��D��RVT�4�C�p�OG�}�ڋ�>~�>+��L����|�����-�zr�ྼ��̂�;�<o����Ho�*� �.3�N
ݥ��J�R� �<VW�x�Ȉ���	���*M���S��=bx��GX]��g���~C�/��rvș 6�9�ds���b�8=����G��o��"�W]���v�}��aahq��ʃr%D��8'��QCS/�?'��" ��^#ώ� �Fy��8��{l��l	���u�j\�7���=q{�{@�殞��Y|6��Ez�ʿ-�3�[��Z25�>q�&��| [�nw�2{���]K�)?����$h~�$��n�T�G+	hg���7����؃��7�$�Ͽ;nlcs�[�G��������.q0���1� W*��&Bi�:�t���T�?n�������T/�	��Q(��3^��*�=P��k��`Tsӓ$�.��S�dN[�m@ja^!X����O�>n��>�qS�ܮsm
ֵ���ˠۍ}�� �yPf����iv?���iμ��!At���½t�w���R������B!������,�����H�RBߟͲN
�F�|Z�1�����`4Ɋy�<[#��A��Ϳ�_�+���ea?�kH[�T���?<��N�1�O���;����5�JX��qǨC�%�=���d�'1���$�Z�qep��/�B�����OVEB�-O���7�p4
˶M��{��\0���@�ZIL��Y�|<�P�S3EhR����a����5�B@��;w�zZ!ˆ�M��*�>Dl������T4Q��ˍΐX����E��d�����L%��Hx�Z�ͧ�P�*qN��;z;f���Ř���;Z�68��� �� \3g�C�_����Nf��zf,�3�3�&vi����vL4 cD���k�7��������]'��u{Zg����O�Y+�(�~%�%�.�xY5�C/�M����`��)6_Ń=`�.�#y���oID�?h�2��+�odw}}U_çJ6`$�B	?ɪ}:o��x:+�WY�����)��8��K����)D��bM|�`2f�]��;'U��M��f�<&	m�v	?y�PyP亜��m��D�I\R�?�<ٱ��/	�J36��c^`Kn�e�����)dK_�)�m�NXo���y|�_�p�����h�oT�&�uB�FH���8
b�24�c��^�5o�f�;��ޞ�*�xA�\s�OV�\�#�bt���%𐣭)z�v�n�.�9qm�[ <f�W�n�F�[f��wn���Ϳ�՗�a
�nE?e	#C�(��(-��F_X��zz��:�Y�\(y�͗&��ߡk�N�f��_̎���k���ʶoN�3�<�ߛ�t�]\�fܯc�69��1C��n�V�ױu�T |�v@ �4�J~�l���_�Af��R��N�7܌���J�S1�T�.�����y%������)f�Z�=���5;�j ��C͹)��]er��Dt�l'g��	T�����NO���]�"�Z�{<0���H1���*�$�Pw�ky3�@�D`ם��ҌI�~z~�bI��t��I�3�f�.�w���7 �=q�v>�}TT�c[>�����5����L�~�]��%����é	���h�>r�hd���QQi�ك\�/o�
������F�N���9�U�qϯ�����l���Zr��5�F7������"��AV1Y�sZiJ���"G�V�c<&�9㤝�;��kͧҌ���d��di�f��ћ$���D�.��x�U��k�M.�N�C㿺�����I,��p'y`ҵVa�
�/�T0��c|��xj�|���9L�3�[~^
P�v�u˺�h	��ll+�-��q=t$ܱAS��uX�ΖF�*��kl2"�1R-HKk�� �Y���l9t�ｚ_ڨ�ڪ�5,]Jpv,h�bF�C�NUP�Gx�5L�D��y�S^�w OJ��A@������������Q�[<�
�`�aH�p��b�'XBRR\th�,�Vx���I����������3d�`����'Nw=[мg.���}����� ��v��k���K�`�bbX9���A0[{��ō�ɩɟ��w{�(ӛ|gq��S�Wk0�:��*bMo'P3M�*TZ�E�	7Bs8(�lu�4e�c�ڐ��&�CQ�w���Lӫ� V�`/J�.sy��0�<�.��"��%e>���������
�	�FøO�*��~�O�����Jz{��1���I^�	=WZ�M�	��A{�YWkx+�<��J�N��2�1(&���h4�Ʃ��d�H5-�V����G�[����c���U�]�q�7e#R&ڕ�c0�[�7IpǬ���"�X&��9#1qqw���0����}�-c�ܣ��^۰� ^����*a�9��[�Y#@	}��D)��� U�2�YTٜ�i��[<�$�(^���m����j������+4������Ԑ8^M�<�!tRG�ꙏ�N��,Qu��7M�x�)������
���2]�>F��+��\�{�n;LFz���Ɖx������Ps��d�>���Xɱu����j���W`�.�d����a��#�������Tb��������H7^"�w�OW�g�Jm;x>�V��ܙ���I�.Յ���h�"57_�8cu2.Y��,�q/iB!^���}�C|�}Q1δ�R���ˎ�.]OqI��=*��kcIz ��?+62ٜ�Ph������SAյ��'@Wj#0`@! ~�F�ܙPv.&�p0��D8�(�^�Лn�g�m���
�u����ϐ&�b���=ͤcw�7'iGfģ<���kKF�$���!h��^��/�
#��h���z5�E6��tX��/z[�D�0�'����G���	�6q�t��)1��a�8qF7j����̘��@�NT��.��``/�'0��"���w:����?=�*�f��\�C�Vl�ii��0�L冫uv�Ǎr'lp����44��
[��}�x"�@Qܩ%{��'�f֬����3�9�8�m�;IQQSL�ah��>kO*E�[5g��J7�G�i":j+Y���E1~t��C�G�0u4���6 �Ԣ���`��y�����px ���-)"f�*)N�T5�fq]���,�<�҇�P���W��=Ev <R��縤�"�����"��j����پdA�6�j:w���U���R���22�b��Nč�H�tZ��M�,#��JrI]{z$:n!>
3D�A�媲�'�X�b����چ�.|���obXZ�+��@F�H�?�4�}�G^�7���YVL�H�۔$�Q�+�mz�E{$�)����'�ˎ_p��2���}�Q�'��������$Mv�vA��Nv?�bz8P9'c����,���W)4�'�MHM��@�w�/�8��X��L��5��l�T�nwJ�H�]1L#q�mϝB����5�v6�f#�����q���'u�}J]3AS9�� U����3Np�2oTM�E6xz�Yk㗍w����{�#MP��0����`}�I�ۿȚWX����b���^Ӯ�M���r}��gC��Kuݳ�j�a���+u5��r���� �
�����9xQ1�F`S�Uj#��$馸.�?S"%A�B�7x���(X&�P��V#8�j���p�����Z�Vldజ6e�o�G�U���;�2�#���	����HIg����3mG��Ǧ�p��E��ճ�yB�\;:�rp��֕ob�	���bJ�8��$�!�S9�>i�/W��W�ퟣ4��.���j|8�3]�%� -�6o0Mo'^ؚ���H{�H*����{�OPhԻ������R;?���Fav��J�O�����7ɮ
���ua�2�H���f��A1��̷&w,�qp�%���<�S��nr�4Ǽ��Ox埕�s�s���K��+���Z2����^�RX7��y7dr~�R�'�j *�Xh�n�'�+�ٙK�p��xB�6�,����#��t�q{RL�0I��.�0����<�b���C,�Q!δ������%7��Eq�Vϟf|4�B0h �'�����R�M?3W�[W����ڻP#8,�����+��C�<x�R�DEG;�/E�hs��z�t|�-�S��u��v@I**Ʌzd/�$ՙ���\�s�E˄�)�LĜ"J���ET�$[�&9r���׷�eL��Qy�?�\ԅ
6��< ��0P��\����^���PQ�6���1z��� ] �l�S@��vR�#�rkK	7��Mq��}o� p��p����� Ǜq��`pl��e�^9t5��q�'3���k$�U3R@�[Om,�'FTgH`�3�]�
���߾��JV�@Ah8;IK�f�cs~y��F����ҷb��k8�*�;D���;���� ��=� �`^����d��6�OV��Z��x��^>X�(1��p`l����;���T�! x�����9�,�tBnU1��2�n&��k��Zư�g�ρ���?�5-г�M��㻊���q[w���Z^Y���φЛ!��l�������pߥ7�F�oI��+Ψ$��Da^���Ɵ��bN�'�^4A�=���W߄]�FZ��Tq;g�[�&�?*���EJ�92�ֻ�l���غ�ӄ�9�U�\Fu������1k���3�t|��[�J8x�lM�'YМ�ΟLK���,6)�G�1�(�Ix��f�*���8^�wiq�5h��x�I�*d��*��`�|�+�4CMv���dBU/�bL�>)'��q�H�o[UC��&��e�MEb_ڍ0ߙN^����֫v��>�w�l6
�'Z$TR�T�d��/Z��%����2ͣ�浧ܛ�CG�~|�)�����r2qs����dg�϶�䷂qBG�ǤAL�̿��F���?ʮ�Nf��g��S%��� �2��2+W���8�pQ�9����U}�ys೰���z�ɟ�w�H�Ɲ�6yB���9ɬ�P��'9襾�'#��&�8�tQWyc@`m�NZ�+\T>f�ke�����l���!�cd�A��ߧ*�fk��<�)��;��N��h��WP&i�μu8��� �R$��)$��m�U��#�N���H@;V��{�"�.�f(�zi��)8��w�,�֤�xK/{�Wp�����n��{�:ʟ�i	[E��e��m�c���=ˉ��͖�|}\R���g؇b��+n��׶���Ե�����}�KFԉ����=�b�%ex�ral}gZ���e�<�W�nLV��L�u��:��V�i�����x6�X|�N)�Ƙǲ�g�|9;�94Y.�\��5X�D��U�?�<Y��?�`Xs��������!G�Y�}�D�{�{ى�;ӹ���t��A��M.�V��j��`ti��8"LV�`M��
�@��F����?� �\�'�r���E�@� ������gԶ�?"m�}ƿ���y��p�.�X1��AL`��qܢ* 6/�B�������y�V�y����g��K�C)6����X�fj�z*�)2�V$/y���J&Z���A�)��O��
�K���_�6�e��5�vZV4w��Q/�f�)����>-<�F���Yqe����1U��UO�0x���n�]U ��U��{$2��Or�����Q���c�-�A;/�@?��g���?A2:�78���|�ld��z:f�^�z�Tpӛ��>u=��r�<O�d��jk��X`C�. LI��tD"��6�w�Pi0nu�lL�����H�L�(s�q�A7���bZKٲ<n5�3�|�%a����mi7lS7�|5���q}/�U��{� L~#�Ʊ��8&�p��=�n_�R�o�ο`_[~g�9��������?�u�IH��7���aǏ���^����{�zT��������o%���ʛd��s�hDf�X��d����ȶX�޾� �����Z�	��Y�!�ޡs��e��VVB>!,�{�����.��56/bi���0��l@����*֬�)ƴ� �e>C�@�����Tyx+Ɲ�_�#{~�v�9�������}i?K�t�̅�O}I�~��z̧e\x�NZ-��F4 ���������;
�=V����ƕ��l��~̗��Y�f����0�����T/W�hY$�S�_vԁ$�!����z�r���T�WY%Uv�a<���� Yǌz�*��W�%vLB:�(=����:�U�(3��>�>���n�[�)�L��h�'�hj�K��%��U +�k��`��I��f�}p\&��+�%@Q�FJD2$��(��?��R�]a��	/�	�9��$"O@�-�d�}���o�ѿ|�(z�b^1������G���#��J���)K������W���K�K�Y��y�כ�Kx��&��UM �#��qe_ŭ��_�����l����ze������~��H��>����)���l;*2�祈��M\x�H5�9�J�/����1�����8r���H�֓��(TsO����Ŧ�o�T��x0�D�����(�r�Q�C�	��4�W���FPu�T�I� �p֭�Ā�V,�o�l��+P��|�0��t�0P��Fv/B�;Ԁ('y�j��_��)��^�:]Y���${�|��H��t���l�HZ�|N�}ɯ��h�3����°Ł��59�l��M��f
�,�'_�&��Y���m����+}�|,�t�5�n5�0륐󱁦���3�V���sɡ��I�L�v��>�,��ԑ)�y���uE��[I?���t���pӴ	��8�v�EZ�u����I���-�U�"3d���g^�T���
N��]a@+�EcѺ�N_3�K*�a��q1"%�XF
��&S|�;6��̴BU4a�Ȩ&̢ �~��$�=����3A�$��wG_;���+6��[�ni%�g\=qRUE]=��J�N�*'@����܋��N"^�fi<��ŷu��G��!�k��A�ިg�����"�u89�皘ܱ�����4������F����3�E	�N�O��)b�li�7�x �	Y�-B���Q���l���r�X���W��ү�BI�3f���R9��`�Z*��j�cL��#���h��?SX�i��{��;Z
:­u�n�ۋ���C�X
`�oa��G+V�۩7��gF���K9j2�K���aQ*;�a1�`.�Cgv�8Th�-n�ޮ�;>=��N@�`Җe�����k�~6�	0�N:��/�;D* A� I��el#��c��&KA`��[���D!P�&�M�/"+$=�S�y7N��bu���7��e�KD��� ��F&�4�ΣR���;�Ϭ	"+}\�RkR���Ƅ� C�� ۱��V�jQ:N�֜�Ojx���nҮm�Yfw��doP#/�B��]<�Ԫ�t�~��(gC��{lc�Ŋ��c|񄫉E�W���_�Mk5�,�w'��d�c��t=n����ޫT��*�ltN6&��a$B.=�O 1�pr^�R$��>�ɐ_�V��?P�AV.C�ᖚ=67v�	M��f¦�Dz�_���$n%�����k�AI�.Zе~(:;`=��:��T���W\�j*��A>��-��9q����Cw�DX�#�hf"�[��J�����1&��sem%M�T}	�ܝ�tS�J|��wc^ F:Ö YIU�&'�JoM��LRJXz�5;
������pA�������o?����;ۊ�׻{_Ut���Ӥ�d�L�R����D!*<`�d|\ 7��{�<��r�1\�c��t��O�������y����fo>��!E	>�S�j���-�#8�Nc,=��
k9���Qux��(]��~>I�݊P�ͫ!���o��g��J�.�O1����wA�)܏c�����98vh�]� ��fg���-�w�)��a��N�"�7[����b�jRޚ.��P�Wb]ʴ����f��w)��Y[ja9d�
�/��^�e<�`���dD5� ����w���)*L���H-�W�1l��kpZ�ypB�Ϻ�WӻQUy��_��D��j�I�30�C��8�,	��K�<e ytO�(�0��B�G0t_�I�������i�K]q�@y:��Fl���Z�Qm�Z�$X���� ��3A�b-#��S�M�_�[�֬�|f�9��o��ʖV��-|�Ve=56��Ɋ��drî{���?������A�x�<�t<�:��vxQ��TЎ����M�c@��f�c�\�85�m��v������D����4F[S�����̃X�
�f�6g�7g�P)�5��b�L{bǜ��&��&d(>����=X0��
P���Q���c=�B�d�&L�n���n�����x�gћ���{#O���ܻ��5.��e��}DX!�I�����4(a`�+�� �
���[A��R��BQd����&}�i��v�m�~-E#W��z2��:�~u�ȏ�\(�
�$c�6Ǯ�0{���b�
ZF�����(u��_��u����;^ʖ��}�9]�n����a_Y嫑����IN쾊|�R���Qn6��2\C��W�xƳ�"�mW�x��mdP��+G�%�07�4��� Gg�1lo����m~��cF�,0'�����i�@p��G�J�ǁ{|
co�5�t�ab���:�Jq�~�t�����e�.՛x�
m9���b��sc�z��7_{�a^�YN�� n5(� �6ٻr���"o�hgF�
�?)�%ɔ��[T�'�G��7����P.o�y�C�Dэn�ψB����k̀R^�j�KY��)�
۷�n;(��'�R3�������-�.��0��s��3|�f��Q}�~�*�ݪ��B�x�"5�xD��!	�����]�#�g��������(��JΓ���D�M��.��υ��9��r��N�F>�:]D%����"�x��M��P��?�/��@���}�^�"�;��A�ѣ���x��Z���#
z�8�
�VĢ4.u�I"��H5d�"��{2�'|�R��a%�aB޲g�s���9�:ӄ�}�ve�A"O5h�),9�r�t�/��X��:W�F�����hC)x6���k&�m��`_�T�N�lUg�:C�"�� m1�	w!N����h�S��w@���Д�H��� �d[d����]DU�IS��
���{�J���.�-A[&��IƗHb�Ӎ��_ZL��ֻ�4�5hG2��N��a�e	ihe������rPm�4��q��J��	y��q&-�h�X�ǩ���Ӊ�|�
�U|(bb����#$Gh���N���-닞q�ܔA�O&K�xʴ��YU��g��t+J����8�C�O��+���WQ�,��	�N���	���y��`���ؼ"u��[i���2xJ1���ֶhQv�Q=�Eb	��@�"�z�Q�;`\@,UόJ�fü��c��������4J���RPD�������%�vZ���E$�̍�1�d���?�L=:�;���̛9
� D��aq�M�9�\Ɔ�HEs��~=�f#�r�b��N,�.��P1�Q,��Sd2p,l*���/_o$����|����IT�	$�:�2�FQ}!p'W���� �
Ϛ���*'�փ݌ �G]D�U�4m�2���,p��3��)$���3O�ye�ȂV;�4�]R�2h<k�K��f�sU�|*	�P��	� �#ӕXܨ\�4��1�� ~@nO��l_#�)>oD;���	�r~��y��OKj��!����yr�'`�QC閳7xCV�����������[;�?�[%��T�Uy�3��k)��)&_}��/��,ҩ@DU�:o- �.*�%�γ���Ja�(�&oJuE�?�cҭ��)��7{�f0�{��FrC��� ��<8�{�M|����d�7wx�$U��#���`�z:�]T���C��������D&���+����P�>�`t;�mhrFX�9nᴴC�V-���׉F�@etOӢ�s��0=��?�`�r=�ű>�6��B�}�p�uirѻ����q��~��{�c��u2���RN�)3ۗ�� ��䜀��Vx�{�R߰3<�����<��q/��F�a�����xT�������$����!SR������L��b�W0z%��6
��	]V(��]�o���A9�$��À�����9(�n��qW�r�%�n-��R��hͺ9�D��I�6&,����!��mr	9�?5���g�Gk�j�j��<I�G��J֛�!l��A������bw|/��n�m̈�6�l�}��~X:
�_��ia��@�v=��?�Ь�j���2��f�/���֒���.�X�-D������<hla���x-;��Df��;#ʥy���6�>!7�+A8����]�U�+�}�4n���1���6�~ip~��k3�D�D5�9w-d?3O���k�D�F-���rx�%=^-�l_��3�CCR�Z�r4.@aEo�2�_	[[���E+���D� ;D�9�����Y0k|'�|�4�����c"Wk�!@���o�_o�T3�b��9�Clq��_>6{�d����$��m��|<��/?\V̨CL���x�
 ����I�j��em����M�}n"+�]%��+	�d�@�orj�����Ĳ����o`����s�E���p��"�0\�x�;�X�z�q�t���Po�q߬���Tj����_��3��|a�Xp�R��2��*1&���l����a�6�?��j�����_\��f�A@�4E�!��I�2�8�Q�m��e�	[�㠻e<yj�at���?�׮+�Ac�^��cSn�(,����_u�����2�(�va�ˡ�J���\zASdH++Ij���M�x-)�zǒYP�QR���|;����G�GvQ��3_H�g�M^���D�̉���áT.���j��e����	z��J�_���͘���g�!��<�FɊ>	k���C�??l�m�`���*�����T�;'<���KO߯;��7�3~�o���G��� ��֞�*�T��H5�Gf
�\O���C*�/��Z%Ě5�o�
�$�uw�� �]jD&)ڄ1�$��<�����.r5ʑ��x�Ԕ,T������q��oK .[&��ǭ#�<*��)�f$"F�˒�ئ��0>I�d��/s��W�\����^)y��rx��K��D�]ڿBN�D���ϸ��&�_�TD��(=O��i�
��@�D�m"� �Ap���Dv���[�+`R�0��p��e�W���hwA)��K�0�*c�7�{xR�/o�f!�*�+c�Q��h���*D�*�M2y;
�aʏ]��(6dC�?gTQD�d�*�hd?.�V� �౿\��*���X�u��]��Sf.����47)(�2g�g��x❏��j�4�x�3?�ut�����.�&�����|�r������~������q�<��
���L�N�Zxp�ya��7J����I���(�N�Ki"��� R !�S�CQ�O6~]L)y괲7/�J���㉕U7�^3+Pųn
�uF���|�z�~'���ˇ�=J�J臂�pKjL�:��|��,r�F@�t]�X�3��s�,�E���2��s�6�/�l�+>K�����W�P�:��9��?y@����U֓X'O�`��	*�P���yU5'�B���
�l���3�n���~��.�7�xЁ�[T����s��N�W�3RT-����ͫq|l?8��P� ������h����:\ܯ&�r�c.�yE �þU_+�*���#GR�C����J�&z��`AIß���w����q|~q�A<��0���I�W��@M�P�X���7VX���u��\���*\�)�v�{!�'��pg
1(����Ei��u+q�j�^Zk��~�Mu?)Â-�B/����H�-�vv��%J8V��(��k/L@���-�����*Xބ%+�D�J�H�GM<�An�����r�����[.���	�E�P�%rl��r�F�
�!�����p F�s�O�ߧ�5F\ҭ���bcu��̭��3�#ۢ��3��}��&�ך�9�t�w��5"�7^ZL�C�	��Ւx��ya��P�wY�7�C�T4��$�J~R 脬�+/��(�F�ֶ�>�����B�*����t	y~l��vd���X��' 7�%+���]�e�Tb��맡	SX(�B���2Q;}wڇOs����������A�|7p��I�rm���xT�l��
�ߟ
�I|W�V���eN!����I�+{��:r�.&ǧM2����Mz���C��d<?�y�n��u(K���c*j�:ʥ��v�^��S���$i�N�JE�\�H��t�̪x"�{��Ky0����yz�?��R�6H��Q�����B���
�T}h����L��,
=E�>�j�6���Qa��	��[�#UG��i
�������x��4��l+X�`��W�^,|�S�_�y�+��.��N�YF�֜~��R,��KP�G��A)؏���X����>�kd�7�|�����~��NUn.(��z*aO�(>�VDޚ��߃ũݱs���S0��	 �5��V���Yhl�%�>1��#~��_`}oh|�  ȡ����G��ג��?z�c{dۻ���iP�4�ü%�$�}WkG��7��$�:*ӮG�I�9��m�B݁p��:z�֏Ä�gP=��L�S*x��yiT�ƅ��s����*u@�n-���|J���1��߯�!�K� q�m��F����h�{>�d��h��ô�m�f5����Ǻ>i�؃��qC�f��y����w��ِh*Zfq�n)�bR�T�L4x%M7�͓���0�@��n�C�̿4O��&",���Et��U`"4���Y)_�1��^��~���b/�<�_1+o
�����Ĥ��N�a�|���R�8���ʣ�F���z�*Dp�pL��ÎK�vr���a�[��:���0[�` ���E6E�%h��Y]�
/�3�\4�����4�s�²�O�*��r��P����2�j|q��'*X�#�#1�o�F�"
�<�z,�7�YӖ�hI_�mxݼ�wxG%��KF'f��:̅w`�sD�d�6S�
�X
y{vT~���X1��8��:�bn��/AY4�"��m���A��2i�"��f,�n�3��?u��XS$����J�*M��t5����3
���M���d��P��K�3�����Z�����u�>s� �[ぉLJ}�!1ؠ�<��pg��ȒU�%c�K�M�1�.��m>h;�vGq�}߀K��F������ ȐB�J)Y�
R���C�]�~��]�R��S����`�$��j����*�����1n��<i%%�kV�	lVz�6x��oB:��� ���p�L��LD3K�`)��^=�LEmGdu��nrn�x򥡹#kz*2�$�K�%뺟�n�ݓ;"Y}+�CY�glu����!�l���-�.��\)�4�7&/r��~����[2o�Sa���c���0�F��H��;S�p�ɱ�b`���n�$�Q�A�ވ!�(@�M����l�m��B%G�X���ɧ�=�kL��V��v���[00�L�p���Ni��&v�T�"KWl��}]�m\�vP':��p��kC&Q���Èb��ܣ�uʋz���?rᬸ��oȟHXD�x�݅����!>C�\"�YA>�fHѣ�{X�.S�u�]�ME�����j\Z9r(��q���ws��$��H�aQwNj���q����p��2LFɇ�k�M�����@�Ԛ!3���F��J���	@q�\�Ē��g��J�Q��5�*�lE�_�=C}�e��,�O�Ϻy�g�/|�1#�F�W�����9wG�A�ߴo��Q�xn��q��.�|nGX:�Y�,�mK$��0Iʞ����j$���Л���W<5zG��ߋpC���{�����.�8���Լ�z3�l�8����)���ONǑ0����&Vy�z�EC3[�	�X���&����1)e����dn��2�����wlvWM�wm�KUb��.�s�^V�#�sZ.�֙�?Z��Q*]aL��B��mI��OgMӈg��J�&�-�!�&>�D�k��6Ф�M7VƬ�;���&����B=��@W �1ԴG�����Eݲ���6g�j�PJ�_W<�]
�dY�7�_�ӔI3�8pa���JfZ=�.7���ҔN���~A(Z�J�Q����-q_�O��uS1+�S9��W�.��dǖ�W� �,�����Khnq��+�� |a�/ 3�V��0���Y�c 0D� ��s�ѯ���)_�������#�(��g���M BV�u��aX4���r[�������[�5`�e��ֲ��A�>�}��[�����H��vz�@#��m��0���\�iĻ2��Y�\z67�T ��-�Vʓ�/�Yۼ�QTj��򰧠��3OA��kT却@-�^0Ao�|�Z�ej^�Xk����S31��@C�x���.��NU,����V���}����|"̵�p�>IΉ�j�ED�j?�1��';g�v2�y?	
�Z(�ej+�<�(v���}1����BC�m��#U�\�׀�{|�Q���}��V֢�؉$ꚜ�1(kْ�qz(V0ˏ�jP-e�	�Ͻ~ZQq	p/T<�i"���6}mj�[N��!$��\�U�.��\�����w���}������qI;�;�[��	���/�����k;&$wɏ�%2NѤa�*S���3皂�1Й�ZI+��������6L{�_�0��&�Xb��W��5�]R��Ì��p�:���C#cL/y� Q�nP�OO�d�i�CHJGW/��s��dL�qY�=��q_*������L�`.�L����ʋ"K�_r�I*�s��{��t��إ��J0���?�.?��n��h�|D���co�!�u L �63��Ȳe��J�i��o�8����$<:[~&�+�/�,؊�]��&?l�fe�۠76:�e�8�A��G<-H�% ���g�H4)��Z��-�P�l���!���xl$�<h������K.�ɩa�j�9�����q�ζ{�b�P�7��i%���O͜HZ�f�˚ߕ���5"K`�
cQ'D���7��+`{8��'��f�B��݉f�*�W�S?|5ЦGJv;
K�L�+���P.���4�cp�G�v^SY|���H�">����	Z>��@7�8�=
����tb�������|Ŗ��o�~IO� �����<�b ����<=��!!k��M#��"��J�QEf}��q ����-�=�C�]~�}y��frv��"��G=MA��3���wm3��|�R�j�g�^�$N%AI�5�-��+�y�j)�Yl t��dpn�N�_�����[E���*�MhtA[3��s���Pb��ʬ������~�
�"�uXp�+I�|=�EG0�%o �1����Nqcc��%�i��C�f���A=�	zn=��e�Gl�v��j0�d�0M!����5��}b�q�L�I{5�⥝�����N�n�[�m�؍Pr�����-�o-����
��!�TX-�W9N�o��'�Xr�����8��\�i����x�C���#E�6���g)p �	@-��\_�iF�R�Ǥ���.���I~y���c���:@7�w�PB�(��8�t���ʴ�J!8_M��q��ҵzI|R/c	��-�>�j\1L =��d�i��n [��:: ��plٍ�~����!� /x3?�8�l�ڀ��٢=B5��Gr���>�O��o�v}�gʜ�it��	�/�]T�8=B1�G��-4�)�Q�Lb�v�}�1��)����ג��.����h��g!�0S"Nf���d�� �%3PǱ���l$�̉�����s��¡�(�U˷�_h1Z�)�Nbe
��/�8���4�Ii�d՜��w��o#s��͉4���W&}�g�!�Ϸ-��y�i9�Mק��Ku�����4z#��%G]���`椘�ߑ��񭥒���'fe����Rr�U&�)ό1��E'Mؿ�^@<`sa@���ӌ��}V�!����Dyʷe�'+)~D珡��I���vE�c��d���2x#�����f��1��ǀ�;T���e����ZF%�)�P!�DN�)��ǟ�o��8�x[�r��CW��u��ru4װ	Ѱ��� C *F�۔�F�p���f�٣����`����͌��[��Խ� ��12|ϋu�8~�yT%25!°M$���b��t>ҵ��d��Z_�h��M�!��OA'Jܳ؞�~���5;뵖�Mm�Dݗ/�=�:�B�x&�K��"�b�aP�P���,�6#G�;Q|��S�	���p�h@���X���M�1.�I4ܵ�K����T�z	��14E���q��x�L-��>��؉B��:\#`ґH��w�ۨ!�몤M	�.!�����p�֕��B\^Ao�����P�����:){#��6�KR5g�yUHXZ�����p��;�ν�y;XN[+��1�g���P�.�/�H(��͌�Ɍ��g&1Yqp���x-��NH��O�u#)*:�%���_���(�0�z#L06�*r'3^�����f�,7"�wc7KE��	(P����"�"S���KT(��gPU����L���"![M��*Hk1 ������I�m��e\s�ڡ��|>�H�v
2�`9t�F�Q"3Z$D�xܛg��x��-��q%�\�7uFӯ2�y���l.�F	�i5��H��S���:�Y�� bs�}�R��#ohC-6c�Nڳ�0��!�#�g��p~�������BsP��vh��K���{�`�f��f���X���W�׾�m��d�.����M.60���)�<g��<����S<ߋ�9{�/F�L�kT�$��	��'2ʣս�^9�`�����E����,�Ix������đ�2�%��v���L����pݵ�|�� ��sK���yv�����y�� +��|�B^g1�J$��b���������|7�ui�	sF�7my�f	�r�U��2s+�w�P�
I~_�B��d��/p���;oIUV�6���!I�	�1)���u�?�{�+9��k�Rد�����o/��Z"'����@�K����/����q`C���K��1$۝���Ժz4?�삎�ֽpT���>w���U����� l��E�W���i-#����]W���vh�'����_�w�1���R]��R#@��=[O�V�وN��^�Ì�ߋ*l�W$�V�r������	�\21��&�&�%p%�Vcj�����:�T��t� ������V�^�3q����A<�T�+3�糹jh��G��%�򇺉Oy����M��aF�+{���a���E�LR�P|<�a6�(����V<��2�����C���NH��E��N��H�$9�i;��^^M�	�0t�^ 70u�o��Μ���_@�2�CM��������G��:�wC㒤�dxl1ݥa����l�I�!���k�Rq��:L�; sL���yq]e0iJU9��w$|4��]А��k@0���+=4��|�p����%ư���O@�}��9�J�&)�;јp��x�9f�|���c�Uծ4��.�~��z�j
0&�z��/3#��Rk:vVl��!^.�*%�xǇ +����l<�	t��j=zf��0��ᴝ%�7������gQ���J��k+��DrOY_ Ez���v�}�=S�� �`N��I>'�Y��Z�
!
�bRG���Y��ޯ�� ͆n��J{y��Zq!�1���^a���|�����t���%�{Y@W�&�*h~U̯��K�`z���m����
WЁwl�65�S#�|�JAp��;��'M��IS
y�!tRGG���d����n5�A	I�&}�h�Da;�	���B�v��~�_�k�V�b%"� �d̓u��x�*;Df$hy�E޷��г}�2�t������aVP��?$Ԟl�ẁ��j��c9�j��#���'ψ�n���u�M���� Q�`2���q���Hl�����+�ޒ����
$�~���)��]�|�߱�3�PT��$K���'�~#����O�s2�eC
Ÿ����8����!�؈p�B��|i͈��)h��9����.�G�e�S��8��O��{��l)�zZ*O�K��A��=Bn��eKr!L�9,����318��w���4���^%+ϼ�����?*��
�вq����S��U�5;�R;�D2!#����G�w��E	��,M�`��}�[��J��d��_�)0���ՠ'i�+�m�=�tυ�p���ʛ���4ˊ0��_��g���Pi�%װڳJlM��Ԡ�
�ۖ��l�O�ե�����6�0�D���I�`e�6����n�N8D�;jǆZ`�?V��Dz����_8H�w/rE�0���D�(���}_p�T���C0[���	�����fh�����9c
T�I[�
���__���~2�c$�Y������F��-)��5Xh�n;:�/�)��;t�]�.g�9��p��:{'%g%�P��F��>l�r 3�����)0GHny���vEd��s y��m��"Qե=��P���\s�Hh�5nt��9�윋v�����I�M��q�aW�W�� �XPrUc�y��<�?�ύ��3M�v�؝ẈO
g˅e�H.�B�aR�^ֈ�*�,��3P��PR�잱�oJ� 8�47��a�&9�ڗ6I�	��x���+7rWr���n�5x�~T+�p��l5���`�ο��1b��� ���~u��^*�v|o}�G�N�� 6���F�M�����	���蔭�pH^GK�'�L��-o�ݮ Js�q�l$΍�����u3%0��Z��Le�ʆTad�;�o	 �8�}&�k����+�"��*涿}��41�W
����	��3"-�.��B+H��$�FA�H�xЎtI�ʐԡ�*��`21¬�umK���ǂF �!��5 #�q�N���m�z�cP�a���s��ף5��S��PG�N���ϸ���d0��gl,�g����\j�;���&Jj*�>N����\�Y�[�c��={[6]�Z��Xs�����d<�[���xQ�_���N�ua-X�$�t,1��VI!N�F/���"pJ��%��]�=��!�r��B��2ԃ�!���W��g���;n�P���ڣ��)�}�9w@�%�������=�C��3�t��]�}(��z]�i7�mP�9�E�UN8J䈄�k��E��u�:�����.�c�C8�W�.P�m��v�sl�m��Sp pІgiQA������h�?沔�Q:y��l�j�;hؗ�S��np9 T;5�D%��F\�#e<��D�P���P��,f\X�0͐�>3qΈ'fᬏ(9��)~OW,Z��J\m<��4�6��Ӭ��5;\��0�mٸ�u�f��Z��:3_c��s6�Hm��!�=�Z!f'�	�[�ԢE�Zʈ��)�B@�	��Q$泱�ȠA|	����Q��3z�|�P����|�x�}��)YE6���M�����40�����P�iu���b�^�V���L��ZXS����g"��j��K�y����'��L��y>��������4X�S�eئ�\+�h\F�Ȣޡ��'��b�g���ȏ���4�k9�j�����W�A~�Ť�L{�H�Wk��"A�I��mIo��?*�L������z�!�������a�>���Ƞ�̏�.BU�WZ���:?X��u� ?;)�bCP%�<󋓤X Lƙ�B���4A�KhK�c�tj�:����a�`�+a��{)�Z3��hv��C�V�1�dG�7�e@�������s�"�[7�/��qS�p�� ����M�ȫa�$����'��lh r(���C����Ҹ�n*�uU�`դ5b�?�8�Pm��"�E�-����3Z�GZ.�N���ң��z�&�����>��KT�Ȳ���vQH mt\��F� ���%���:(���I�*�{��N� /2B
	y����q����v��W.�u�~�o�w��=�R���Q<�>3�w��?Ikp��@IM��v�Y�2�5�d��d��\CF�,�!u��A�������x��T�4Đ�a
��UX��(Y�x*�,��=?��#�����YO4�h[�͙g�t�iZ�OL�y؞��b\��@0������O��0�@
�'`��?n�(oӹ�-_��o�0"�)���@�*a��2��yo�~������ㄥQ�O��R�^a,pqq���x�#b����V�7��鐯7����7䐴������&�\̚E��b���9g��UE���ü<��}3��g�[���e~������O���)}Ӱ/#dk��
[�K������H�q�գt�����<���݂�� �PY�1,\�ps�~(��8_�RI'�)��k�CK��%]��|�Σ�N����j*�0K�S�i�I��.��VcOM�zDB���36)�t&�N��q8��n�i&�g�2��Pl*2����
��Yceba6W5�t�Q�T��1�oL��"i�b�s7voG7951��W��\��"bHP	���I`�P��	�Y�R�2�0um���ڌ���i��A�G0v��܎#Q�Ҧ�8l�%`�
p��w�%@����
���Ϊa6���9��#IAWP�B.�v~l/��F��r}��@�-5���R������)#,g���m�9ݫX�^�'�f�Ϝ��K�v�ۯT�����m�ϖ����a�F�����nt������OM�T�����j[ș/�LdW��E98���Gj�r���.%�iJk�eZ1ܸuf�,�8M��D�q;�\�%��C����y�C��x��������K��� �j���L��Ϋ羂����ٲ�r ��)����ǳ��2��3�]�)�:'��Q���?���0�M�,GH ��'�4j�q�����Jd�W�g����-v���ƃƴ��
����;<�A$-���T��*�p�w���x��<f+v�j��'W�=zn��e�%�4�W��eŎ��'�{�/l�Mн���_?��
��d�L*����ՒS-XhkĄ�@���t�|a[A]�;����cl�W8bPļw�s^X���u�%̦�ښ'�K2�#�{v�^��?,���G}`Y��@��.Bt@9�ۯپ�cLtg��(��^�g����������1M��V%l���d���	��m��ζ)U�����
�ifE�y��M����>��&n�K ��οx�a*5�jVp���7�r��� �d^ؕFh �{n+��"1PK?r�� �k#���!������4�@A���G+�lյ�!���Ա+C��F�>⨎��1��*��)&��G�-�4n���w�3�!Y��D�Q���oF\�	��c9���q#������x�v�{wײa��wu-G�3��{(/	F�Łr�|A�L�#<�$����̖���E[tʙFeq��Q�隕J�;*�va�M!.-	�w��En���H�i'Aݢ&��k����$1�����(���Mz"i@i�P_��y�����R�<��c��|`� ��/���ޑ�EM�O�]</����/%��}�e��E�IB(��e���f}����B��,���o�q�g����3�B�pK)
���yl͂�<���BK`�������n�
R��m¬T1Vk�3Z�q�Ò�YUg:,O�����ȵ��O�><=���Ҍ]Uf��g���Z��� 	�\�BbU^e�=I-���!�L��C��fE+-s���#�g�WyQj�`�w�������\����+q2 �֘�U)�d�r%�s3�KE��O΢��Q��5��o	�͆��S*s��].�a���~0`�6lsQ�)*���7@Q'^�����C���>.�K�5�:˭?�0u��1���/fp�;���+��s�p���1�]܋#]�Ê���_���6�NP��²U���=����#�ץ�����t��/�ۜV�ҍbp��j��E�J(��L��:6�`��k�G�"���3�CxT�n�,ن�f1�l��ȂD�H��� &�!�@�ă�h��Ȉ꧸'ii���{����?}}��O0�S@%�D�*+ƞ��\��ғ3x�?�R�nw���!��|���b�݀al�@��J�j��W2�<G�6em}�<6�L�Fʑ[���[J��U~8���㶶���L�
��,���i�q�0�3S�ŷ�����=�掓/wz� t�٫�'+��r�~�{��L^�����k���N��"+���u����0����@�;�U80�|KH�&�V����\��&A`i	뼉-�W~f�teCX���!�yC�dn��\̈́Cc[2یHg���rn�	���	a��&��^gH`,�c���'|kGd��߫B�}�-W4�#��M!��]�%�K��z,x�е������-����z^Z
��|`�r�_���@��]G�a� ~�qvq�*�%��j���\�#�+Em')Ft��P)cA�V�#�{�-ܷ.t���K&�+��lʣe@��K��џ�[#���wQ�*�ge�[0)��y�U�/5�����_�4�T�<ֺ8�HSp#�10������|Þ"�>�}=�s��њ��O��A��҄bH�*�3���1����8 �m���Zbz!�dc�(� �yR��5�/�
���'��~l��V"[�$��~�M��RKh���w8��̐�\�P����XYSѿ��lhw��5��nj� ���:�ꙴl��([]%6�r����^��{��9|5F�692��]�jA��o��#<����紹O��g��Β6�ʭ&M��.J�=�`�8!J�%����*�>)N����2�_|Δ��W�WRM�������%�H��������|0,��dwg�6I��+2d�6�j3�1>�El���)aQ���1�>��$����!��Ew9����i�1����[9��cx!��9���"��#��3�~�n�:�m|���-�%�������1Kf}��UA��J-���&�����S��^ބ���%PK�k�\����c+4;��aj@p����� �!��dD��4���L�x%�m�sc9(�;��!�{X(���A�HF�O����ɚ�b�(� �KQ&�2��`�L�t�%��J���i*?Y�,�¥�	����G2R���Q@j����u[�5o&"��墂DCD�v���Dn8���+Q+ā2����*6�f�-��0��-F0�3\���mWh,
 ����+�\��f���4]m�x�A�5�Ӿ���tn��-V��� ȸ4H�3!U}��v�W��`��J3{6��4���fU��9R�K�Mhs��Uz�q�g ʕ����,�}���P�,��x��@��ʘ��g�tR��8���"P/�l�&/K���Zk��l���o���:��-�{���Y�(9ϐ����F��N��p�>��(�A[[� ��xd874J�z{D!��e�	��Y��劾b>�,��(h�d�*�]}�.ǐ5�=X|���=��	�gw`����y��t_��;Qo�:7�k�ki��JQr�Cx21��r�D��{R����*��ç?#{����D�En��~@�h���j�%)!֥V�o<X��(�֜Mx�~|$���uH!͇��4��I�k��� �>��h�0�@�D���W���\���0X'��¢�Ahw�Us�?X��iZ�?���������w�Eu�%�[*¼��㏠�B�[a��o3�2��Lqi�(*X2���S��	�Q�4��L�ˊɮ~$.x����Wdy�{�B#�0��&�P҂>m��68u�/�<��2�KNA�:mC~ݚ+�շ7���8�ր�͑�.�x����l>C��]��l��(�&�~�u���4i�F{o����-����p�5��d�����JY"hM7�cZJ�E�'5��`?�b�Z�{�X��w�����;����zh��LO����S�[
��C�e������LBA�@:�����]��@�}��G��.��(�<d���WW�۩<zs��~	u�uio}�u�,ڟ~�G~(�%C)���3���9ȇ;o���D7J�'�n�G��M�&&�/XSt�->> �J4Oj�O��QXR��:̴������#�����m���5��� �����jo��Y��:3eS[�5(���֝��	��i�*>�J�# (���c���-��r�L�����42��9�6n�:h:��Q)o�7������w��=�b��0t�����5c�t8O�>bq�g���G����n@^��1=B%�L��+R�4�/wx�/�J�~�ƻ ��zn����S�u@Fl�"U?��I�F�9�������+}2�{�7 �saA�:�@�?B� ��n���R0Ea#I4I{y���'Z��i\�j.&Go$�I[鹈N���>[��\]M��y��p����=	�r�[ 0jI��s���*�P��yA�[|�N�O�+������zk>�����ƙz�n�ə��Փ{@[c��n_mH�Nd�Ԟ}�Ś�3L���MGSUD�݉}�g��5��g�-)�XE���"�ڢ"6t˰R�(���}�w���P/�w���ZkV}�{������ R0)r�$6/҅��͔�|�j��f�������㺹�V���(�./���e��y�5�q��wh�	�����N�)�I�2��{�vU@��H1+�W�+pbRi}�jav^%����ԙ�!r�52���v�

�=c�uaH	�Z��. U^�:{	Ϣ��^�"L
���bS�?�C���]$�T`V�Iy����{���y&_Z�sU��Njڜ�-�98@!,с�ӫ����7k/^��leT)�0"(�ҡ�x�f<\���)��	h�e��([ū��a�b�m�%�;�3Ik-#�^�("f�}��Kd��2Md;~��I!�v�(ſ�_�3"�;\cI��q#p�V�H�$����i�"耜��w
���6�vp�{�~����)7Xk��וB�&d-A)@��kH��F��}���q���6&LCa�>Ґ�jG�
� y����9��xʴ1_Kk,>6��S�9݉�Ϩ���WB��s(�����[P� �Z���x�`?�����a�)t(�6��6��mW�+��R�L�mi0W�WR�?���"������I��4���d7��W�x;Z��/\NC��Lqd��/��k�*�K��!w������;�Կ����]��}�oID�z�qP/�|\LG\c���YI��Y�3�٭�J �h���'�Tnl��6�kO���b�0��qvk�z�j���l�ʊ$��:�l/�9<o��Zaa��e�a9p�ݯ����7��H�]KB�0��]�Uv%�*z`bf5U��Q��S}.+oŜu��k>���dE�u����we	����J��m�r��ք�a1�⮻�!(�����9�B5�x�t�2�LH���$;ɧ�H��m	)~s�#�QG/s�j�9�k�8L�%PtͳV^a\��f�J�[��	N\7$0~Z�P�����C�b����{��f�yѼÙ�Sg5uG::)����}��g�Ι�Ư&v�\$�y?Ö��WE���U`څ?��j�2�!�}Z����wb��3����~�pX[^�vhj����"M�����>�8�#-M9����R㌔�bf�v��S)�[����Ez_'q�1� ��KϬ�L�I��`?�&S9�pf���֪�~QabZ
���j�j���)���M���0Y�i�0�1������52�!lY�_�3��m�Hr���S݇[�v#�b4����$^��xU���]����+��UW��f�7Yh�:-x4��EQ6���L�;0_�S�����ɸ�PI��Y�mg�����?C���9Z��(���"k߱<5D�Զ�q�İ�Pg�&�D��q��(���C��.������냬�$����d��M���g_��!��0�p]��p����F������@���lD�p�Ο�>J�{r���ԧ�K�v(�ͩT�P�e�c���B#�m�z�ZG�B�\ህw}��9�����R�Ѽl.��r)�A���׀i�5����P�O�������Q#�d�\C�)�o�Q�(�C�G�oe�L8�����t,9`Jh5�pÎܔ��9-$U��W�����nޠΈY�����o���;��=q[�ݻ��o��Z���:b��u������E=s@�}A>�20�r������>��X� @>�fjlY'"�p�"2:�^�i��᳠hAԔ�O��ł�F��2��H�_�0�����	5,0�'�xNK6��J�f�z���{PO�3>����P�q!D]�&��'�2'�T�x]���.&����PAըϾ�+�HY�������Hw{����*/����ȺGwPo�P�$j�`�um9���z� ��؈fZ��>��9ڊ�*�f!u}8���<���*p��rˑƨ�礋�i$�0�Jy缈�����`Y7�ۂ�"�2�y��&�e�J|Zl@���8�Շ��r�UL��~��&������[4(%��7'�+��tj��#Ox����s�7��{�D���!.O�ː�ї���)Ֆ�F�I����8}�Mg��~W."?�+$"��[3�Q�гvq���%ǹ����5��k#���	I*(7��m(���:���U*�.h�{����KF�xA�#.L%�H�ddi�l)�G���x�ְ�<��?�5�]���4*����+d��9G�x��s^��^�O}�����"�8v�`�x��S ���p�̊f��>�;�!p"��+��R�>8�7H�d��yWdkI���o68gW�aW��3!�>�Ҽ��[�|m"�ϸ��YY���㒎$̢R(>V�/��g�r���H�t;�Q&	 ��3��jp���Y��kd+3�J�h(����!^H"[��R�κ���!E|��x�k4�HE��<�I�e� ��f�Rr��S���`����ڄ��Z)��'�&н��-'��!�K.��p+�9��eQ�w�G��D	k5���L���Q�aS-2�ҍ#��T� ���9��L�u|��C/Dv�Ub�B��zQ�jN����;	>�> Ul�SF'�E�w��~�*צ(a���F=��2��W��գ@r,w�N��H�J�;]h�DT�=~L���k͜��A�:��{�Zm���+̳���n�k��y�$�b��0��5�6��V�����??H������Tچw�h�����ivFs���[�~!�r��aO���޸�m��A��w���x(YZ5._f*����Cuv��~��D-=$�v����~��k"G��q��,En��z��Vx W�>�K��n�@���y��U]����X;�R�5��Xe����-PZ�I!	L*;�z锘L���-s<ߟ�b�YK�dY��;E@i�ق�#�.W�V����%�/4���`h��{�R�{�R��H7�n�+��Xԟ�:��l��I0�)56o�N��fy|Ê�L�����XJ��$��k�Xj�/<L��J��o+�%/�ȜZH#)ukp��
'�U͠�Џr#�lh�KV6 ��Fs�G��~4��Z��㐴Ӥz���L�%�=f���G@�HőT�aX���)@;ǔW2�S<�Zk}H:�uZI�(��m���	��->$#�yW��9�-[*~��/��4OȾW�R����Bt���{�k ��&�F+��H�q�3��g9X��~���&7����a4t��|��I� !a�����j �>K:�c�nL&JP�_Hc�)��p��ӗί��H+���G3NB.����,�9Tb'�*�n�G�sڎ���o�R8�Z�lk��B�[�����&0�밓����M�}w�[��ЉXri�1`=�7���4%��32Kk�sP�}y<S��.�����s�t�=��g��_��M�I��$��/�:�)����!;G8?���oWy���;R}�\)̝(3#-?�&�u���!E3�����m�MfQ�H�Ğ�-�`?l�$��u+�w� q:ާ�u�Ȏ�G���\���-��4��r�\���{�L�����h��D���b����9�h��u�;C+��"�ViK
�W�T�[P���� ����_yze`Dm#����J�<�Ҁc�����Yxry�5W"tߡ�O5g�7�;�[�`�B��UnU*��H��wq��<q����{#��!�.Vq�� Y�5��t��k��qU��8�e$z�M�(��)a��+�ր���yє5�@_�T�����ېg�'�� ��Gb���%�TjȖ�%(��w=��ܤ�͎���5d=׏Ӷ���̈́�4W�l�����ꜴבW.J�Qs��)FN�k�2�}'1�����z�ye�n���Mfc��(�S�d��0*���n*;��m�^)��$a�TS\tSHv��'#uR� S+r�Ec�!�&Ř �Z����%s��J�����6�Ρ�Knh�5 If�����ML�&x.�ZI��		9��{�|u7���@�G�4<�Op�&f�x��x�D���eP��iô F*`G�`uL��}���!ů�|^[�VX�N�MwC�
$�g� z��->t���0�R��S�i�J�:�fH�-��i�f0ܷ&��V�^��>�7z:[���}��71'�5��X�ՈIN����7�.QJ�$CC����NvY;-B���M'-��'tsKg�|yr1����N���K�2�Zבk��g�Ǜ��٥lH�bY��j�ߕ�0j2-B�FK<��t���`Z�ri��L�7���`�}��ϰX	��*�Q����|^���IP���c���`�[���r��ne��#m|�!�j�Su�/a�'fn�+B��=AgJާ*\������_�KԣGb�E�1�ؠ��p��hg;�.ּM�`5{��l�TO \�ÿ�̔��`�Q����ʒX>Cs��8����IΪ�����Gۃ�����4����YM'K��1p����Q����z�W�&b��Xf
 
"5�"we�����`�����
�"h/]n�J��¼�m��M��ū&n'߳Q���O`�<c�+ ��T6j3ͯ �2񊼐p��]�-�p6V9}�V�H���(T�w^s9�c��/;Ή87Q��S�zS�jOz���Do��e��C���e�]� $u�> Y�u�a����G�͋�גZ�NwL֙k�7$�����!?���4�
}s�������bk^oɂ�8���j����T�\�]���Ƭ���
~��5�쏵������k?����2Bl�������Fh���W����K#l��p�oD.��|�����E��0>�� �9�O��t)bۄ)�IEWM�_�pY�N]ƸʤO��^�m�G�����P���+�CI��5�J�3g0YŪ�-���U��a[����zu�n�C6���ζ�=d��ܒq�Y'�m	 �A=�0��G��KS��kM��B�M���O\Ar0fM�����!*�Xv��m�<�Y�5���`�M��~��1l��w=g���ݸ��Y���C;r�4J(������n�1}V0�Onc���*���j�DE/z�,C�jn�3�RoV��neYd�����r1<���ׂ%�B֍�sR�>�o[�8 Q����<dSGu�<��;Z���ܤ��7!N�;c0����{�(Z(';�x@O�l«��Ӱ�{+Q1��j�B[/�TP�^�:y�vU^D���q��{�����j',f�����/y{�ڻ����rݣDqE��C*3�
b��	���dE�`�k�<��X����T�k��
y8.@vU�+��E�[v9���k�[P�m?��N�嫰�d�YߥcQ�i(� �¬\��B�Rf<����R��A$�S=�0��汊�ĺ�E㭩�*TW9Z"�(�$I�~@�@�}�M�,�cB۲���C�v�(���vz�Z��i�_��]8�+^wN���=��LT6�C0m�Ѡ��΄�,�w��Zn�w�r-�����xhK.7d�	Z�8�qg�����3����l����/z��#�K'R��Pd�(�����ɡ?E./�#�E����o��P�/{�g�\��1|���B�.���/<���Q^8���Xz�4{���J���P��d���v+��GI�o����x&��GГm^5ڝ�����H ݝ��A'��?�i0L��H�(�����58�o�Y�'�<h�cJ�#x�'c�v���+�%�M�'�[9 �W9����U��M�:P�30\�a�ém���^��*V����G��-﨡������ݻ����'��ٹ�cP|1|z�-�Ի��G	��I�M趜��w����g��4g��삂�9�a��Eգ`�^?r��CȖ~�m�~��l�p��)���3����رN��c��Wj�����@ٍ��0�7��t�*L`��E��o�x��u��8ͧX];aN����6v�1�G�Ϋ̫V�yZ�<y��F�0�V����ε��-4ق�[Z{ǖ�.n��mw���zI1��jJ�o� 8<�t�P`f|��ʣ!�TS����w�i�@����w�>�p�	$
oV�c��ݠ�q���@���S�Ua%X�L��Kw��T�B^���,�=�v{����g��*𧠬��&x�%�w@yg�!+��r'bS��Z��.A2�8�~���g"�wm���eP��)[���Ӂ��y-?"�g���������" h��6	�C�-�M^B���mB@�(�DG���ſ��R���b��^�<�8T�X�xa�螂����`�.�_��X��VX���)�]���q�|<�87�)P]�nw���fL� @�?ĩ���FK]���ⱝ��c���s~�v�Y�"ϙSk�s� �GY׏�C� ������j�N���w���ȕ	�k��'������u�w�}J�Μ>��ڥ�����bA��{�0�m��r��@N{�I�M�\�k�N̺��]*�G��C�No޿v
z<h���o�����?��lNy�JB�ge�F'�Yps�� ��sէY.Y��򡰄t�|��/���3e�5o+��	�A�9����w��6G��-�3ɏ��6���j>���vD�qr��#c@%[]���p�K>x/)`-R�nc���P�>���1��{5t����IW�?��d�@�,���x��BG��ޯI$���J{CY	������[w�3aQ�KŗNP)�t��$�X����E�D�����Œ�mr`��J�}��(5���/*Ԏ�s�Kㆴ�����F�e���89���>ɧ��L������w_�I�ؙ%�-W�-��qJ͉��K����usj�O��&�ވTgwd/7�F.:V��U�D�m@����Yx��%��TrD'6{VHgI��Qf�/�u^^����|<q��
����35M�̷�����fO{�k�ؽ��L������R�Ym�U����D�e:5� �T��	6�����Ԟ	):
�B
���_�F��ٸP{��=��5<cY˝��=� �~J	��=ji��"M��:M�}NQ^4������xg�=H��Z+S��B�i g�֋�|�x%dgz�b�ww��Q{�x@��AR��� ���+V~��l!&x/1��ܐ�*���Y.=;�S5x���xR�6w����O��{�Z�@$i�pw��OaMkg�})x㎊M��{cI�k�&v��'N�c�߀hO��m(�W�Dg�v���:^y�kcs ��
��>*�r�"�m�n��0{v��X�g�FK�idv��st��9�@�@��T�>���K������@�z�4<��r�|�%!�1����^��wb����K��r�R��m��]q��v�a��u�I���ⳬS���Y��I=���|H{~@�[��Fy�X©�_��{��Ø|@q>�ysr��g��K��P]�*�B)i�@�ҭ(��g;�)�C&`��}`��6t0��1�cFl.����á�L�֩b�I�����V�MU�,�wlߚ�"�g�a�\{�Ǯ���ϟ�B�G��P��>�����je�O�B �1=r,�z���bWO�2	��+� �ո\����*��~4���Bl���(��J��|zH芵%}�_8��0�"V/�� �7[}��'AR?s�r&���]%Sk���P��p+��G�7��z�l�j�6h�HA%F����n�!��tX��z�C2����V��C��@�������>�ìd��	���Ǖ[m�J-��q������z���Z�i��m�E��T�ڑɒq<��	@�(�����١�5-�:{�7�b�^��Q�x?��Ї�\I�lF��H���5�C�8&���՗p����,�:e�����|u�{�w�@ }q�e/�@��4mIh��)%���"Zȵ���ve�h..h*j�h��D�7"�����<�4c�й�o`�z)N��p�%">��G��U��\%�$�R&օʊ���aS��$*��;��mBm�/��YMģL6|��4�AOn��7��?�'@Q�]|��s#����&���u���<˷c��uj�oK���G|���C��~�&�؋9�M�[Q7DGOx<< �gڞG-�U"X��*��{05ʒ�~#[X�F����r�����'�Q�lN�D���O0��zh�"�>Z�0�_M\Eq���Jw)��z
7O�k)d��0<�NO%��-�&��}���<��xI���Z�]���r�n�pw��?��-����a��0/���а4R�s�È�8��tUS���Ļ2�9�N��;����8-[ai(jr=�$�%���2#C���>�� Z:���u�G�.y[)�����2�:��oʀi�4�x ��>6z (��z�{��:L-����\H���Z�O����?}l�mҤ})=O�S��r��CkT�м}l��	�Ԅ�{��~�wx��
�)��͓a\��)j�5'��U����t�Ήa�v�q�C���|�7�q+��@L9ֱ��T'���K�!���%Tģ��DBw���?�AC�Ca�]��W�?��P
|�~8�?Tܼ{�I�ŕ���_��*}G�9u�`�9�y3�v��_م&�A_v���8�T����^V������R�L���?�Ѿ����o�U��,�����8�42Sy'�,:��������S;\�9Z�{��_�n?��h�=g��:�E2ӏ0���I��?ߌ<.�U%6�Q6^�����v�Es ��4த���e-�������'n����5�pZ=.M0��-���Q|�D��$H�'�� q	���y�����F��u��l�.�D{ֻ��0�:k�xi}&�xH��с1i�c��z�����:�ud*���)�X��?�/��.���~�@���W�px��`;��>�&/	�I�c�ۤ�~;�Y4O���'hUh�]uһ֍7������%E��i�X���6�U0��p
4�̐Y�V)����F��yA/:Bm�1h}��X8V�<{=]d�F�&����3�3����� ���������C�،�C��ҘI7�Y�DVH��q��$G��ȁc�˩�VS�"=���Q�X�K��H�ep��@7,�K��Cb��']�免�hsu�|��J�5v�*�_�@&��=�%�[|1�ھ��K��}kw�0��������,Ҋ#>-�3��;����4�upЃ��q$��蛿s+�?}B(Tsp�.n��r���sN�5Ra��(Dt�hW��U�̃�(��Sr�[�U�U��9$��J/�Ed�'j���k����X�t��kq|'�J����H�M�'Q%���A1�۠(�G�)oN��~�f�zdV��'��@S�9�)�yZ>�{���Y{宽֪:'��,��R!�{��KNe�[�fv0
��#�qg�m�8��iֺP���{z��Iw5fAŹ<(g�r�P���#�:EVXGy
����-�������6ށ�|
�5�4ٚ� CI���֮Sg��-�8�lƋl�\үeJBb~j��Q�-?�=u����!��q�.\�_:S���t{;C�1��/^��$+M��tX�ʱ��>�=x��}��FT�Tc�hn��&��a��d�D�`��~Rw����U8ԉ��l;����$��</I8�<��Vk�PMZ�K2K_���-S"��f�����pp� 3�kd�i�OFk�2���0[	�ac/���a}.&y�� w/B�̾���QE��'ё�f������-zz��R�E�wi��9@�Z5�U�j�2��E��lrVN8�D꤂�������y�Y���e�	6�ù�>r�)���Iߔ8���o��v�ꆜ�D�{D���z��3C�3dv���I<-��d� ���O}ʜ��yŠD��J7w�0�'�Ս+p�"�^�>Ҫt��po�<���d��Z�����g���v�<=%�����G!�'u���Ʈ�o���wђ�̼@��]��X�֔:o�D;�w2~R|�%n����kȦӲ��{:�k�\�7J!6�5�0��԰;5u@����&����v)��|�:�d�k�O����rs���l2Ǡ|�&�4T��o���g-��ŀ�]rT�ږj�
ܰ���_]+ńX�lHkTkj1��(�Yy���	|�{"�ʧ��;h=}���$ْ
m��MC+M�$my'��ك�`G*5V ���؀V�
�8m�A���@ch.<Cy�{�&����_�p���+L���Zo�`�5�t���VN �}���������d��=�i�ƨ�����/^�U&'.���W��S���v���L81>Af�i�& a��Dfv�JT�骲�J��ģ��%�3o� 6���GFKjt���4��*�̾�W*h�Z8����Z�cJݡ��l
��̄�`��M�$U���X� �=a;nMVz��L���̇�$�^�s�_9�K�����C"�Z@5 �9Mր=mλ�3��c
b��������}�{k5��%�ٞ{O��z-��@J���޸'I���(�+�qrw��u�'�fCF�y.tQ�V�Fj�������B��6�u�=�V�]�"��"fJ��{��N|��|B����F�+�Q�Oqe\=<��*�b	�Β3
�dy��I��!(�G��y?�e� �!:�ĥ�����o<�U}�/��,	�|[1v���4� }� �NLO�d��t�-�m'����&-Y�!���%����f��PY�@�Ǆ_�_:]�u���e�jd�F�H�C{7�y�E�����P�;.��������ߡ��7�Ō;&�_cj�u<�eF�����
��̃��W�q%27I�I�#
�� ��i?���_��<�X��CIo�H�����-f]>2��&�U������{X	@�LoPz�\�4?łɮp'`�f��,��V�]D0�d�
�n��#��~���m�k��NcR���q��p����ޝ��j�٧��s��F�����'��� ����M�Pk��%����f���L�@��e�JRI�x�U�߁S]�`�:؃��AެU-#�]� ��|h�!�b_�����bo��-PO#dČ99B�%�29������;|��[�f<�����f����#��
��mc�iH�j���jZy�u;��P8��L��L�Fa'�!w�4�m:����}��44��"k�Hlה�K 󚜀D��$��+0`��9��3�E�ߺ�V��rp�\���֌�������.B�����k�Ҍ�_
Z �;�sH��*�J�\�o����T!�S�ߤk��݇�+�௙mp�r��d��R8��V�n���>��ˊCU;O�Jp}=(�;�(�^+�~ڍ�𳨤#��M��~ʉ#���P�(����]U|IِT���Sx����G�9�A�ǩ�l"��jY� Pmr�Ƥ0N)���1����!DS`Y���r��ۢy�c��z}9\��H
��d"4L�5���eG�bi.#�Xt�w<>�� �g�� N�fh�Yz�(�r���do�6�<�P�_�;��J䱱\qˤ񞂆A������`�(�%�?�}E�R�M�^Y�7i�'��5uY�q��{�%J� Pu
JL2��v��"|{Q�!��=y�ߙ)��4����/�[�`��P�ŨD�X��*��B���ׂ�O��?����(��B�[�=�����u�TX)[J»(�������Y���q�	u���f�O-��t`)��%_�'\�C:��4e�?��>�����kv�b��ץ�L���J�E�dw�7��v*e�Ȩ���4�HX��M	+�d]tN5�/F��I�EWi��㣧L�Api`�O!�*�@2{�V��k�VhG"�Zf�]�9���^�z��ME�}�|��!�����P-$�h�P˟�lv�U��]%h���@�eDmq3��47��O�� B9 ࿄V[a�� �ܮw��{{TW&���=h*04�WT��sso�;�O<.�2����E�]Ь~�_��s�7b�m�NY=&�8�v���Y�
�A�}��]��K�k��r70��� F�����fVI@]7~��f�����j����a�V�i�W&�6B����D�1c
��)��5�_�����������Mj-}��|��D>{��%N|^I����-����W~B��&�:�
�tZ��}�)��2HJ���X��?�U(G�pu�Mt�V�}W �3赵�;Z�.~:C�y#%Ƴ�_XѩA�q^b7�w�~���p��sc"�ٲR;�;����׼���~�����f�sQGo6���rR�G�A����]���%����Pv�7�<�=�mǒ����a��Gk�ZSQ�'\`��5]BNA�����A�i]�!����FԴ�2S�!pAS�xdҚ�!��?�f���b����	ctT�sbM���=	��پ�_-噆MW���$��:�S���^�!��վe�>��b˱��τ�XzHb���;8��,a�s�,;����IX��+*��=*�4		zs��9����B :�Bƫ&~5��)>Y4�.ѯ���u_kӲ�Őza	Y�0b�]9�.?�7fG	�%N��df58��h����K^����Ɇ8��EP�=g��u�c�C~k��v��0ɓ[!�]����Q��u>�6���*��ȃo״�M0OU�������e
ڙ������t�v�{�:vi���ӟ��w�-�D.����XP��W7RX��H̰_�T�u�n�a�1�zr|_i�Z��qa$�_�Aج�p"Ao�;�P�`|�!��3W�y�Z��Ԃ����N�-�E�F��ku� �E�>��ǀLcV=>�iݛ�����@m�<��[�L
R���qEB���?}_3�I����� >�b�r��f���憧%�b�|��ٍ��K���k�;�!6W|.��������)�`���UfG�S����fy%�O�	��*���M���������<��p-~|>��T��e-���Կ"���\�~U(,f?R�O��M�A�8���8�9����bg{�T<��x'������1�4�ԇc�P���� ���|��?�BK�ad/�-��ž�G��/Q�4v�x�K�� ~�\��5�m��a�4+LD|���x��}ͳAy=��	�e�W:�b%���"&��d&�W�v�B��#�C�zj�t��1f�PI[�I�Y���k`��ͺW�iX�5�to���p5ֺ�O]r��N�l����s����A��Ki�s�!Y�*S
ʹ�B�����:)o��yv������3����K�.�$��V�]خbQ�M���i7��������Qz�j��ҨN#��7(���O"=x�Y嫞��I[!k����a(<�әO����(-��7���M֣V=X`j\�Zv*{k��'�1}I�{�w+�>0�:���?ǒ�#B ˺��҈g�����$}��%#�ƫj��9]J�9�/׬f�?e� 
�,�_6��~� �e[`��)"�����}C�������H0����|m�X��҆��`P?"�^"rp�_kI](;��������}����z���� �5��s� hc�A,�7x�s+q'*>�3�� 'b?�dw��;Z��M!�D�'i�'�X� �]��������G�ɢJ/��(�H:�W�'�x���31��Ps����6��^nN���|���H�B�*G��|1@��rw�U*�L  d�B��n&5,�/)G�6�S]R�e���W����!BUo^0X�/�4Ͼ�l��we�ܠx��b�� ֺ, MƖ�M) ���	j�dhG�^l�_�ng�%J�i2�`��w�0g�~$���خ�a4�Pw]��݌5�Q!l �+&�p�mȎƻ+�s,M2��2pش0-�IsYI�4lr�|H2�H����c�
4^\O������N׶�"� �
£TG͂8�k[poL�߇��6N+#��P��u5������!��?�K��� ���lm�iC"�J���K�DM��,^kQ(wr�aCcyt��h�xo����6��,���]�Ν��	���x�~�;��w<z�J	��?\���0�Sz�j�\���<� �)AY""�[[�J-(��	��ҷ�̹uM��(��V^u��+�bD���M� K\c���wb�t�z��7XԲ�Vx����Ц�@e
E�N�*`�Y��.	Ϝ"F��''_ʵoS���9�h���J��.V��:�i�^�	��4�*;_���l�G.�,� {��nx�������M��(�'uc���]��+�SWu2Y�9k���(��PC-:�|�+z<-�W)CH��՞ذ����I_�����,`͓O�ζ�����y���섘�����pN{�j���h�Z	?�\�g������/7}#�@���o�Ťa{�'S�.-�S!l��Nk�����z�z�2�������"��B��#L^��,�  z��+��#.�_��1L��wO�o-��bzjŢ/E:
��.�Un�!3�Ђ�jO|ř_Z��
�",d%���l���p(K�g����1�4W �
;'�Y��I��^-l<�Ԃa�^�p���e��{�A�?�?ǧ0"�_fI�9�����?��S��ؘZ�}?q+��T����v�9@ds	�z:�[P}�O�:
��0�D-���<ןڸIR��5E�R��\�o�-�ͫ����I��	N'˺k�d:�K���De��xR	<�w7�Z踶ъ?��,&T�{Ag�܇6�!���~/�����R_��a�u��D{~f ���X2ۏ�X�F_���4>�U�����=�ߥrݏ��2�Z6�W
��3*��w�G���mcb̮%3L�E�1>���:���7����g���״<tu^�c�~��;+��VmB�OTq����(j�6TEpR�-u��*�A��QF+�ĸ�b7����m��@D����^�9��5�������������l�, R��5�0�چa�Ň��3��Ysګ�M]a'u�E�}��ܣ��e�.>La�DO���
������ҕ��B�f̺�o,}��N�N����y�z+�;m��8�A3��iĝ-�ŦQ79��G���a+.�;W��R��5��|Qu��/�*J�s���^�� �����y�EJrL7�_Xh,��	߮Y&]��.��_�n�z<���Y*��ݾ1M�sW�<X�7�@je�;~e�s%���N�uG����[�f�6����Yd)���������8̑��)��w*�����83J���n�#Ȯ�Б�#6�"ĳ<'�PK�Ѫ���j�S���ö��
�ZN}N���L�	��T��2ժ�I�NK���߇��j5��i��Ӌ����k1_�9L�v�Oc�u����=w��U�g؈�q�(�cM^v�z�C �VF� ]	cK���#\��&ԝ�������kq��Ί=�rǎ��3oY7��\cU�G;.a�U�Y�$��'�D��:"����9
���t�P��Q�dM���rS�a{w�?&���ꆽ+�����b��wTQԇК�ƀ_Bd=��aɬf��s5/1_����d'��RC�D���S�^�n�釾Y�V�	��#
tbYA�H�X�9�9���̋|�<!Ћi���s�b�߄T�m�0.-�џw�� Z93q,>�r�B����!c�Z!�.���K?]՗�%��V(uS����� r�J�ͩ�=3�������KH4o�wϤ��ޓ��;��!7�:}��|X��%oMikL� �o3ᡀ��>�(84��'�8[x��r+ �?+���}��
����`Y�c��
�|4=��%�A����/�-)$)\�%�h�i�ĕ@M�X҃�T�0��:sg泴?��:��ZJ/�g�&���w��ɾ�S�k�{wM2��e��� �:_���ׇ��B�){����>��-m2p��r.�p �q���m�K׸� �b�hobt�����}cIi���Α�����L�,��v��N\>�:��$[cM�,�X�����e/���*�_AG��Q^�-��Y���pxd5�l���+eS}�畱�h�eɷ�ST��gC�$6��Uj��9 :�U�@�)���6�2߯	��MJ�����~�;R=+Ct�{l~�\�}�x~o��Xӆ��6=���9z ��2�X��t�eJ'��;6z��[�}K3��X��>�+ՇD#���rS�
S^�[����d;lq��~�qdR���΍�Y�%�L�y��x���W���E�FW������Uu�G�F��5��<� ��巘� ��������BC��orz+'g�\@�m,nܫ�~9/��l�T�j2� ^H��n(�i�uZU����v!O���4�;�у�=9a���
��u�� ������^+0��9�Y�
ݱS��P�pY���~7]�З����J���M��~Q�%mm~V�$��8�J�}�vkL1��۴<����ψҊ�u��蘓�} |ԴL��L A��X/��ju�L#�D:�?�Ҽ�1P�R��C���u빃��)��J�Y/��Bq��$f���y�Jj<?g���Z5Y�(B
Ҕ[��g����7��1��鿇�������$O7 p$:��2>`E�s�U���xY�$!�H���'(V� �����>9}�k�ġ�'M�O��KH��>�3��!�yc���>��y�:��1wߍ~Haǰ�}�X0PP��b�5�WTB^r7��$��M��8wP, Ⱦ�<���o����tCDNEzW+�nMz�\�T�"^B�����ۍ[~mqN���f�v.�Ju�m|j�&۹�㞲`�t����9�q��6�ԥ��d�q���������]RmE�^��pN��+��e,�&�"�]n��g�;��|�e�o�|��4�A{�2Q�a^�k�����8�zc���d�ުE_	V��`�&�P����F2�6lS�NO2�2�[���줯h��W�ZZ��]� �!VaG���@���z%`�h�Aܨ��d�Ο�ځ�F��q�h��؎���*T[+`��JK���q�z&���
/�b��ZL*=	�卻�%�̬����	��Єn,�,�b�xz�[jOR��(:�'�f�~v�4�rIc��W�rKI����bv����Ya�O�X�w��{�Qz9v�B j�Z=��(�^���5u��f�|��
:`knS{!�9W���H(�����4}�-�k]T �e�z{[,#	C.��W6�Q��0��sڶ��\$��A����Զ�uI�Tc�7�>W|���.����{LG���2P�[�M�����/T\,�>�B������@�K�9lg&�6�0rM��WN����* 5�fG�lE.��2�Y�1�'���v�cnC�v�֍��x��?;�L?l���ڂ͍= ���K���k]m[b][�!�����؝Պ+��G
��8v[R�WD�J�m��7�@��S���o���~��&�t�2�X���.l�U�xӡ�|!
�,�߳������*aeͻgr۲��G^�?0QS��`|�-K�Zʡ&#�F�!ġZ��j���𪊃e6D7P�(g���`�IX�i4l!�~�m��Ce'{���v ?wkp�*{��V%̠>]���Г�mR�Nʆ�v�I׼� �i��]��,�/��]:�LM��?*,�7x���m��.�U��3��s L��X*�IFO�������~�W8A�W���a��q���'f��lqv�8Z&��-�<G/���y�����5'�j8,1 ���mtN`�= ��^��=�1���2� �s�%+�?�B&xF�,l݇n}��[�����գ^�p��I�-�a� Wmè�/Z]Nۃ�X	��b��$�CV��_<fUtM,R��0J`A��غ�SO��X鸵1ۨ�!� �Rה��f�~���X����Lt����u�A�mYײ8���!�K����ڃơ+G��E>I �zJ�=��������ƻy�e|���F�=�3�������X����:@�7S5�[�-hOWd)<���o[���eeҟA�Q�m��b�g��e��	�N� �K�:Fa�Ԟ�5�.���)��|����~���=��������:�$U TC@�?\��(��q������#����r0�j����	1���ט×��c��+���f9�?C&H*����Q(	��t;�?p��2��We�f������ip"�H0��)���e��r1�m�b��	���`�Od=�����o0:Q�BY�?�E��a�����$���js�D(P���1��S������U�|����@]�M�3%c ��Ty�_#_�K5!�6�i�x�9�v��ЅMC0� 4�v�1�2�.���� .*����2���zi.�\�l�@��M�f���*�MԚhn�����$-�f ˂ڝI]�!Y}�����-�e�2@I��Fi)��;�P�c#��mr�)��b!ʲ�Pm�kӱ�L���$��c�L����YVFl*��np���-�Q"+
F{г�g�[�+j5A��)�V���}^�V':]���^��Y2zKkC�x�k��C禅e��R��%F�Hc���?.���A��vP�|������F64\듦��n%��G����W%�8��!�/�Sô��i�5���y���~�H�٩������ &֦�--��7L���5�C��JĢֳ�W�Ú:��.C,6�Ɠ!�w��FL��sՙUe,���s ,ԣ$��]�1A�@O�3������/��kU��E�ژ��-h����ҕ�WS�R���7m8���l6��r]IPɡ$#�KG�lvH�AJ�^�G�v��A�W�p�N���Y�W��:���uMIJ��B�;��mrNf0s:�{;Ղ}�C��
Az�T#/�Q��--���e':���]��@�er !dɠ��;.�!:�d*�������~�h<��~EIr�y���RM�O�)�M���R�_����0.?1���m9�v{`(��j����^�8�����I	���*'��Z� �����W�զ����Ȏ�3�_KAx	A0�Fi(*����$���U��7�e���e?��[A�]���z�H�����v<�z�&X^߾d��?mY�����723{�7����`@�O�5q1�޼���8ӝ.�,����.���|S(&T���N&��c-���D�󲋬��t�~�F(T�)~��T)��}�>�tT�����@�L�/��(�DcQ>�R��t���dCְ���/8�����~t��N���Ѣ�������0�@L2��)��ԕ3�S���Z=�n���t=h'��T��Y��ʑ����t�L,�+��P��T��dhw��M��t�~����8t~\�_�1�h��t��Uĳe~;D�����{SI�a�f3Z�[�L�n��c�@�x�9��j�l����)ͦ.����!.*L�7�!���������o�J#@��S�c~Am�lR��"��6�=��O�a�7P�,�ނ.�兊�z}�̌d�E$��v����x����T>~�2G�h�t�����P(�^�S������1�`�}J��$+��։�}o

��8/������ޥ��3s{e����w��i��σ�KEm�i���	���v\�O�ɺT��Ĉy�ʡ�@J�[=�%k��Tv��y�[H=���Ex��?C=4�f����.w�٪F݋�cPӦ]���.<�\{��
y�Kː��S�P7i�����B��D6�O��+���<�
�X�2��E�f~����u4��vD�{ν��W7���}\ɁG����N�aD�0�>�� �T<�C+�L�hQ\� i�! ��R���C�E�,P�f��58��?��0zO虏b^�M���J��>L��1�5Ulp�X�����[Ͳ�E��g��˚+�͓���8�f�L���� m�^���OJ��{L����m��C ,���b�����9��q	X�����3w:[���J������Uh���z��t@c�^%�le��D������VK�ꪇ���鋡�Ћ���F�$%7رZ{\�#0-®\?�!\~v���j}�g�7�� v�Z�Ox�L[˾)��Y��f!�+(4`d��D
�Hq�6m��:{�/�nD!�i��n1B�Jޒ�3(��JOݍ��Ş׆�����a�@�T	�t����h
_��+la1YNQ�]R�m%��^d�h�4��+O׋�-��C���A�Z��v�R�z�7���
#����G����v�����Y=�c4`������Ȓk�:�g���g������p�&֭���b�N��ҵ�o���o�]9��ŏ�0�DxnളL��-��22���-
�]�G���)��a�|P�F�;��E�[�&� '���-t���+�DF��_��*^Ֆ� ͷ�q�ƵLh,'����i�L��D]�%��\1܌���:�'�`�\?.{X0z跹ܬ,�=����`� 'O�;)tgS��雳�Zշ�Q��y�/���eѾr�V~�P��l/h4�ݫ�j��u2��I�{AN�k�Ņ�lC�v�=��tV���D>,��k�W���lv�Yg*E�ÍY\H@������vQ�ovLr隆�(C�g.t"u�H��e�+�������K���t�5#E�q/�r��f3{=g(������Ȼ�!�Q$��,��s7��0���Sx��v�H*����4V*�������SS��;�fh�n'�q��=��"�����5F߂�bf�������4h
C�M�y�cimP��#��t��E;���&{��HC�#��@��lNT���d�a������ �TY9Q�@��Ey���7t���gbmV���;�m0�%��W�+��*�	�zd���ީ�>Bh�H�9�@�~�z\T.|�E��$�}���kc��N�;c����tGJ_�ؕ�����{�rD;C��x�<�����N|��҈P�2���h��(�&�[>a��}�W�"Kj��k�
42e�R~�f����bsS���>�[L\��M�_Z�mZM21@��B����-̽��Ҭ�Vb@��&�he���C��ƿ�i��*?��̸I+�[B�]%7��f��5�9��?}ů�����r��^��u� �%��#A���� 𔀜�J��1�|yh�M˙x���i�)
yp��N�B]i�~�l���;����8����0hGzK[�������hy�+���o,�h��7��"��ru����ns&�#2��I�/DVѵV��4_Z+bP�M��QhrqD���fvH����.�R
7��.	�c��&�^�x<ń������O�`Kx��4�j��x@�z�Z��[t3�Qt�+mh���S�nNc��G`W��I;���%��?��q��K12�=-��飁|�����@���V�(O�MWς��/��&qpF�<�Hh˿�|io��_���Ҥ;0%���+e{��vǯEBR>Q<�#� �^�葁%�ڸ��w��$V�c$��YdU��֢#�ΘI1a� )C]@��\Z2��X1�a͌"���˧���F3���΃��n������U��^��,`j!V��CvtW�h�wɣ�����8hϓ��L9�����X�),����G����L�7����$+�����I���u�����s`���X\�����^
��q�>�C��F�%E~���6{��/��b�ҖLǤ'g��g����J!����xZ��-i�P�ZOS;�%&���Oi��|E��دi��Oy��:��q��K�]��&f-n^���<�L�Lz�ے����=���@-��`�럥� �X�'g��R��0[/�Չ0�G��?_�X��|��薧,՞H�gs�cF ��KL����8��h��3��d�"Oy�K#�w�X��c��0�t�n�`�4P��+�@�q�5k��,�v!Fo�eQ���B	��f�?���+�{'/E�G���46_���Ur!=�w���R�i$.��Aƞ�g�m$!�*��$akkyL9��|#�l��j�h���:���I���E,*U<��9�YQ�����~��/��cz�L�Br�V3���r������_��~��' +�
�f�,~�z|>�|2��^:�H"�8�B#�I��R�1��H��E)6hW�{lY�@��Z���G�Nt�@�ʔ�X���6Y���F��;sʅr�K*�p����m���i_832�Ũ�2�īi]�B6��g����MoK�%�$�7�?�6�w�
��	~���p,2׶�O>@n�A`�ե�e����*'Dh06�*�R�nG�ڨ�z
�N����Y j�.	���J��@ّE�d��*�+qUG��8��wL�N��Ѯo�4���渆�]�)��!*ƑB �j����?����M��G�ڷ��^ⰻ�F	�I3�6R@�S,  ��<��U܀)gr��{7�8u�
l�|$c���'w�����L�4�sR�!	��5�䀥�l�Cm�^��ΨM��F�N�7eb�HҶ���e�-�F0]�J-ZS�ғ��UOQR�J� E�jb� �@?�c����X'1Snh���n����_Bڮ�h�E� k��`h�2?�B?^cʔ7� 	��#�'�|�ZZBO	����0?�~|A~
0��O���U���Y4�E�H�`l!���T�a�u�
KP�	F�\�'��4Z�t�Ad}Y�U?a_ay����\|�O^Q��obuu�x-�$�Y��>�Ԉq^(P5���Pi�!��7驳{�����!����Ę	�~��!�#�w�N�����j6�dX7�9bs�L���sdtg� �69]fpg�L��W��!��d|*9��E\���@S���2�3h�������ۡ񞄜��Pr�CNUnD|���4����Vs� ���K\Ӽr��s���>�I��ޙ������ؖ٘��z��&�V;����� �#,O^�G���qTĪܫbu�4{6Ha�����.%�o��J��2]��v%K�Vb�}�f�|9���5w!P�pQP�ӆ�黶^��&��$33���,��o�����G�u3����z����h�:���J
�l//�Kk8ߦ9���c�]��*��9�w���3����� ���]1&���$&�I&�s�� &Ğе�B{m��`t�hE���<���lb�,J��a9�����P�Z�I��靃eDa��w�o�R�^�b�쉡��������[Ke�4��a2
��Nm��x�\MZrMj%3;�&�j�*z��Ζ}��n�N��8�!��J���,o��M��f�{���Iz�_0fw�	���X�$7��� c7Ѭ4 ����{�	����xA�L$o�P���en'�U�k�J�KGB[���2�R���5/�9�&��T��n��΁wz|>�9j,A��Q���8ɇ�c�q�.�������
�*��"E��3�i�)_�L�1�Y���G�Wi�E̎8�z[2�!�O���J֖衃p�c'"a��8���������7��8�0]�i�n�]��ׇ
��g�?zl�a�����A܊^�Z���y�v���p��̀���d��~�^��1y5�1���m�DoP��G�c��5ǧ뼵_�S-&oD�.<�����^��ፆN[����ޝ}�Um&��e1� -��v1�r�s�]nBa����24���q\��8X~0����/���@[.����z.��Xz�jf��"� E�t��8JUZ;U/�ȫ������j%�3{����� >��W$�xD����f�6+6�*U�ȼ����}4%B�����s�y�#/�'�i�i��C�+�l��Z����3�z���MM�I�H��>w��c��� (�r�M o�@���"����T]���s9I�v���%��ɇ.�q�B����E*
@Xk��zv��M��~A�H�3��R��o?��d"�-��j���y`��+��Q�AD�&�������[�m�s���X�`bo��e�������r^T���"�E �];c������?o�a�Z�E��G.�ܢ{斀d�	��؊���%o�5u��^�rY��E�@mc��N�O?�c���!!�R�9���q��Cj$	� W^����(lT!Zc@�������p_��+ m�8�:�e����O�� �W�� ��WWꄜi��������"�2!��=G�o���@��*��6��֔o���*j������Du��0%�����UP��|1�_A*s6x��ht��f�=�E�O'��9t��ˬ���ۧ�oF�Z`y<]<giE)��
�Ú�C�,(����/�[_���_KV��6�Zx��e/�<���'םk���Pm%Ykjv�C������%�Ǘ�~ � ���Zޛ��pԍ���Ɨk.�#�+~k��#�Y�`��Ր&q�A��QB����S�J�DC�p����Y�n8s�b����o��|	r�h���W���*�Z=�(k������:�;���1b@*d|F�/$"��^�X�H�����K���Vܮ�����
³$s�;:!��-\t�;��=�|%�J*��j {F�:0�o���R+�]T#�Ʒl:ٳY���w	P}�DCò\@�>2(��'G�ݼ��#��8��a�����^%�_\c���,�r�����"�r&��\�q��mz�yqS��G����Q�XqX&���n���L�>�M'm���e����Pf�H�Y7����iM|>Knl��K����]�
�DNQLEw�Yp8~Ƹʻ	m��d�?m���Ȇt���b2\2W�����'tQ�m�ǻ�����,�w��8v�yD_E�G�̥�cC�|
'�V���5�h��*V���=�p��V3�.�0.m�����[׹6��{�[%F�s�8��� [�������oQu�FOֱbt��˖�&>�!e��0K��Q�H�k���0����{�(��?e��Tv��s���!e䘴����~�`���|���am�J$��hm�0r	�HRg�@�@aI��%�Db���ؙ#s@�;�O"��SŋƑ��_	�k� "ɣB-�F<�`":��Q1�9#��@aK��������^>C�0k�ò�H!$��zW(��c�Wd�t�b ��<I!���%��Z�X\�8ig��$;	�����Fg�5��3$��Ev�yv:8@�� f�S���f��I�ˏ��4u�{�����&k`��W��w�)���oL�I
���M�q[���-W���]��v���P���N�G��Pv�����m�P�Y|��|��'��:ɨa��[_�%.���r�����Y���*Ð#�n��R �Bq=����Bg?*"���#��B�����2�@�ԀA�\��H0��$�F,L��
���<3qO�5��l&}VVB�cͯ����}��.D�E� =e�"�<@����~�$C�64�.�z�j����j�dvl��s�����.Z5>��x⮆��R=}i��W�ɶr4�VLx\.z;��hH�&��c�-x%�.���e�:����됫#\�xi듑1����I3�F�bLF�F�v��Yoפ[|��'���R�J��Y���1K��Ώ(�Hh���=����� >�ʮ��S����7�U�����|pQg������A�x��N� �Pd���^��D?�7�)�D]��Eg�U�w�,scK��A�9Y�U.�xԼ�{�2q=\4��a�����4(Gb�� cM�ZtZp�T�)��3�� ,9�|�~n'0�ꒀ1���ʪ�Wx`o��H`fZ}����<�\���:� �*T
�V��:���Z���I����a��\�a�8����	��p��d�ZP��p�|�Nyed}�j[m���{%�/��<�k��3�L�=����e��d�C)�����U���>�|��xf��#���C��v���S�ök���ٵ������5(o�C[����TW�,��ܘYN�У&�Uf$��Z�����T�!�:-���rT���c�kG4V!ZD��V�G�d�N\��/<��؟�i^8��Ii�g�\(�_�W[`Y���QV}���3E$�}nI�V����m��{?�<�
%����Y�X�LJz���$��g�+�(M݇D+	+�z<��1P�>^~i�Dlb,�@<�z�
sz֐��V��⎊ȾTz���EaڷZ��|jF�`���1��=�S3�V��Āɪ�v��'��k6[��P����0�Ji�w��ǫ ��U5 ���)s�jѭ����%A�v`��,MO�[
�G[�^4=�HՊI�������B��0���/��L��)I��㗋,�D�"�g�Պ�1v��ܚݴ{��eg0*'!VN�֬��̦�-x�
����u8�$���5�C����)�
����7�Y�]qB�.RNe��i]�U�'a�E=r^�g��h1��f����ڪ���ɆS�uQU���9�o�����A�~t(��j7��S�4��=��?a͑��I�zi��2�-����R�@�4�%I\{�R`�1���@�]���:9���g�����Z�&7P�N��ۦ��͕־�Ű	�͂��|7�!�*$���`�O� T�r[��ـY��͜�8k��z��l��C�+���5m:���r���n�+��}?��.B���lcɫ�|}��m�=^j�����#ܵ�*���{v�p���J�B�;&P�k�%,R�zW��/L�J:��%V!�ay��a��	�0^5n&�+��U��|�1R�[����[^�&<�1�?�-����鯼�yg�z�5��^�bA���H�͵USj��!0c�#����	�P����k�b�9}N���n��qa6�Y�U�n�*:`�f^P�_q�r�	�:E4f���ƹ��hJ�%@�և�")m�g,�i E*� �-%hg�"�kZ���#H����΃��rԼp[hG�e��3���ӗ��t�Wp�M��a�ʹ�D����?�iJ�A�&��4d��z�H������tt�
�������q㭢49�󖍱$nw?N���~��`�5E�ݴu����־�ue��g����VX,t�C�qsj֬����o:}pq���ܚ(:(���4�|^C{���E���E&y}��j�����PD�\z4�]Mg3u��swK����+T�!����`(6[�+�5-�J ͎��Й1�@���[O���-�­u� *�
�����g�$њ_3���Ǻe�f�,ϞA���xK��`4�U�����V�
�E5{P����8�V+�Ȣ����|���DW>,��v`�WM&4P����Z���]M  �<E9z]�6��v�䎏����=���	����Vo�7�=g�硥3rYUb���:B8n�g��'Ea�GK����f>9��GR�(wdT	��@zQ�2I�)_^e�~v�4&~@FC�F���!#��I��@;Q���to��N��8��
��yhZ
Hn�S��5U�J�1"KVb�[�g��6����֖�1,�P���~�X<������?S�K����%t�2����YZ|��:;���a!����-D��5�ǵ��m���	�i�����5��/ܘ,�B�K(��;>� Բ��'F f
4W7ik�Z���@{�(w�GFM<td,���1G'�����|~ε!�E�����:"~��oh=S1�;mT�5�$��'�.��q׎��{N>"2�[�n�Wm���#i�b���:\��tl��RI�q@(��߰�*<�xK@��.�%D���i5a�cɝ��Y�����m;!Z�h�0ΉR��[l��pe�����;y���=@)�K�C�>��{>d���/�G��G6c ��ڏ-b�"r�h	���9�(�=|ȑ�}���h%��$�>�'�L��yÍ�*毩�s�B�}�{g�C1������1/�G�hU�X8d ��J����Y#�R��q�l{a�m�Ǭ
oD�}����k=<M��̢�?��1��wV��^��Bk��,ӿ����(���$�@�DC NL��D�0�����'ɩj�/]�W��W�w�@z�����e�j���x"	Ogv���ЂJ\��o����{3*>\�N%؞^ػL�DJ����>�HR�||�H��3(��v��$+���y�
��v�����{�1܂^� ����*edd�R���L��i���r�RZd��b�(k
�B�"��up��pX�aX�wK"��yD�F6�P]�g67����H����	^|5018%Zy��=���:!;6�"����B���u�G�q�}�ʸ�XDV�����;/N7"�	g�E:� �U����C ����o0��k�i?�*�h2g;D(�c9jΡ���D�A'��?E�^�}jj����Rqm>'3��?۟ЏR!F1���;�|:J�&��75=c��A�~�2�q��]4@�æ ��r�QR생��g�w���8Z9��U�
w.z��b_4C"2]����.�-n] ,��r�\�RaB���FDa8sZ���hQ���~6b[�U��NL�ü��'V��`?�hD9���U���l��47�$�=����d�l�5O�����^���,�@yX���;]�9��־A����N��M
iVZ�����(���h*.<��kh&�v'���i)�ReN������j�U
y�����0#��B��f���JTq�>�]+7�A2b��cg܈X[2��E�g�~�=�;N~��V���]L/"����d���bA%����:ݺ���NM29v닋F�U �!��u��3��δ�$�5]h1��L��0�޸Z�!}��ApA��~K[��)+9+6p��,�����Z���_�-�M���/1�E+���{Κ�+�/�!�lC�eMq�8�0�a�v	��rT��e�57��;ş+���R��p��ĥ����V�������<�rW�ɋf}�k%�?�~�
����� �Q_�S�l@�:̙э�P��Wf�ow�z�t�FS=��*F�r(�!�@�-!;3sG�����_�p("�sJ��nW��6İN����g���8���(����0�^����e�k��^���,�J��U4�r�b�pKE��AfMp�Nr��-��z50=�$�l���py�!!Z����h�ԕ���8��6�l(�=| �/m������}U�H��9��� ��c���������Εg݇�����)M��O`��4[
���&�㢷�=4_�-q7��w�ɍ��0��2{В�c��1��nrf|�*�町���oF�٧��6�-rRPlq���cG�^.5��F��qJ��o�]l��:Մ�)il?8И��d�
8M>�APX����~��1�¦:��'	�1����>���:��A�(�@�G�����
��J�<3"��;�WY+G��9�Ψˢ���A�	���V��-�1����IȠ���4�b&/��t��Q��Yk] �'� 4+�S�&�,w�V%�}9M|a#1�G���^�*�r)�W� (����=k�/��]0��X�����R��~�{��_q��ѝ�(0�p1�c^�~�R��>�ٝ��d�mV0F� ��Œ���ͮ���b��l��]\Z�J�t9�.N[��N�9*��!���0l��r<��WN�G]��S%^�3q9G�Z��%r$��B\�|@��\\hY�=�dm�?�ً�h��C��"&��s����p�J[�@ ���o�`��A�9����Q�s�`��z@y!c�xFoߪY�e��w&��G,F l�Ĭcg���m��@���
�%�קNK�����ڊ��Άn�Ԫ������X�;%c�R�@�E
K���O�M	jE��i,�o�6x('�'������h�f�ߥ��3��5	e�+�V���MuUs�%�!��8���X�*���a�э��q>�@3�*v�O��涙7b�$͵��1��i.Sϖ{�\���(�*O��ǝ�y���L�j+��k��a)��tB6wޣ}�I�t�.�Ǘz�h����RX��v>.7k�By�R��f�Ϡ���r�9|��>W3�f��m��e@�rZ�؂M�,&A��?��Z`�{�<�p�5�#�egx�œd�?��cL���&��\䭾*>�֑�W����('Qi08��[%�+�:��%y`S��xT�s�ح�����L>������<	������޲�/�o�s�.W��Cֺ�	��%ߓF�9�tc���k��f=5t�M����G�~[���d���ffF웻�Z�m 2�Ba�ǲ���^㝟Z-gŋC�4����#�dL�PF��!��G�ʹ8�}r-�l��>��Ϻ��Y�䡬|�9a�Yl�L����O���..�*������3�gtj�M�q>_N��M)H�Wڈ5w!�TDF�}Wl��u��g�̨�F�A���Ug�RK�:�F�a>�G�'r1T�#��)gP2�6���{d�F�`q^��k,eǾ\׌��Ƚ����hD����)��{��Z�
��ؚA��*�72? >\mXt��������dM�v�3�I$+�A��|���iB�mu�����v�W�E&xd�A�\������9&Xna���"xq�:�Ə,�'�uL���t���(��F3+z�����>�I��Zy-f����͌�r3�	f��F@i*��K�aʌ�/:.�r���J��{P89W�8i��*F��3N&g�9
Om�xA���s�?��l,H�4|��tǋ	����}��w-�Ï;��M���?9���WPP��RhC���A5�e�I`�T�����^4��R}�?�zn�lm�b�&�x���ɕ�|{�2V�9���4;LI��9�����(��� ���VZ5z1���/ݢ�#�j6 ��;?^�Łf�d�{^�
ķI3X֛�=���z6��U�!&,�+8e�u�3�SP�V���-�춱�&`1X�&�t4^��U ���o����4�����	9����W�h��X�.'hE�b���tu돭�`�'��/��>"��ٰp����W�ﰔ6��z{Ʃ��ok�
_]�k�ixw����{陪�U�R��g�����I��6�	^N.~�s��Z���G�{|�iDۄ�_̐qY>o[�7������!��̺��׺."�䧦$'P
(�T%dID�ȯ��Vo��j��c���e0�"�'��ڸ#S�n��ؙ�>�>�n�>���[M7'$[ݳ���cG^!Ժ,�A0nb1�XJ�w����<��Δ=I�����2�����^��4��m�C�UN��U���8�Ͼ���v�p�Ev0�X���u�C�A���a�g��OJ�� ��Ou�B�W�Vs�Ù�����Z&���(E�=��U�Q��y�L��(�����Ipԝ���٫/M2��ǬH�RG+:( �'+���`6Nq�*?����6�sC��̨�[5Ar߹��)��Ȥ������t�G��eۅ�����?����'mdM�G��f?Aգd2/>�lNP�ͷ�s�B���|:��;+#�7�F=hĚ.ޔ�i�T���K`�E�g��J+�CQ� ��f���9�m	f|Y<ڌ1Id>M1�0Vx'p�����6`c<���6A0�HR�^ �Om+��H+D�����R�c�rH���ܖ�8e��jL)$-oBek�'%�mLx��-#�7?lN|�����OQ��.�q!����]���f���"q�C<QP�������¯ן/����d�2CeI�2��T��'��ؠ�q">�7����BB��{Z��!�N��(� .Q�G�dT��5��1U��)�4���D ��D�9^A�Pڇ/&���>Ý��@�B�Iawf�.�'�R��E
�����|�&{���bh7��e�^u�����o8bu������A����q~�^4������m2�T�>JM�ᷝj���c�yD�f"���o? s=�_��z�ڜ��\�Z�ZT���b��UZC��)1H��W�	��6e�o"�!Y.SN����j��P�
s:� �.��zh�Z��*�Q�N��?��=��9:_qq�&R9���i�A�`O�y=�3�Z�W�l)fWT����TÈp@׋ϣ�=�g�i>��o��������K��B"���+��W7��(q4�ڄ������.����-��?"�bw�D+M�k ���jiE��F3���H�m�������?򛑸-?2_�m=�I���Nii:fY�X�m�R�X�Ȱ�����U��ɜ}���d�<��R(w:�$�~�3UD����`Y�G��E��og���NW��s<�9z��\�oA��zzb��j��R�j0�[3��� 5���\���ח~��[�{z��S���g-��t�A(ց�6S���x��j��7�1���ʂƉD2��\��QL*#Cm�Cy�u�������m�G�J�����i�F�}:b�4=�_w�CYB����b�5����*�X�c��Oh��R�z����#����@/���+�T�򌪭 #��jCA@%(��[������ݦ�{�����q>)�Z���ӯ7�oa�l߻?&eb�;���Wf�HK����S{�U�,p�ϴ;t�|��0�Έi(T-�d<U0/l����}D�zD��]	�dZtq�5�xgJ�mT�Ө�0�lM�H���R��+���Vn_�STbYcS�M(y��1;e^�6��uP��"`��g�(`�[�
�fL� >Y
���{#�s@�	���kq���/��ސ����oo,��?�EW��Kh+��<&:��,�v�/:��4F,�ߞ°#ZmQڼ"����m�*���_突{��,^}E�uO�\��,�+<GUӰZ�v���+��û9�r+,�ڙ@�`"��ua�s��l�A�2�}�O]�d�\a� !8�b��uU���>7Uq�\�;����.�׳��?&%�j�ObV.S�L��C�sө�{�_��iMvJ����mJ������6=d6�Z�W��&^�[_Q��Ռ�	��5F�_1��`��N��㽩���`%����6Z-�]uƯ��H�(�iU�B�^b
#o?���K ��Z]0�!|G�����N銉�SeԐc���qU"���Ӣ�Q��%�3��E�m�ۚ%>c��FӃ�G�l{i"X����U`�B,掭f��x)���yg.^�&o�%�f�+GUZ
��i���fX�?��Y�z�<s�mD�Mv�AA�p^aJ���,@����/�(�>S���ð���f�\�[G�(��簾q��w>}q\��I�K��k�V^~
����݃��+V��
t7gPT{h4E��W|�d��A>$*2%��_�N�� ���� ���R�������#�` Kffu���P�>+�,mX�t
�u������]9� � u]�pN����A|$N&��Q��*^,LnI�&�����������2 A�j������\�Q'�T�t���\��IUJ�1������wm᜜�$�D��~���cߚk�Hm��nӠ��8�c��Eg1��ON���Xl�'6v� �!{�(��`�,���XN�* 7�����,c8溺��o�M�쉍8�ޘ��|g4�M�Czm���|���oe���LYK]-�&���y:r%h�:���gIU���m��A�Ł�1�E.��LĸN�m�.�7���@%"�;�;��!|�w>����Y�1�}Ĥcǒos��ؖ
i�܄_m47��ȉA%��*�c�����b���(Hx\ѵc�ċI���l+���{�$�0�A=l�6������z��er����<�i�$:NQ�M���6i1��T�V�KNCT���L��s�`�Ӽ�=�']~�A�bF�s�= #\͑!���I�Ā\�8UL��{���E>�S.���-T�ĩ�B"�{J���Fp��&N)s�O����Wǟ� �8�[L�������}ߠ=[ǵ��Q����3%�4��K4[a������J!���!��$G��͵?�������zܬYH��K���8�9!��ג��,�v\χ}鑽���ӯ}�T��.����O�2�����!/��uL��������6|vdy�.�+��k�s�x��_�)O.��h�k{��ꖈC�q�h��	Pc�Ƨ���#�-;�D����I���g-NZ��C������{�;*:��8�C�pmؠ� (��|�M �\�3:1���#����E�]��>4ǖ�y�!���-�T������ a�h%(-|�r�\M{ʀ~^��p��9H5&E�� u w�Bo��M���Tܤ1Qs�!-���^��pe����*�vX�Q
������ �ب�UrZI�0��x���'�O�o�t�?��2'蠙u;s�`_�0�K��Y��Bv�e��ʜ��0�i��uz���I˹��� �3��k��ZqxEWC���w|z�X�|�v�M0�����#��)��F����"�.Z����W�"��&y�t�c�m�Y�o�ZK�'&{��$n�8cz`�O���,�J����<l&&^���0�������w ���Z(a9�S�\��SԬt�;"�ȓ����i�t��@X�k� �Q��#�
z�F3
O�h>7=�.s�/��x����[2F��l�>�Fd��)kD}�f�|�|{Z�Gd��l􌒙����Ծ�����^F]���Η\2V�eQ�"_�� K����L4~���`��`9S�\�ڹsX# 3e�4c#��<b�/<�rZ-Qd+M��\�)������	]ݞ�^x���%�r�-�$�w�4�e�Z3�vb��b��pO�|ɡ`�|�G;����ɘL���WM��p��֦M�ׄ8���yW�3�uܩ�l�S�:�X����0�/
.�}��7��o�ȇȐ�6I�L�\�����+��Q�I�i�z���	�jj��+��rV[����B93��d�Bѐ%|6�m@EaT �]�ռL�;�l�[;L�]���Y'@逻	��
 ͗ɮ���0N�F`��!OKq�<�f��c�;P�v��2Q{�Iʯ�S�Mz��pm�w=��H8X gI�-?��/Gw.�E�ȳ-Ax�M�w_lNP���ʚ���r����^Z���g�b�_���|�n�ٸ_��2�E��@V�;9�۟��*�υo������{�JHlzP ���V�E����0�o�Mj�5�a���$�U�f�[�4oVEf�M���@v��=)(�7��ʶ����~�!p�,�'�z��'����v�:4o��BF胘�����O���@32i��@6ĎC8}������������7N�Y��7Օc�`b�1cs&�"]�d��O���c�4�<��]2�Au���vU�����o��?	�(��"��h�M�qRdr�9�mg.NmO�uQ�[�@�Μcyޙ��Ż<#B	aa�����]����Ն���1@}J��u�R��	�B�!��\��Q��Zh��[#�2�]��
j*_�6�Dx�I���
�̬����7*��'�.o/�h���2���4��(�����2�2�8˽�k�8����U��sR�tEX[6���]I:3���W�AP|���)�=g��"��	J�b� ��cl�~��BB7L����mW�3�#�+"Wti��<#K)��ŏ!�U�2Fv� �a3٘)�\];޴ȹ�6���f5��vz/�*G��
Mu��❔D���� ,��+ҐN�E��R?��]�U�*FhF7���:J^9=��ĥ����v�Te��?a�.d�l�cU��ɭ4�%3����d��\�H[�pW��5�[/�C�ܒf�2O��D~�_R���W-K�գկ�S��B_z"�@�Z���p#�d��߱Qu�U�k�T-u��� aC���r�B��J�ש�Q	9zTt W�l��'A~s|iH�����p�ϣʿ.��q��t��g˯�e�e>�^iAa�"U-<D�Q�b�/@���|ikEG&ˎ���5��  ?�Ƅ;�L*Y��7�ʼ)�˷0z��;�$@�� e��0�do�2[���Gܽ��yI�h;��q	j�JJ����:g<����d&�(�j�10�n�'�T)�
�1̥Y$�ה���M�N	����s��77�ɗ`�v,��9a̻tp)�!KV�ar'�d�AU�ꅀ4�� U����:zd/��1L���i�@�W������(m��%�$���H^q��/�����[;�N����l&�*��^N)HܕY��ҊWC�p��6U����"[Ih�F�������d0�'�9d�f7�2�B��Ϛt�Z�w�D�M�X�em��s�Y1���>���4�k���4��0+�8�l��â���(v���Obr�G��v9���z��7��QAc�u3-��|H'p���p���m]B�뎋��do�\ 1���f�.��v��j&"��R�M�I�
��������$���Ǩz����U�Z߲�V8�4XEj����sJ����M�{:*_xB�9��L��g$Eg	R��;2IGL3��5[h��MP+��6�^e���ZVo|���Kd6/\]� ZW�au�[X��ߐ�S�9����P��p�z�ߨ���s>aIcJ��1jfg*��Z���l�\C7m�(���\)s޿5=����ʚ��J����g�^e	���S����W!+���><�}L�@�ζ�y�ӆ�.&���K��w9���ģ���B��`*P��J�&Q���;$3e��﷼�N_\���������sNGbխ0m��Y!��n�6� �b*n(j��X��1�a���s/�Ŵ`���(��E\�I�����q��H��-s����<��*qуk�ӛWPW�)�q7k2���ً�%��Q����|��'�:l�G��!�c� *"��2��%����Z�f}���ߘ	�@i���L���|����ͅ(��Sj�$���������
/:��᭝?vaDآ�\����+���+��Ec�mq�=�7�]�!��7�FC]�|�ұ+@:{t���� G*�#*�5�qCrUV� I��
�{�1!	�8;��+ه|%C2j��u��o��+˽ǐ��#(��^����"�.�|,"�?���Sl�h���n��e���X�P���m�j4T��� ^͜a42�N\�'w̒�ӔO�����2x����V�g�s��b����Gku��&���n���`��a]��i�l�[�6�?���΢`�m�[�C��]b�MńW�g�)�?
�'��;�7 �t1���		Z��m��%��wfa��T[A�j�Ʊ�������4�"���H�m���RW��������L��jͮ^n�X�<��/���B����V��I���[�W�*"����-��*�f�l��<�"�VE0�2迁~%�h�ҟ+�UH&�����I�^U��F���=Pgb����7�+֨����[�{��w�����O�К�Ew�ҌzAz���dm�@,�ݗA�h�!mm|0BY�c��Y{���L�4���Qς���Gi��ͤ���۶�� Pƍ:ׅ�܍�:��r��x���hq(�#Ѫv������>H��:G�&WA:�r��ŗ���b	岢��ǵ3��l���OR��O뚿�./���A��仛v(Q�� ��`��T̀$!M��Hu�j/$E�@^@�/�&)��v��Q4ǟ�Fo)A�@�wm�:��+[���Ip��L�]+����-Pa��3w���7l�z�������%�߀���������
Vp�H�� �U���9����Q���4:[�
�_�z�	���F��Vr�.�4'
�p��F���d���[�^������F/�1V���V�(�28�vn���`q���P��6=�-&0��)d�Y�-C&��r+Ny���c�	a;J����>�C`��.��B�������c�T�ڌ�O��	�ioFtQYg��}�c]����b���MD�D_��ODv�J`*��Hf�b���*�_�v�����H�s~�ݥc�F�q�Y��m>��*�7�2>b/����&N���B[:^���b�C�7ޔ	J'���$h���/���w�$����e��?<�=.��c�Y�)6���UZ�Wo���J��[��[J����ݸ��v���� l~��«�[$Ə�nxe�+�Ω�B ʞV�֛߷*g�=�%)7��w.�}��HO�s1g�-���}oө�-�	�a�"G�=蓊V���́�=����r�TFU��)4���l��4Җ�Z������X����o2Apr�z�Gl��=��@��Q��G�%,�3ڽ�._�ƞ��/G�1h0[)'��(շ	mt|�n�lO���v_�d�H�2��{��🰐�]=�#�5�v��+��l{���:��_<!�{�?�p���:y�`��[�Vy�K/~��yn*N�_x�������f�{U��3E��ē{�I��!��!��
B.�@jT���	o;��]��e��;;���yeYl��/��f �y����嶡	Y���ܓ�����yN��f�hp,]���K`p�	xIz�Wh��չI��$c������T��Nm,�a-{΅�R'\Y�dT3Z���� v�"�����L�S�����p�W�X�F�hx�@w�n��ͩᤲ
�KK������~(����q���3�q�-$u�ׇ,������%�-��D��]��,,B\�`N7A<!�0���	���+�~�rk��>vS���8+X�8ĥ��߫3�&W(��×�6 �̌����<C���	h�K��ƻY���1���͢�1�i@F�f��t���b/v
��,@.�c>��2����j$ε�$ѩS�[yg�~���l�����<�p�?�k�褃s�b�>��5Ђ�	�?���K�������(���f
� u	�ac�yYq'
�����Dn.V�P����w�KO�L��� \ �kЪ=k�=S��fC(;E�!�v���ݸSlm�A?�-�tY��۸�ω��**8P�B}`���^D>v�E�|*�2�e������/�Ũ��Ao�.,�x��0�x��L���XF}�D�YU��P#�U>����x��z�%�ۂ#VŞ�{�h툫ʫq�O���J���1�#���Z-\�ާ �l��t#2�����l<F�Ls�eRJ=���p퇷�繜HxXF,C9ε<�%jbT���:��^�39�*ˡz-�B�[;<�u���+�f��iPX�9p�9_�=�����@�
�"��m�=l%�#��.H�)���;@ ��$����`I�}�B�r�� ��aݘg��&�������O~ȸIT%)9�wr�S��=v
Y��c��GVC�ώ�f�^ix�$w[N�W'C>�g�`w��=��ȍ.�-N<�x��W���D � ���6���M,�~�rz�m�2�{!@�`��C��֍ɶ��P��)ݜՐ��k�,Wyi�th��{G�D�9H_�P��a~��pQHh+:?8�)���ܤ�[`+Fr�DN�z^G`<��K}�&��2�UA"��ȉ�"�e����o�bc@A��9�~r�e0�(0NZ6�骗���"(*�j!yI=���N�hFg��	����u7��2�Ǭ��>4���ƛS3|����k�4ر�J�A	���U^4�UY�~�B���Qϡ3���<xq�L����"�b9�u$*Ą�7��J�|�^^��>��bf]\'��>'�y�D�cm�U��$,��a�[�;Re[�j���d1;Gkx�2�AD����^Z�|� U_�/�c`u���m�6!�YI�Cyg;��: �4�w�(T���ɜ>}d>^N'�Rd���G�锚��Rh�v�'N��^q>z=�d�;_���,���D�+5�i�إV����;0�s����3�Kpz�|��!IT�iGh�	��f�[=����_����얮|��{d&XǶ����u�:��w�l͚���.��G���#��Z�B��7�|�Y gI_u�i�/���y@��� 쫔���Z\�;�uw���r�[#N��{:.�N�ooY%0Q�z(ݔA(Ar��������n� ����Oc*'Fpn E/
3�4�;T"�Wɿݭ�"J~�q��4^'�
���w�
�iD�����Z��@�X������#�)O/�����(8����Մ��#��<�F���
����)���%�ū��K!������v�jޥ\)�`�?�Y?�ƥ
sN ��Be�"��������+в/l�6ʈ`j�����x��}"�oKmdpzO-��ٴ5h�>�{I�����Z{{��w���l���בl�qt.��cqM̘���Fe�a���W��^�3'����������Jn'Y��U���9��<�;�H�A������^��U��.�6��\�@NV��_6��mb���y�k^�����S'�Lʐ�����yaZ��5��W��ڹʗuzܑW��{ʨzKKm�z[I4tU�q1���4+�\�@C)?���(0���An�����u�W;�]�Vu���� ������c��Zl7��@�c'^�	9z�!J�kB
W��WOU����zML$��"���z����RΣ�4�j�j��C-����1�&��U�>���H��]U��H��#��vW*$�7�`��{��$�bۂ��1��ԥ+OlEx�&󡁘z�b����]<zp�o�?_J��v�ly&r���~�3a����h����6 �%{�lH�SDD��e�D�X�6p����H��Ȗ�3�ӕ8^K�$u�q�����6b�Fp��\�����s�~�(��{��C�''(_��uɡo�:�P9��yU��%�綛y�:��rV{y�)�}��5?py?��.��WiE�C��z�[�յ#hʼ=����DIM-���e�}�΄gx�`\�,CwgZX�.������=�a���'�Cn�U�b�AKu�9,�Dh��g����ʨ��uU���\�m}���Z��ͳ�RsySd��x3&��>��u ��
��'=��l#�%�9��j���
?z�lmK��� �fB���kڅ��pR�@�ڷ��,۩���ıx#c��Sb�O��'>�6�\�]g���cna�����̀��L�#}����`lY��k�0�1�E�	R�뼅y�]��&
�J���
�]Ρ����W(��p���2���QLշ=�$�7�sG�4��4O�f��9��3E��Ј+๙`�}�x#?���m�C��oc/A��Z� ��������Z&| ��ϭ=��	�N������x�⿦��% V� {j���Y��lpz�SET8�ao�ݻ��1)�<(������M����N:E��u�<'�����Q�-�����m�:�̎F4�BBψ;I�*�ϟ2G��t	B�Z�x��`���~#���<����@R娹H=Щ��X[����G�����X?vJ!���C>�|J'^:ϱ{��M"�P�$�-�ҔW2��8#�-�����l�� n(�!��wP���� �,;kљ}uX��ɢ4P��%n`ΦG�A̔� y
��(&�6�7�a�o�
�U��!	*D2K )��N��#n5Q1��m{@!���"o��e:+eG�>Z�씯��7��v#���c0����\�H7���
λ���>w����\�
1^�:��bjuN�hng��Q�G|����n�(��n"E����gz�C�85���*�Z*�'���|�YU:�� +���=.��ԕ�*\���/>�?&�ȵ������������+��3��K&O+�{��,Jl,W�ڣLT������i�2���$$TN`� �H������t���7o�
�@kX��g���Y�#\�L�.8w�<��;���B( nŧ^�c��bT�D�;C ����:��S@o�g/!�ְTw5hbE<�C���D�r$8�L�SAp�[�!�h��G}�	��E����*��|��\`p>�&F�X1�_�~��H���9�r؅���TF�ٵw��5����7S$����\�/��:�ׅ[��.�[7 ײ�����	���C�ü���r��Jm�s�^p�GoO}� mlC7���=��
�'r.Po5*5�y�%N]���H��ca]&|�ga�gM®� y��q|�<���aa�S��*��)���!�+�l�i����3��hU!�R�`n-�v�|��켆��n�d�mD5�S�!R0k�D� �n,QB�0̿I3|��魯��(vH�h�ޔ����J�ҭA/��G�)�@{�5�Zv�JEn"t����:�5SŃ�������_����9jSi0�XE�$"��<��W�o�Zf��ض�f ���Kk�ˏ��I9.|��r�$�)�l�o��P|N{���	5L(�35�i����Z�����9sA�L;Z�,>�d6�$zG'gOϬQ0�4���i��lQh�����sWt�-bh7�r����XD�Lb��o�v�!h�DLG9����`.�4��t���P��1c�(;\�ĞCT�H՘v=1bl������ 9��ݥ�+�z'��:`��za�/۪&���=|�AI�U�o��<J.����4���Q�T�u��-��E�>x��\鲣=[��"��{�W�mM�c�G9�(�� �w� �
S��D�q*���i�(��(AU3 ����<�`{�wͅ��c��nE�8X�,�|+���������Y�-�ud.�t��!`��w�a���OQ�̔O٧�*/�(���.�g���l�
�]�2�P�� yn�o��SV�e�_�N����(
���y�T�e!�S-v�Wt�߄��s�z��)��$�;ԏ\G�� Dj0S`�l+��3F���.] Ӻ�h������l�Uҽׅ
nO��v&h�3�
vo��1�f@ �y
�+�qX�;�oF����d?Մ�<����;+epE�P⇆���-"Lי����mB��D�_f����R�s"]��4�n����U~EF���b��.�@�|ˊ�Wy�l�����a�] z���Eh+�W�#��Ҥ,�]�|���^m�U��	9�+ �J�9�o�tJ��;��jS�\B�[ߋ�>sZ>4�6.� �K��_��W-&���(�/Թ�|?�k�����}i�i���]oԐ�4�bݫ��K!�6��__�S�ȯr���0����3������T�B��p ��4ɍw�53�2��g��_4T�:%��p����@Q��sc�ਫ਼�"v���yZѺ��GN��wn�_s�E�W#l���<��t��OcJ��Yh����G�#������T"�g���$����S�x�e��8��=[���BSWx�_앷��P��W-��lII�WFÙ7�h[����*���a~�����;�A�m�1n[癓�����C��=\]��w� &�k�A���5�˩u�Z�l���n�$~�k�5[�"&�}����b5�"W�*'><�1��0p��r���Щ<�!��H�裷Q�S�}�aoS�0���墉k�.��z43�]OHC�Om`lQM���2��'K�b�j`l Q-�W-:�����=9�0���D).�K��5�"b�����p�l�T�H���A�I��ԺbF�N�Lcr/�,,����-F��M�H.��x$��#�d�44���o�	��?�w�ŀ��Q6F0b�`v�z�Fz�5IN�o�d��Wx���Er��S������B<+J:���+��qs��<��mA�������&gZ��� �'��!�-y���ۀ��1��2�~��l��JH��s��[������˛����؜NT���=~g��-���`]=G8��bH�,� l2���$��28��0^3���(��h7�H��e�|��&"��a�$�V�∡"�p�G�p��L�V�Rc�S��[BU ���sb�bf�-�c���s�x�u::oe��ծ��h!$E#Ha`?%,m��Aُ^� 岂׾��$�z������wKV����P���F�׷���'��$��e((��Z� ��P�hs���B�|��A�c:��[�T��K����ۋ�6��JW��˝��6�Ӓ�r�͹�֟yJB��90��� �'�R.�������側?�Fn�j��O���� A�4�G�_l\�+b�G�CN%"LXDD���*���`K��W�'N �<��$"���f��)bG���]�����JG���oc�����P���ͻf�/"@�}Mч8�C��n�{�!"/"LG9ϋ��;�,�w"��{Z�e�UW����X2F]Vc�\�����>���������y���@U��(3x.���V��<�����Qy��E��#���_سj��p���r����������\ƪ�h����Un~=eb�7a�ĐZd&	�uw�(�1�X��:>�l�ânh9�!�t�1'���(��\�17�3k�/� �a'Z���It��Q�]�`,83�C� �Sk��mt�s� j������.��{�9o����d��Hk�s��X�&��2=��YGq��b5�o5����q��~�oϥV v�Z��k���]���g��(r���lݓ!}D��m���J.ܰ�X {LǮ �m+<��)S�!�Kv����w���_wYb�V:�׳t��Z�U�����{C��̬X��.�<v�+k.���i�m�3pH��>��9����B����N�8���v|���c�1�_��W��H��hN<O�,�#N�G?ǈ4��i�;���~�����2kϰq���9�}D&@_���*���[Hȃ�2z��V�6�sX|�3U#TKWџa77����l�bMc���|�����ʤrCh�Ҳb��	0c�>�
�I,��W�3#�L���&]Eǡ֥�t���r�P��	�M���*�t�g��q��))#F�O����P�5Z���{)���T|o2XKh�8u]=��|�-��>0�zK�#e͡m�0�x'��������ȋT����9���p�;JQ�=������x��I�s!�x��c$����r�ZqY(��'��b�����N�I���/�9v���j��_���?m0s>�����\��E���} �����Ǩ��������X�d�Q��Ft�U
���G>푘orFYCx���3�T�v��g泑�h���Z�����-��G�MW�D�����%_���B���vy�ρ�g�`ii<I��.�1��¸A=���-ѦhjW������2G�ͨ*j�P��5����x���6��A��m�ʬ�"A;`��;��_Y/}��qµd',��LƱC��p�qm��O;��/��wuV�P�!������]�Wm_I�\;�f�!fIW�'�q��O��S<_��Hk>�0����7�^��쥀K�uP�
ʎ�����,�	�i��)�
)/9X���J�8�b�upD���Fi75# ��[�f���l�ɵK�A`�6����@Z�ӫ뎤�wbG]	"��jVW<��b3M]�Α|���z����t> C�� �� ������;a��3u6E�u~=��}�]r_���dMDm��r9n����S?����n�S{���Ҙ�6 �w:܁yp����܆�x(/��k�c�Fo'�X��,�S���lR��l�e�5Z`Χ��?Ab �M�u5ׇ�Nz��؝NS^||��b����➥b/�8J��c��-��f�f�R��Е �%���M�P��&�����~��S��ሚF�q�&n�j&�!XAE��(���!���&��Ȃ�Bq���B#۱�|)��?h�]���*5x���p�讅7��9�U�o<����>�$���l+�M=h���k��ż�O�̗-Ц�D$��+�<����RD=�9���+:��ТI��2O����l%@����z�<��D�cu���JV�ɥMA觝.��|?����{�bT���-��D��,�^�F�e�udZ��n������[�"�G����4*8��r3�h��9�#�z�.-b��ȩÜ�V��3���)�������ԩ���މ�����G���;v�K��wove/L7>~�rv��;�9xu��%�a$�d�y,]%�<����7N�S�!���rw�_�%=T��a-hB�%j��Z-Y��gF8]�XB^�^�v��z
<<�-:�a�?'�Ŗ��\��t��[*n�L���O@�}q�G�f9}�^|������IΛ���x�	������3�^Z�4P}1u���C���*t�\��Y�Ȉ���ܭ��9���=�)������qA�D��u�27�6��s�}OiU@ID��_�:�׌j�/�&�%����t�Wc�x鎽��hRw1t>�-f9��e:�
y�#ii)��.�3�1&��e���%��T�����R4m�=���.��t��m|������4 j��͢������bb���mKڹ!BB�'}�qJ��κ�r�.����ry����:��T4 y_��sW�6��wпp��{d�C_�����NHj��I�k[�B�툛GV�V�h���Hr�ǳ(�Ek�:X�A�D8Jބ����	}t*M�iȹw���)�+v�:(&WI�ʘ�� �H�pT�R�D6�V�c�7%��+�8��	~_�þ�ʕ.���!�\��70���!�ⷶ�J���	9V}(5[_�Qe�}��(�n��4d'{����o�|�CuΔ<v�a3ISEP�F�TQ*V뽳��7'��XeF߬����d_���ء��4!�)G�^��V�LT��e��3=Y�MA�ۭ���h��O<�i<rX��I�wY|����=�i ;�	���f,fb�&���ҡ��z�#��
hypN�:��TO��1��qE�?�q�:���ԑ�3A�a?��O%��<�����a�x�	^&����Bh@0���ދ��ie��ν<��ܽ�ٞ8��@�'n�B��UP5��2V79���i?r�#J{K��/1��g�n���{��O���O�����ϫSs$����3�k龦r���,T`�24�D�Ik`<neMF��Y�8
kU�h��'�oh��鰟^;/�N�X��aN�	g�x�ɻ��������Ft���Ƣ��Pa,�Ao�΢����~4���n�p�4��FRy�4v�l��R���TSur�REª��г�v,߭�?E�GLuFK:W.��2w#��"M��br�?����j���`�cP�����3
v�]	���5N����/���_�JJט|�{����E�����9�1���^����v���"�W��w��hu��[�'l���r���0�� ��PΥ�Z������\3���zG�
���%#'*wީs��uK{?OsA��ҝ�b:A�OH�ƞ�>Fg�=��K���Qx��5��s��B�����!($��8k�xX[5��D�jK��36���%6eU:)kP��ʦcbOzO�:o����v����䤤��5��#�'��k��U�?��>1+��A_>��(��8F�	�g�I<D������.Fřϗd���[q��(��^��J\Cw�f=Ҡ���8tA�3�A�=��a����d3d���a��L`�g���C�\!L:���
�|#B��]B�����eHz���9}
���n��&��~ۀwA��:̳�-h=�R~0K�����v��LiM�R�?05M�����:x���Y�u��'��V4���a�����KL��.��ݯ�u�N>�&F9 8٦�㗠Ȅ�F����Ч`��ƌ������:���.���.�z��Mz*�}4�FMq��B �c#8�=̀�������w�q\p ���\��T�h��ٹ�X�d� �u�𺋗'��.�����);[��EDZd���>���p�LsNIo��us!f��,T�Ɠox�o������L�=�@SN#���9ȷW㣨o����)% 9Y	��\�Z:r��'v�E��q�J.}���������wo�#]?H�G�1�J��v�PP?W״{�S���EP2^����gcC�I���γvc�AMTb�D48��B���M4<X���ؘ����hS�8�L���Pg4�j\�~b�'��KW�.E.��o�*��ʫ�s:vؘ� ��5f�o��
�Gk���[�e�Ҹo�4����>�͗+�~��&�2�GP��n\ L���ҝ4W~��d/HQ�m�L�<����>������[WR5q�a��)�OJ�%�z��o��Y�=;���N�~F3�K����v��-љ8 ����:�K��9�3�"w��R�z�g��{E��Z�M(K34��5����*�깕��W�*�\��j	+�1t7���΀�~љ��5�Iߠ�z�I(Ls%�ލ��(0�nҕ���
D�]-@V�M(��\54�=QS&��jB�XU�����.X�o����_nQ�i�ud^�J6��ɾY¤8I��$�tv_8"�U���A=����rҞ����˙ ��a��"3�1��\V��C�xyŌ�J~$���*-�у)`�M�U�2�*�D���@0T-�z���nQY�>��DS�ȏ���\���ԫa����?�b�_]s��~��j!t����moF�������������-.H�Ē{��$�7=̐b�� \����x��x�K}���֪Y�^ns���'w�kZ}-�7��CL[3R�ȳ�վ�[H٫�"�X�Qǧ&NW�[^��h�j�>L�5�VJ��恚��ޥ( 0�"�Q�Tc�$q��J]GD�/�e=|���u�*��mܰ��9>_�1j�0�1���׺F���ia�� ٨��M`@*���� �d�q�q֬s|��14�7_����[��܏�(>ౝ�q��E#�᳐��f՘���p�u���6���� �+j��M�0q��y(]��g��~�7�B� �v�M삻N:���F�O;m'#�����RA�m�R�p�f"*����}B�ڜEʥ?�ceYs�ֈw*=���.�4is,a^M��Q�r;���o{FFF��ܩ�\���\���w2��1���� ��ۯ��X�޼�!\��{6J�$�Ϸ�`���bRVZ,q��Ŋ�e��T���ŉ��4\���5����V�����q��\i�����ܒ���aㇷ���/���߉Q������ּ�.E�r��~*���%�� �<� ��������K��&��j۬�F��i�Ԡ��F��c�=A��(���E($�݀ �)L���(����L�E��F���Kd�#� TN�e$�#Ӷ��vtФ&21�O��`H�1�br�1%7�)��s���)��O�{ф�W銈[ǩw���>�^׉��ؔ�Ҋz�U���#L�R�pgzk�Bݛ����#����MB�ϓ�	7lof�F��q^�X�����נ0}����+��%=��0+���	o�\Z�Y��/��6*㊎g$!~� v�#P���&�Y#����,�ڏ�$��C�{f[G
@��c����R��:M��Σ����٧.��8?Z�c)>5��4׮�0E���xY��s[*���yeZlt�^ڜ��٣�	0��Bٍ+����i��hZ��*ƮP�0\�x�Ql.��.��X��������qKXT.�\�U�:K3K�SCZ|x�8�N��(�����=m�*��>����bpZ|5����%S�LH�GC[��7�>�8h�p��Tbt��3sN�mZ{��?%X��υ��xA6���s<BH�A��m����f�	�>aǇ�!�3V�D5ד�L�>f˅^v�k^�'n����tr��\"5�5�f��ji��v��]ظoW,��ɥ��[MC�z��4&�Y�<�����%\��ۿǾ�[ԗ}��T�ZX��!b�������ѻ`�EUB��I@��a���up���$��e������4H�g
i�y��f���r�6l��Q�m�9ߴ� ��j�����]»���ur^�r[��G��XGؑ�1�� WkO(��L�VH�]w���;�R��zt����'SD���,kC���D�	7��f�e�a~��ؽ��-l���}n����V��wq��A�i&��p>T�g�T)o�Ý��%��ǻp�M9��
#4�Y��c0~W�I�dV���7>?�S���/^4�����6�b.��x*p���S��%�r��=�"GdT�ןQ���>eO�zP�U!�NrW�۷6��؛4�3~w��f4P�j����`ϼ8C|��K9�g��P-������Pc߱5�)C��?�]	�h�x���z"�����.c���04	NU`�����pl��y���S�%+�"ͮ�M�(9�Zt_Z�m�ӯ�
ғ����L����C���G=��0uK���g*�SJO���<�q����P��9|���!��.j0P��>	�8�_'HGjo�������5�B��*S��iп5�9��7���1�4��E�y(ޠ�N���\�it�	N t��H��1��!��l�1��ɽs \����+���|OFK)Fֳ��<h�QwBs�=
ߖ�<�y{��M3� o䕲[1ûp�oAc�h�J���7`x��Y|.F'ٌ$:OA>�f��3K|��8���������w/@��͘�5!Uc����#(��t)��@�}����Mr�[��m�u�ݎ&rFU�4xP�L
$⻓+�^6n��C��� ڙ�Q�����)�>4/�@����N���M)C�b�г`+��+$���BD����s	_(��y0;�6���tc�\��- h1���gQ�}Ħ`-V	��/������7���W���Q��8�t���
�T3�^�ѥgH:hW�-5�o��
�&�@��Mz������G��'�-����]����?����&�`!�}=�7������YB)��3be�ɉi�������	���r~��M���Pm���w�GV�g�|�#h�#ȣR��������7���&�S��"��1*����)σrs"��_QYڙḍ���s�kL[�Hw��Md \�T^�A/���],xnU�^�i �X�h8o|��
Zl���s���梒�C��
)2'�;ա��3$��t�����Cc�~�LT�T	�2uq/v����AsSJq��j����m|b�9���]@�m*_��n�l�`���	���V�������o��ep���J����� >)Sx��φ�&��h M����WqJڢ��a�C2��J�|#!<A]'��:�
=�L^��.�-��v]��V�/!P��[a4�FͣyK�����3�'a���(�N6���H�Y�!,��2ȄGZ�&���o������;5x�l�k?��Z�d~�p��2*+*$8RU߼��bnx�� �ڌbq���U�*]��BL�a8hk��oÁ�1��oHސnl�E���j�i	ܐ_ˣ0���块QO-��Zj�`�% �wI��o�?XIh"!Xvr�_!H|ؤh��&O����x�.#O/1�j��D����@�;D���N}�v��\Y@��%W{�����Zz2��>�TB�i���EY[����Y��_!�.nq�2i� �=�G_�(u'�u�)$�	#���%կ���,���
#c&I��d�zh,�Z����չ�b:��"���
Bop`N���K�0��K�Gc��r��Oe��-q�dq]����'���W�n�S����_�l�D���N<�rz��:e���	�0{k[�K��u0�[�{8��b��ۦYYe�7���]��$6�$�+zu���$�h�H��w������ �i�?KQT)���ؤ���i��N�$�nY,l���c����{�=���\�`�T߰�"�D#S؜�v��^�*qS�bi�F7�[Gm�	�㬹����==����M��2�\��qzK]���!B�%j1(�M��b$���R黑���D�辘�3/;�-�s��RT؈E���/d�D���'!�c�:��qSZN^������W����Das��{ci]!i�9A��εw[rz����C��fP��J�M�M~S/��Z��G��_������\����~�eH���L��2Ë�xn����bZ���k@�"\S����/���"����h"��o�8�|��4��`�{9�$-&PC�}.����mn�}���e���Q�<�I����߅��U6o������e��K�zJKC�	�(�堕wݽ�Z�v
_x@�Oⱙ�!"O�
��d(�S��Z���Nؿh{v�f��b _:%�0(�nJ�Z�?A>z¥�*=��ol��i��<״���2>�Yړ���Е/��۴�`�"`ke�}QB���D^<g�.�M��NuIʃ�Z�kך�~��ygw�L��3e�a~^|�&"1=뿩���.3��PA�p�2��!�,��-<_�0B��1�N��ɋbJ��S�tL%K�>5˖XK��A����c�'ɔ��PA�+��<$$en�S���s��R6,?.U�.��,5b5�:DgƱȾ���	8��������kCݢ���M�a���͇�/�KhK�^Qnr;�75�?@�C{|���G�<<��-y��o���-���Dgi��T"�V�7�n�m2K�~���~�ܙ4��!cP�_ܠ>DH��JsӡMT��w�|��J������=���-��h����<GKZЏ�^�$�������C�6q�q��-�ʽnK_���t��Z�z�V���:�K#:"��Þn��lǟp����"��A1hG%;O7a����%.��舱�H��x�c=5K䑧)�b�@��
��`����(�<m��lrN*���� �k�H�|e}�����YceY�9*C-P�CŵG2S��oX��H�X�R�\�V3����2H�H�Z���s��G��<�gY�?Y�,�o}��oL��t��(��g ܄Ů�r]�[�x�V�;b���lU�)Z�[ V�Hhd�z�$� �P�)B���'L���&%���gr �U?I�f'�G�O�F��A��t����$O�,r��ef��a9���=D��Bet�m����1�1�&N��}���;���Wa[=ƚw��F�32�.&�-��ڑ�EG��G�?z�8Ny]_ѹ�0�Q��eX�:AӜ�,��G��˸��d�Uòr-��\n��$�&@�Ź��Y��O�'�V�\������t8hB�k��P�4ǲ�� ��S��{ʘ��.Fȴ�k{AN��A�LK��w}����
K}Ѭ"q�i����4B�>ly͖Dm��'T�'�ETt5���[���?���S4�S�*�tla�s��;�H���%�r���ӳm|M[���������E��{��r:�`6��888
N%m�b�ޓ��~6�n< ճ�[��]�`{�%�3��9C��~���G��R�g��,'���r"*�H��߷�u���0 �O��Bԣv�٫������K�F�c\��m�	ݩ��xl�^�l���K��2����rF�ߔxj���Pn�	�����o��2Y |�-ʀe��n4yYhs�*��r�0��S�%�B�nN�����/)��
x�6�����������B���%7�Λ���\��X�#�"Ү���A���#�����7��^j+N���3���&�)�EV�g��d�tz튱o��d��g;������09�Z[�ᔔ�,_q���̓=*����R���Y5���p���5�͊_���r�a���-��y����U<��7��[�h�Vѵ+k���T�����;JS¦hk~��)D��Ȅ2W��@�y�zA;�v�%�|�k:���H����vk�Uֶfo�v���~8d�Nkdz+�2����.ro:m���d���f>����Qӎ�-��n�Ѷ�����]��-������Y�Ν�˅n3�=��4I	�V2�jI��9fٺ���  �b$j:2bi0��N:���[�w�W��f(tU��g�5�mƌ9 �PW�r��H{�I�P��������#]�����,��Z$k����z]�ZM��yz���=z=�x%y[�7)�]ɖ��� A�@E��Bg��}L.,p�����&$�� �Kw�y=����%�����I'�J�F��7r��?I�Z*.���8��֛���Bƃ�%���Pre�8�CĠ�Q�q��y`�#ק������o�V�<�&��������+ԃ9��pF�A���EB"�$hZ݋#V��= �A���9҉�<�AN��
�C����)�K"�n�Y�d%0�B�a�m�,���w*�N�(p)�%dϤL���|8��؊��^�n?�g�FI%�$��-�τò'N�������L��8�ZB�+l�g�w��Ҍ7;�
E�oۯ�LS��������d��o���R`EB���HV��f��f4��� iA��ڭ�6���!����'�v~�O1��R�E�1�(�W����p�g?n���5�R�Ǚ��U�+o�*�ݻ��k=%� �u�b��ə�I�~���e���Ւ�\k�?�V�$�0;��lmR.;�F��I�8X�$���@�;_$����R)31M'�5�/�w��'���^8�����>�c���!�˫�yN�H����\08;�Ʃ�J>�Rd69�%��,9�2�W4c���~������b	E�0%!�x3��4;��	�r�z�\� ��m~�L�������B�0?]�=�|�!�O��Y���F��3@��8���;�����J|A}�e�G�Qx�ߨ�P�z��a`"�{tC$��
��-.��2[r��%�ȡ`hK�.�:�l��l�>�_f��fA������^��'@��;��$8�x매��|«�����1b�R��\Ohii$^pv��a&6�l[��$�n]�ݚ������t�x�&��)%��.�y-q7~�3�|ґ�þ.w�Hj��@Q���;7�N��-c�����?������#�x)�S����\���P�B�d���<��~�m��"�yڭ-Z,��󤓏�����&~!�u����=q1��Qu9�<K��)����������<��{u9 ��w77�ܵ�b6��ջ 8���Hg��i����^��z�g�f>�+������L�i�K����׸�#��h!�5�ɘh�B��ɩ��M ���kJr����u��(�ùʑ�>�(@~�ȵϪG�eWޣim?����o�z�����V���s�m�jQu�>&a�Q<�3�U�F�FJH��^*�-b,���N�I��P!�Zs�*<�G���$�p�&2i@�lI������М��F�zK��P�(n?fRɤ�m�)�9�e�e�@H�'�����_%�t��-c[��.�&�b��RI��9���mP	��iN�ӼJ���5��5��CQ�c���d�D�>^���.	E
�ֵ� P��Ro�w�v9�����E���dخ'�9�o��N]�%#�������~H�vsYƏ
i�SC�����6�lN��N��*#}�S`8�'.�=+Ugk�;�n��*o�KC�Aoj�,8F���H�Q|��1�ě�x���ҫ����v�	����f����Xs��ֳͿ���a�KdLt��=�H��ڰB>�,�O;��%�N�+�!�H	�����ޔe���������z�|`$l�x]S����-b r&���t�Ntw�@yM)�X�5�X�C)1�=]CP��u�[o�[A����(H�$q��Db��_m9�2J'a�mm������������]<D���n��.d�dgvݎ&�3��mO/5q���rFc�6�=ne&���|J��ɚ���rܨ�~d����;�ߜ��1a���}]��7U1FԝR�V�FM^q�RP�p@���2�y{oHd%�T�b�*&ZK��(�P_��
�w��N)jk�s8���$B���2<B=<Q����]瓱�n�W�!���$���*���m�"p��SO;t��� ��^�u&���4{��#5��ߧ�D�M�+�����`��0��t�w��9�q�ȶ��0�����iqZ�����)���D�Mw���!�g��Oa8{	Y^	��V?���9���Yvg+.b�|-��� �p&�Ѐ3K��S�8��M%�`��F�P�d�x�=��}Ky϶�0\�H��[KXx�=�;,V��	����m�d���L|��"�t�1�� <tt�E�+t�7�X�֔�����Uw�tP���]ے�tvߠ�#�����JG��F3��9�&�C�Y.ZWgh;̑�z�#�U4��a���2��*��x�e
ť(��M�T'텘���J�a�/4і#V�&yv�^r[ķyV�3an���s濸+w��?�0v��hj�I�xL͉.��G�����P)�_��aAl�׹?�64��J�Wͺ�Q0����w�?]a�L��9�J����ϏX�ٲ���UD�c���������|33���}sT�UZ�3�\�
�q���D&����7O �3~?��!Y�9���a$I����c�a&\/�=J�!}Z����P�Ú�kU�X��|�w��z�� �2)8֡^���Ns��������P,�`�*%��$R�]P���)@�� ��Hiw[}!r�
]^���T���2���3딤�N�d],��P��İoucMbϤT�:
�)��%<[��rx`��3�J��>���6ڐ:h\���y�&�YJ-Kw)�����!C�X��)|x1��~�7�Y4@���r.�*��6��ڂ��g6�o��3K�\�A��5�nv��ش)sG����w��Z`���WaX
���%z���[�[n�j7Q�y�����޵�K�Pa��Ո.=�3�-}���y�����Y�W@[7*��B3�Ъ�8�H͕˳�P�Ad���t1=J���

����"���,���h��T�pf����/,��:��FcߨȘ�9�;��;;���+�uxF�%��xzJ:y�w��MY`�l��/����K�R��.���u�*�/mEA����2%�B;����U��;\v:D�~���{�	h�����HK$+�}h���C�"��q�Ò�h�:9�&ϊ7�&���6��'M Y��unJS��7LO6G�e���,a��'�=f��\
B�) Mp|�=����	����?��=�L4Ԣ�qp��vE�������&�����m+���T���`�B��1�ne��y����#��Y21d@_Ӑ���x�Y�t���o����?� �
�����OFK�+���[��� ��:,�j����3�e�� x�5���V���<�G|�&:����p7�v*%r��7]^5a�q�i!����2�#���GS/�gpN� =@�H{�6!k���3��o���l�v'[��0�~���Q�Ѓc+�/R�]��F��9����^nA�׸�&�j}��}�)��!���cUK.|M�2�ͩh#eY���_��F���x�T-�5F�7M��}��?�}�Q����<�w5��7�o�o�$ݍs��+az����@ft+�OE��z�����z���JH�$L��s�~����0�_���Կ�SW��>�:��e�oj���B���6�Y�X��֗��$�d��Ƈ�u��C�e�T#�nD�cƤ�t�Yv���
�=-�s\�l�`�D��>#�*o�)�x��L��Qo*4K�\�衧��^���A�u4�=�� ��{[
�_�����y��{[Kz�L��n��>�\�R��TK*A	Mw*�����Ii��;%w<�l�$Z��"���2`�>@Q��gP�,��/������@d�c]���DK���*w!��z�_�phl�ܷ</��2�@��5n�B{�Z�Y0�=Ў!��@�y��0����?{x%�1(�T������"��r�a�:��a_�V��d̡���vL)ч٢/LE�>�OJ����1փgN:n
��>�����[�e���;gn�_rT�7�7zy6��JJ��d{���
���
��=r�h�q��RORl���_/�b��NV̔�<�t�/r�(5��W���.�(�Y�-\��q��+{!�������(�t]r(�L�ٽ���b4x�٦W�GY�4��hȃ���KVT�!D��2ܖ�f�d�x���LQ��N�1Y2.�Վ��Z}�ROM��3���6ȯ�Ӡ}�2�.�z�!�3�Țm�k��O��|r�o�sֈ�3�v��[6f6l&<S�� f�4���q�-�pA��QO������M]S����R1z39~��?
��V�\�<=��}=��URY�m�^xlQ��ku���5�E�y���M�/�7{����l��a��S\��b���o�Kw�e\~�#v!ދ������U��s���Sd���W~R����z�8 �X�+�	�����jb�ů�J`n����\��YZ�Ҫ@�B@�F�wR
��XV����c�5j<��� ��9�ȼd�� �`�,x��{,��ҿ����!Jxf�",lQ�	��)6Y���zs��?L�����-��9��J <IcҢ�tp`{wyrwǓ�	t��w+��u�-����hu���|��	~�i1����P¥�r��� �y�}�S���-~��Nyg[Y�8�7àN�a��.삭|�w�y��'���!�t5���`�}I���\2^�&�3���Z�� R$jw�+��srp�;���J�j��;��%ɺBf����?>nZ�Ep\�Y����[t�o�p�>���M뮒XG]2H�o��?���ttO�W� ���C-l%-ǑRpaҀ���'Ò� �,�pX�&s	��+�OH�"A�֯a�[ ���"9%���xv0�B�|� �O�Z_�G��=�&���ᶋ��xuk��Q�´6o:)d��j�����������P��3�_~#m��z£���e�Q/2	��L�r�wSX	����%�e�̼�10*�yn�����
���FPecb�,zf�����>�x�h�:!��26j,�TX�f[6�����YTe��+.�wq<�]�_���8�V�Y�V�J`�E���Jc�8[-"g���7��8�4�qI���ܠ�3xol�8ڽ�8Md68��IJ2u0�W�Ғo[��#W���FB#���f{S���⴬��T,�7�� bH,����v����|�ߕw�Ă,|�*���nv�$s��!8�$�TVYb)�T\�&��FHv�z���xH#�'no����v?i{=��me�9+t̜�I�ÎSd��D��U��>\�d62B��m��(�
w>;�F��;�^Ѯ��+Nr R��V��W���������8�7C&W�
�>E�Z>xj��d0�o&-�(Y�W
�M��E;廩��Ax2c���G�z� ��0_�ж�Mh-�7�	|����)�g;a�E�V��{��<b$z�$��oI����T�;�q�u	4��R�3�w�L�UK�X�H��}���|�E}�NH�5cIr	��t*_�;ʴ�y�Z�f��R="�3_�i~)n�*;",EG��b���Q��	Hp�����s_#ֽ�~�gu�
��-}\zD-h�Q񦼚���Y��/�#���D']m6wM؆�[�����P��3�L��E��v_��m����OX��!
�3���sd��7��:�e��v�d���� ���AC(���@�7^<�@ZS-;�a�L�p_�Wh�ڽ^��A�/�UE.�h ��ڕ��h��=�����brd����aR�����[ZH�5�[�+����Aa�����C���[�V�2�7�zK��J�ۤaZ0��O�S�h�R��4�s��OY-b:��dLܘx9�.�0���>S��@k�`i��q�vS�ֵq�b1p	�U�4���(����lΛb�UnV"��M��z��5�`�Dz�)@ =ϯ ���޿��5JCvz�0 �@%E�(�3G��F��B�u�Nva��Lͧ�ޣb��?����/=�ԩ,����܇JOpu�dH#v��]�z��k��K����{u7��J�����;��qv��q_0��.g��D}��I?��ј�dO�i�o��,�m���v���R
�K�P,h�2V$
;��3�N���9Ǐ������%ݳ�&T��ᘱRq���n�g؟���5H���}�t\9B�3�>��C��,~�23��ko!��ͮ�M�&U�I�B�RqLj�UB���8Ƿ}>��)�d��rN�R��T@�I�ٽ�~��(n?�ns��fף���h_��e�6�?�����D��
ɞ���r���Վ�Ɇ�>����K�i������ڞ��P?�1{s�6����ޤ��^�3XYY6�|zx��� qM�'��V����ODD=��[�$�zp[���a��+(f�0���r�O�L��4eh�'fQ`���N!غĞ_bdc��'��F���ܜ�Y�592A���
ee����bh]�n @�����ِ�"��Y�L�i��9���K7��>�4���T}��}�T�M��k� |EU�n�B���$���Ƀm~ӕ���b%|��oڭ���(,vC�����s�Y��+k9��NW�����5=�޷�?2� �v�/e��vyNF]���]x�����W��}�������r�)���b�mϙc ��n�~�� n�+W$��}]@���W}忞=%��'�k?m����Wۊ�ǂ�@!l�\n��u��5d�a�f �����T%�σ��}�;n�7�UH��tI��M{���g*�p�b��[u9k�"��#����<Z!����k&�E���T��*�������f�Fr���OG��V�3.�ɛ|�>���&4�oQ�ٰ��� ��z�|<�3U�},M�h���f7���b��+��?q����Faai揋=S���@�V�fF��!Q?[��k�����{�4����ݝ����|�:+��̞�q �1-�o����&EpU	�p��b��kj��шr�GvR��)����1TBۗ%mFyVКp]���_��@��:�h&#���̟BM���
����&���#���Lj��\
?�2���~���4B�����R�� >X߲޲ݢ��30��C����YP�F$C",q�7�$�LoR�����o!NH��%�̬�H�y�X��Ϡ ִ�눵�����%����if% �5�_Y�W�c�#o��^��D}��{TF\*�������7lZ1D{N��Z�K=��1���D|W����؄ną�T�rP���̈�:OY��ob8�̟Ne}�UZYg��DC�Z�C�`�='C��T�r'�"6ߔ�sd��>���U^��AK��=B�z���5B��3ɾ4���Ϲ.�u%#�n�W�3+Ã�CO�j �u��Vў�Dͤ�H��|S���k;�K��A�kj�T\��{S�<x������ܚ*���UU!�.w��^5`?�J�O���s�L����k:�Ӛ!�k1�6�jg��m܇}����ٮw���X�A�i���>��������x�U�`c�馘v��cH���w,&�ǅ;�7,���%�&��NF�J�%����@��)z�K��uB�z/��A��(S��c��}'^_�~@9qO�Q�L,���T��-cJoU�E��J�Jׅ(�E�{�
"�B+�.\	��<�i��\��yj[~��.��c���˺�D�}��'/@�,r�r9�|��\��s���y�S���T��:��~&D*�h�-_�[�������,�3�sC�����o_��u����O��x���C4����uI�,�¿� �	�qMG|Ȝ�9uਥ�F-L�r�ى*(�	�}q}��n�W�s��r�P��ۘTA{��ړe\}
ML�I1_G�7�r۷J��d~�6Aa�귡�Y��C�6%UL[�o�Vx�_��o2�. �R�>6Xb��6�+�g�Fs��s\3���;��������hL+�{����\��<4���O��W�a\Vh�b��h��}>�GǑ��j`����j�WO�H�}{�t��'/V�yP�@gl��1��	�~N��C��� Ҫ?_B��{p/,����W@�n�T(�>E��  yɃ
�f:�3t��Y�A3��ʣ�Y�<}�o��݇�[�;O���}P��D�����m��[��;tLoc���'� �MA��J�^�J���|�8�oO���l�+�憽?+�!����Ls�Xg����Q�wm��]��M����D�4���b�����a���\��_E������FW3�����VSXt�g����qf2�j�vQ�]IZ��)�T"�����1��
�F��Nv��K���dc����V����cI.�pe�٦9%�_v��6M4���}���\qhal=C�QK}�z���1S
iaY;I`QG��������Ov�+;wG���XgޠQ�� Rx ��M�;�[WZH�^�J���\�|��0���q�Eߢ����8nK�⮳�x�+fG�3@^�K:���a���b,���a;�ލ�4Vl;��3�H��b�RS���Y�= �'|�_B��6Ԟ��p�����ާ�̣��UO�:<2�2�^.�f�o/��w䀖�(�l���y<�bn�Ym5�B��}Rx� ��f�Q�P����Q���r��ނ���ZƘ�i,��t=��������E���\K ��֑�c��v,~D����*[��'1�4K�P���{:Ek�T���g��6jНa���7к�_t�ªn�%|0����g�[r��m�� X�h ��������o�� I^���~���-9��۝w��N��Ct�yDOe+Fv#9�4Ń4OS���d�Hg���T��� y��t��ZԮ-8e�n*)ݲ��q���S�i�%�2E�s���ti�����7��b���Yq�V�m\�[��OЛ2�ߊN�#�V�+>���2�D��������1�O]����~\�Rszb���qca���6�U'�I�n�c�_��cst+i����#O|�[�5�bp�����U�I3�O&�cS>?qm��uK�՞���bQH-�1yP�/�{��Wcf��v�Ii�aW^�c�|d�>�l��s?ৈ�U���0dQ+�1�@�ႲȽsb-&�*%��֩9A��$�*��yJQ�؁��C��mŹ�շ�q)��ឌ�o.}��N
�zpȥK���aMw��V
�� ̦�ia �Gٞ-�X��E���p�V�*�n�5ɕf�w�[�e\-�a�0��ΡH�����r�־)����G���~�MN���2�\�sL��h��uL4R�ꄫ@m�)g��/9�"onjV��Қ`�A񩜍E�v��i_�k�3u��J�\}R��h%�>��i�H�X�v���	g��4duX�$̀�	(ӐT�<��u�h�9g�	Q�U�	���NY�ki�a5a=$"ݜ�$%>9=h��rpւ�%���a%�O��ղ��,���� �L"�4��v�K��
6��\J������M�+ z
