��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2c=�Q�	��*��������z���7���TE�ތ�2�_����r#t$J��p�+|�r �H�#��K�6����E7ԛ`Vi����0�d�?�ܮ�6����W��U�7w�Ȳ���=���+�
�r$��$���;]A��=�gˢG_S&Ȥ9L��V���\}�^�L�(��넇|�uʦ��������¼(@��>?�x^C��E
����w]��_4A��x��ӡ��������2=���$��!.�@��m�\�3�b�]��h��rl�t����-�W�I �頢)�ǘ^H�Q/c���A}�[���P�D/I�6]M�\�w�\���-�m�Q'��* ��ĸ��W�������n�P˔�7[e,��΀d�p��FO�����"5�Yr�W��2�0��سI�[����s��ݍ�Ѩ���ϩ:Ѿ���Yf/�q�[G�ȍ|�Be<�j�3;�x|X�Z!f�fm�H} bBܠ.6X�S��J�5�yIm�F�7���	bJ�W��e�N�$�E����<?�Dmܦ�'Ѕ�m&�a�8R�%t{t�e~9ڴ�s��j����4�������rй��W���Ȉ�xl4��Օ.}��n����D�E�����:l���+CS����X��XZz*�<!U�A-t�MI� �,w�B`�S�1H��ֳ.%@��[��K�5|�|�6�o�j�l�0D���`{���;E0�^J�}�ݟy�
#���������_�W,�:[޶�N8�cA�Ͳ�E�郭���.��Y$�7l����D:��E��*�#��O�l;�E��F���\�8�'Â��}b�+~h���	��< 7�e�����P�P�|��G�M�i8���P�tP�JA2��9fTʽS��$��a��!Qݦ�V�n!v���G��No�CCe��`­yd3%�>`dg��Beb���N� H��~�n�����垸�0X)6�����ڪ�;�;��~��慄�x�y�蠠�w&�q�@�ƃ��
����U/�YV���0X�v��VY)��Ő�kɴ�+��S�_�D�R-�������>;VR2�➤��X�X�p�*�w��,��&�S;���h�:�2�O5O�%�k��c0�Nُr�A)
 ��0k�À
V+�����4۸��1 �=���J�]��qD ��|S����ϫ���d����+�v��P�]�ēF��
)]{V�)ʢ�r{�)]����NggZ�=�!�H^CEথ�BuxZ-`���x�ۨ��mW�y׫�>��LPGC���[��X"�1@ Z_9�&|uxgq�	D�m��0w0O&�8�^��ț�����!�L�tm��<�r�Zٿ5O�0�Fr�sh��m�hu��70]UF^]Yi;�t�6��.��F�_�� O��t���S���l��'�&�ۙ��P�r\���G�[�P��b��j�e@i���~��D;�N8!�U���ۃa8�
 3
x��mLq����]k+Z�1�R6����sH�$�T�DW��ºe��e�2��	�y/%�g��)�"F��u"q�sw�^�B�������}�Xu�����wq/�[d91l�����2x�j�v�iF��}�oϓ�YG-�cif�=5��-���#d��WD�J7$����%�T�maEZ}��ee�Ǆ�'+���=��(��ɤ\MP��m7Xs%"/_L�Y�?����r@糥�E���|��w5'�f�d��Cܪ�\)�Z۱�F���Jw�y{eN�<�g��k�*&�n�A�D��<7v��J;b�����LRh�I��TkNY�e��O�E���-�ˢ��kS�dO9^+/Ǟ)NX�lhk z��?�@eZs��mT���q����?���XQ�(�}�#ɯ0 �)����b,�۪��1�BE0m����Ό䙭j���(%���X�K$T�"?�{�cGn�l#"���2���6M#+��d�;���Z�p��Q�w�Q��0E�8�q�a�a��[�C�v�Z�c�����������y'L���[�R*7�e� f�>\@�����>�w�D@�d�*�جEr�'ȡU��EN�\��t����G�{�ٚ�:7_����H�$�=�/,*I�ؠ٦�_�����Fp�bS� ?�BSu�9�������,��6�k� 恻�v8�j�
0i����0w�#[�g���.Z���ڍ��Tj��ӟ�Ot�c�0j�?c�MzFJ���7d���!v{O�����fUM�ct}' i���f�.w��ǂTK�{��rˁ�G�i$ �R�;��c�SH�MŎq�w>8���ޚ9��}z���`&�,����R��Y�lǉ
q#8�n�#GtiQ��	��n��'F��O,�d�p4�iH/xi���w��o�*pU"D*�q>+!)|�g���B��B���%q^4��泻,l��bB�0E9�����]����v0oC"tA]^ #�?��&�%k��^Us����xc;ƀ~�Ek G ei�
3'5��GC6�an�iK��Y���'`?	��;T3��s�Z*���攽ba$�yP�lG���!yy�u<��^�Z7�I�#is�Z�vop���N�]�n��#�6�2��'�$�H�:]�&�$��~�0T|_)�;2�5��'�半��sQ�FQ���ɠr�3��r����O݉"�b�T�������8�T�l-�
ϛҔa�[;D�r<W��4�XݺrIE�+|&a{j��X�M	�%҆k��y�̿�ۖߠ\4�(��ي`>߿g�rB����V�_�3	
o3z$	���NS4M�W'F��<=@�ﱕ����1>*�̝���o����X�	.Zu8��(ڶ߲�]$oܱrk�̢���*�����;��忔Z]�����?vl����w�*�k_�V�s������u��J/�CVq�$2
��]Q�P�m�5Vl�[��C�*�BK�4��G�eC,fUL_���a�}kq�SV1"=�� ��^�x��o�lW�]NVSu�7{��A����\��5}k,"8b�Jl)���*.�.����s6�Rjۺ��0��Fa
�8By�򆁸8�p��f_��O-R��ћ��g��A�uo%�����g0#[�HF�5�1P�આ����@���F���+��Xr�������]H_w�&j7�W����a�Oc��/�����_�d: ��&�mlYW��0i/�aOVg��� dͳa�Q%!A������$�>�g
�:W��5�?f#��dk4ى��K�u��Ĵ�_vd�}��t�i	W���)nf�<�&ͅ�����!S[s�xiҘ�����zX�������N��g�k*�`�̄�Y`���;s`:���	�%�"}�8������H�k'�"Z��!�9�)s��h[H�4�tD�b�yE�0��5#��l����:�� !��h��mfU]C�������R�<��H�߬c���j5�O����HzY���~O*U�(��jy9P�{2�G�L �1#�h7T��ͨ|�Wah`e�/K��q�R���S���6i�MI2^�hs�~�<��w;:�����$��l�����,t�y��6�����[좝������oՐv�8ՙ��.a1�V2��eN���K8q˛X^�|:��>M�TU�	�Ђ�������^{Ma���ԫ��K��,�V=
��b��zVJ;�ވ���;(�͋~�UH��L�VK֔�Lb~J�J���	�iږū/�K�Yw��0SP��W��ڡKW��U����<oG�bY��`��E-gy?�[����I�J��9���_V���Y�Ml� ���d!�#���=�tT��(���
��Ӻ�sd�ܟ��Z��r�ӥ'<�KZ�o\#�Q^ܮ:q�F��	�(�|b�����^��"��Wm,[����ǂ�Z�m�tT�TןG}a���?�_N#�yi�D�Q�䖽���tҜ�D�S�9����`gaϟ���&i����o��������S���u�l�{��jA�=�U�tW�Aù�g��D�����'�@L_��@�=;
����[�Z�"���%�-���w�и���G$�x jR �c~X�+.s�Z�>��M#�s�M)J��-..IU	�у0�0ڐ�>�W�Y�|�S��1�N�M�XQ�9��:s2��CL��,��;͐�����Yz%�J�{T{?�����U )�~�Lo��ֺ,H���CF�G�i��lpy/��ЬFi�y�R~��/`��9�K��1��-������T�חf�7<��ϋ���֪B ��z�*�Zj�/���z��gWfz��{���S���j����0��,�Q� �����S-�Ƣr�]
$(ޒ�NO��b��_խ�*�֠j
Q�|���'4<����̿��p]W�L�K$��
H|	4~A�����{�ݹ�Ј�uD꺇���R^���mR0}���ǘ*Kˑ��C�f�
���=m��à��gs��cΓz�IF��������`�:�L(v���	�G��Y���V��:�S���ͮ����ⴼ�j)�{.P�+���4���U�ն���^j���Of�c��V����[�8���h����]���й6��|�����B�@���Q][��S�L]k&扲dQ|z)��8}&�O
p�'�����;�X���	��%vv�/��nL��u���J,$4��f����g-=� �����}>淛���*�V�ա�v�8�R����rU�w�	�6.7,���ha?5� ��UR%ժ����tc#ډ:!�FLK��3ĳ��㪘��|�9%���'�ff�'��.��5n�vlh�ULC1X5�h+�h}�����^���p�����q9����'�h�/zSb^Y�����r��b4�{7�*Su��.,m%����İ��4�����Lo��e{��A.��u4�l����mA�� Wju���a�'�����m�_PaM�E�Yd{��u��\ל:�����;�1�&�hU��~��n�N����|�iWמ]#hgb�v�� Vx���˰<��x����e�� �'��R�f�+8�K��|R,�+�Pkն򤦩e�
V�J�V�?ט�8�Zd6�����������0f�ǉ�*����c�aa���;}�� ׼��O ��/p��b�7�SNpY�11�{�{l�����'FP�f�9�~{�Ń�YFP����$��AO��JT�U�<J�m.!����Lo��`_,�qDFG-#�}���N��_�@��phk��5�\��(A�懙`-G�l��gx*��߹������w'��=ǟ�ȧY����_� �-{U��?_�Sޭw�{>�!�D�l����OOZƳ1���e:�Y8�N���N�QW�����*��E�U�`��]H~^xN�{j@��c�F�N���!�%�)�W�`\��^�rb(����� ��qv���H�_�b7l�?�@�m�G�_�>A��{��0�k�j����rE�i��'c˘F�:���$�ˈ�/9�
�qO�U�ˊ�;��e�)�ǌ�ĸ�	��^"%v ��wVm>�Ҋ��GS�>�Y�+�جT�h*��{�dawH-���´�0��+�WdR���r����Z�b�Ԡ6'RR͉̅'�Au�R����&��)��4r���[R�@��g]�A}iZm|��YHJ8�|�`�������G���w}���d��KI�D��&#�5��b��&:���3�<�xb78�ׁq:�3��H6)��q�Ɣ�G>,o;)׃��MB�7� 1�>H�1^�H]��L�:W�q1�|va�pcjW����rc������85��4����b�n����!�.Nn��i�9�0L��~�Cȋp��,�ӨI�n��eF������ɑ`���� ��y�ͯY�r6�q�q����a�[�Sr*[�%�n�����K�$�?ِ��j�w�ֲ��|=�9Vכt�����|`\�����0kM�#�p�D;��A�p� ��,�ᣀ�O�鏋V>��S�KAb�q�޳��Ml�)o9�BsD���2��٠HO���σ�9�����/d��m�g'�J?�����?l�Q@MU��MfU�p��z�1� JO�T��J�!�v3�jpŧ��PW���d'�u��L�m|��+��T禅��1\%|<�:�z su�oo��'Z)��<�^jf�^���`��l~i��'��E��~Rft���V���8���V5��â��9���}�!�t#��T��Ӊ�0"��=?�]k�`�����w�56�8�k���B���nN��G��;ݥު~P�o���������٨T��*������ӕ�ٹ�K&։�ļ�ՑjZ��7��jU�[Q�f���ɞF�z$�e4��4G��]~�+��n��ŕ栭�*Q-sN��R�v{�"��a�3/��xօ����:�m���ʥ�o8/ ��k��4�/�G�N NN����y��/�o#��������'�*������bÊv,���`�tr�����d��s�����E���s�<f�w���(s����w�)�ZC�l^JＯR8�Y���x�Y�[���C�����7'��S�U�֓o8!�x:�N����KU�Q�/�ֳ��[K/R����#�����%�7k����WH���{�n�Z��%݆T�Ûs��>R��x�`���t��[[M�n��Z�^0z揹���3��gZ�_v�E���lӦ��3�-���C5��iĪ���<��{T��ڼgs՗��T}�T�9+�����Ⱥ��q�����Bf����B���Ӻ�5���^����gq ��,������u@Pe�~�`Y�[��[��P������2��L(s�/"�"��0!	Ζ���P�`7cvi�V�)�7����S#'�Ħb�`��Q�,:�{�|��FnN],���oA��A�s�� E
�`d��xsrrݝ�{���|�#
�O %z�y����,'�_�E	Dj]mpR��v���6�Z'a�ù8���fJȑqu���	�� 兊����ω��Oi�/�|�qk��>6��oy��2���mq��=`zX��`*e��S|��C�Z"��/��q\BYR� Hyfn2SjK'������bv�=ʅ��k�p��q5��̒WS�����x͈�����>N�dϕ��1{Hhbv`��|M�W�6T�+�ƪ�ާ�b���5�¢.��ZHm]<j�����?3��@G'{�j���ь���P���� �_w��p�K�ayx�(�f�����ۈ�BcM[<*i�P7Hx���U���QIꈔ=m�Yna��k-��J�5�E�Ls�5~^�uT���C6��Y�1����0O�����|�F �t���{V2S��	�����E��f�H�]��G���	����l��I/pZ����t��,xQ��H�`SVp��B���tZ��>.!%m�$h�IC�X�\a�6�8i�I�ˎ�6F>��3�3�"
�16Zn<n�̌���Tv��=���u���(*���NF�I��ފ�נ�lx� �C�೘[1�]��w'��7��Û���Ř���&@���������z��R3d�,�=���@���5�P�nZE�>��>������T�&��.�vn�v�����:�5S6�s5��Rp�O�|Y$_��a��M��3e ]��o=�u}�߇]�X��K��n	Lv�(^���Lw0hX_�ߐ��.�[����%/ꭣdj��g��\��'���rI��p�a�I�ڂ�d��3�4^CNTن�e�d��Ov��
��w�U_ª� �{ktb7hy�Y�zM�O����XD5��%�����4�D�$�@��h��
J	��~����da&m_++�ݯ+�����|ج���g�&/�Ц��������`&. ��k�� ߽��4G�bf'��c��8����z�`�d������8s�m�JL=�f�s�feG����Y����h�>({?86��0�������]5�R���!� ���h/�j~�U%ݻ�Ά��G�J���?-*E4�ƴx0���4�j�?%o_�jb���F�dP���h}�M��s��|����LIw��s#��űcy���F�@������s���w�� �H���=�}�ܞeI\e|.����T�c'�G�Ŗ��
h0=>�5�	j~�A����x�{�SMe�	{� E�R�{�lV���R����5�(�:��?�]_m���5�0�/�\Xhs��#9��m�< �?�Zo��y��
)A--.��&�p^/�W�~��6ǊiP-�ć�'����Dָ6�c�[���MTZz\%��~s�#�]��u��m2��?�6�݂���{F4�N6%���bz����5��1α�T���X�|94�=�+�]b�A�p���ݯ쑐�@4)��:�)��9��t&�vM���eI�?	��!�'�z-"㉹��J�\Z�zj�xh_���L�c�ڨkĠ�����*�,o9�@��A�)i����|~���q�v��=L�6�
#Pt�y�@DrLT���w��܂#��pM��r�aBx~�!=�9!�&�E�?ǵH9��e#D�ՅÍ�2׫�"�w~w��>͹bU�Ӂ�5�XO�r^'��c����7S��X^S�·��:�ɟ��S.(V��(��Ӧ#(�{�R
��M��fm�o1#`�*�!gJ��n�jU�K=Ʀ���������Ӌ]+�P�|�v�pC��=Ӈv����#�rE)�J2a�m�CS����	QJ}����=��hLǋ�&5�|����JȺ%- ֒p@r�ү�`5�D��K�;���Q���'�cੰ�� .��)K	NOhŶ�s|�N��|k�s˚pP��e�rM�<J�����4�2�.�x�n���hd�H���� �jOl=jOC[�
+{lA]kC�
�M����������7���&Ҥ�3�tn!���r�LDM�]o�1
8���+������(g"C��yƝ�,�A,]kZ �X�k���s��/���3ϐ�U�12wa�T3�4�z2}$��6�r��1)��]<�~$_��h\!s�Krڻ���˺V��A�m����H��j�鰩��[����!���ҧ����cd�Lx��|Y�e�<��E���!gvs�aOk%���{��]��ި�#m���=yA\<��P�6�r��tPTV�;� -�=��X�:̎��wG�qa&dbn��U�cyʷwW۪�U���؀�X< t+Qk<�z�P��:�G&�B&{�C�*���0-�	�#�������.k����������ʴF�t&tS P��2�<��>ӥ��`�\�8��8��;%��u�e�٫W�<w��~�����QI��+EA�H��
�����1u���F���J�0�/��������S�t.圏��ѱm`ya^4Q��KJ7h ���[P�R����+mٰ9����w�8�Ƨ��)jX�T|�J�NT�u7;������(�0�m�t%ԼM�;t{��b	��;io��&���Ⱦ��}\1�2[��=˽W���`��#����l��Ү�j�g�"�.�S�ҏɚ}�d_sȋtlj�F;v<�pp/��)Ό���JO�*mE�ٷ%R���s�