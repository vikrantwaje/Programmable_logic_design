LIBRARY ieee;
USE ieee.std_logic_1164.all;

 ENTITY mux_2bit_6to1 IS
 PORT (  A,B,C,U, V, W: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 S:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
 M: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
 );
 END mux_2bit_6to1;
 
 ARCHITECTURE Behavior OF mux_2bit_6to1 IS
 begin
 PROCESS(A,B,C,U,V,W,S)
BEGIN
--S_STATUS<=S;
CASE S IS
WHEN "000"=> M<=U;
WHEN "001"=> M<=V;
WHEN "010"=> M<=W;
WHEN "011"=> M<=A;
WHEN "100"=> M<=B;
WHEN "101"=> M<=C;
WHEN "110"=> M<=C;
WHEN "111"=> M<=C;
WHEN OTHERS=>M<=(OTHERS=>'0');
END CASE;
END PROCESS;
 END Behavior;
 
 LIBRARY ieee;
USE ieee.std_logic_1164.all;
  ENTITY char_7seg IS
 PORT ( C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 Display: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
 );
 END char_7seg;
 
 ARCHITECTURE Behavior OF char_7seg IS
 BEGIN
PROCESS(C)
BEGIN
CASE C IS
WHEN "00"=>DISPLAY<="0100001";
WHEN "01"=>DISPLAY<="0000110";
WHEN "10"=>DISPLAY<="1111001";
WHEN "11"=>DISPLAY<="1111111";
WHEN OTHERS=>DISPLAY<=(OTHERS=>'1');
END CASE;
END PROCESS;
 
 END Behavior;
 
 LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB1part6 IS
PORT ( SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
LEDR : OUT  STD_LOGIC_VECTOR(9 DOWNTO 0);
HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) ;
HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0); 
HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) ;
HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX5 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)

);
END ENTITY LAB1part6;

ARCHITECTURE Behavior OF LAB1part6 IS

COMPONENT mux_2bit_6to1
PORT (
S:IN STD_LOGIC_VECTOR(2 DOWNTO 0);  
U, V, W,A,B,C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 M: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
);
END COMPONENT;

COMPONENT char_7seg
PORT
 ( 
 C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 Display: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
 );
 END COMPONENT;
 
 SIGNAL M0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M4 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M5 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL BLANK:STD_LOGIC_VECTOR(1 DOWNTO 0):="11";

 
 BEGIN
 LEDR(9 downto 7)<=SW(9 DOWNTO 7);
 U0: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), SW(5 DOWNTO 4),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),SW(1 DOWNTO 0),SW(3 DOWNTO 2), M0);
 U1: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), SW(3 DOWNTO 2),SW(5 DOWNTO 4),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),SW(1 DOWNTO 0), M1);
 U2: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), SW(1 DOWNTO 0),SW(3 DOWNTO 2),SW(5 DOWNTO 4),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0), M2);
 U3: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), BLANK(1 DOWNTO 0),SW(1 DOWNTO 0),SW(3 DOWNTO 2),SW(5 DOWNTO 4), BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),M3);
 U4: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),SW(1 DOWNTO 0),SW(3 DOWNTO 2),SW(5 DOWNTO 4),BLANK(1 DOWNTO 0), M4);
 U5: mux_2bit_6to1 PORT MAP (SW(9 DOWNTO 7), BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),BLANK(1 DOWNTO 0),SW(1 DOWNTO 0),SW(3 DOWNTO 2),SW(5 DOWNTO 4), M5);


 
 H0: char_7seg PORT MAP (M0, HEX0);
 H1: char_7seg PORT MAP (M1, HEX1);
 H2: char_7seg PORT MAP (M2, HEX2);
 H3: char_7seg PORT MAP (M3, HEX3);
 H4: char_7seg PORT MAP (M4, HEX4);
 H5: char_7seg PORT MAP (M5, HEX5);



 
 END Behavior;
 
