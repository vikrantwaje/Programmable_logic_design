��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�6�'��wm�3q���3����ci�>Ĉ��fo������Ay=4�)�<�P-���Q��F%ANA������lbɞ�<��;����9t|50��d4��y�.�:� {��,B�8�/��
C@*~/��JB_l�2�/�>���i �熲���]lLO���!1I|��s˪��i�hf&���:]�L���1Y(����Ѕ�b��$�0�6rm7��dN�������^G1;�u	6U�J d�L�e�{k�f�x짟hW�P�^�æe����0�&��y4�v>��:w��m�+�P���S��l�\�$	�(���z#{g~nJ�g�%L{:x��A��;#EY��(�a�$YBB�Hؖ����7pT<��S�)G9 u����L�]�ʶчr�d3NKEN�p[����Kj�G�y�R�(p�GSK1%�%o Ā⍁� (��ry�	ԅ[y��,ޙQ�����8	��%�?�����g�}(B�q?�Q7��I���28ہ��^�k���~I��]%<؀���R��0�kA���@��,��C~D�1r�Y��Of�J&m K���WH�|�]�7#ж�c�Ԩ8�^��s{Y�0:S��,x��^��8ց����69p��g��#�'@I?�b<��FK���CL�}�h�����~�X��A�7�X�4�p��A��*i/�kv=w����9�
��Bz��;t�6/	�%��b�)8�nH1�j�W>�+~�*]'ed굘*����!����q�mY��~�� �7pҁ&u��5/� &KFQdL��į���� �	��b62n�j�������:�����[��ݑ�����+ipR��a�fj�Q�欮�mg{��5T�j ��ɋ�v>�_��<�f�C?Tz\W��k�>�>��=g��"��=!��¦*�]y����㶺�-���O�s��jQA�U�ڜQI;�1��nL�:���;Y�:��c
(��������bzw��"��s�,����!h�91�8ǹ��:\3}Zv{E)�
e�ڄ��J���Nw��ؼ(f��!�Ԑ�g~�K�a#M!"]�dLm�gy�*2�.)���EI\yUn}�<.R�Q���0�b��^`�#Q������(�v��z����%�?h��,�S�A%k&kځj&��u��P����k8:����(��Gn�'��=%�mBd�\���u]�JZk�J�� �<Ȯ��$Yey��s@؃P݉>���z��*3�w-.�Hkm[�t��q#}ԉ�䗬�#������Vt���S�DE�g���,gE��^J��oIgc�})k8�,�!����Q������O� ���W�V}��,L273I�p*��0����WD�6S��?��!o�:ْ�	������~�N���h��jf��:*A 4=�eNhL��\H����#��~����;$f��ՙ�&��5��A���W�����>�S #�����H�O_0�;Ϛ�
�+A 8�2��ƍ��
&ĉCm_�\�Ͱقx���I��w�ǆ�A�'�F׉,%�a���yi�����	ډ��y���a��@���by���ʷ�a�jx��'�r+"1�Q,���h3�ף,3�A=�b��``�H��ĕ:vs[`s�������O�DG9#�9�3�Fs=M�Ÿ.*6�����{�V���h�sX`���Y�tpG�r����2B�W����KɘW�Tf&VD򙠈�ߨ*�?��iDe&�M�tC��:*Ņ: ,�̗��R$��S���v�ٱ#��Fj���{���FX��F�3�v�f�\Ӽ�<�P�t���R|�4�`��r�tr	%;�i�����i���L�g�$�E|�|�6����s�1_Y��Кf��s�4�	ql� ���0i���ݻŧ� ���|8:���b?��r�rG�-ۿbU+���UC�F��	�n�<�x�`���iQ�,�hd5�0�3��16��h%d�Py����wz�Ա��v��i��v�T�؈b�{I�ST�d��ta=�It��X�����U6w�خd�F3>vLs�>����p�2��];H� ?N?+��|d|b���'�&!2��D�L �f_[þ�dbJm��|�j�DD�_��C�`��9(f���q�3�Ćv�g�ȣ�1`/Y�+_�y�����=?1�ѓf�u��U��p�L�����^	E�]��΀,��o��#e��~���lJ����R����?J�x���n:z$��v��)�rٗ�#�S�rd�آ�u�}�+a�F�8��%D��1�
T�u4�VD��(��hO�漏5X��3�LFY�!<g����`솨�⩥�����0��ӻ�
'�=�i�e�A���a�����v��C[O��-�П,�G�8y��<����[l������W|#��[ҠX��Z�`?�N-)��[��:����Bs4���Q�s���6nX�=H��E��(�GE�z�Mk)���k}�@�o�_�QK�9O��]�p�H���k1������`#�M����q�&f ���O�б%A�t��V��9��*�L���]:�B�@�I��7%{;�֏<��>=�ˏզ���͏�V<c���,I��ȧQ<{٦�1��y�v��xHw���P��AR�N�6�|T$���b
�,&�#��"9�.�J(�������yh��g,�����2��x�}v�����e���]����P*���R����\R�(��&F����=IJ��.t���T��D���/��c�R�UY�R�����{8,-����E5�]�'��7���I9��ͅ��7��:I��z�u�o��L��Lu���Qh>��f!�*��S��avc���"kM9�[����Զ�|��xzk�p��c �ׇ-�RgF)��!F<2�SU�5���%�u@ �����Y�PF��>
��?�����	�-Pɑh���t[��~i2�߈�}:.Jҟ�*�(L�j����Ȇ�׹�l���D5�+��PFh��նq��]�+v|1�rq��x������'�>\J���D>�*\Kh9�����E�_ޒV�&Ym9�fۏJ�٠���nN"CБ��K��#��U�*pm-�t�������jt�;�V;��QM#��F�@H�o�&q�Hf�O⭑�R���n���wԱ"��u��9��?������B�,@[��D�������`�N}��?���E�	hųZt8���"gr��I��O^~���
�?�V��t�-�O+
w
�#�9� �˟mu��ÎO��vp�u8M���Do<׽���]U��͠F=��EQ���p#M�৹���U�'��3ܦ�y#��Z3�P�nRzD6`He�td:,_u9<��1�u�A�)?�3V�/�C�i��&������D�0y���1�m���V$�M��J��t$�੉�6E��`�&��ju@	�I�����,�6�Ɲ_.�8G4���CM����~�6��!#�>Q�t{/G-��JE��~^���d��
 8�q�f��1����Sϝ(T|4��r���`^��*a��<�ϧ���m;:)���Κ�	���F�4ߥ9�]�N6��S5����Դ%t^a���xO-ޮ	�V;��Ur����b�Vҡ���AMu�O��"/'*�Z%��м�W���,u�~�|�@�fgbL�^�u(�����p*CB�hs�J�8�	�|�C�*i�����9���<��yd'С:+��|qi���ib�8�)b�����+ﴅ���l��龤�,�ڕ��n�sp��Ӧ/����3��s�%�m���F�՘��!<HYˣ�T��6Z��,R�7cS�V��wy���{�嚛��(�Hh}�����b]%�p��w����2��[jHK"��'~� ����|O���S�W��j��a?���&�����T�{h����J�Xj��n�P�؊��z�{��OJ�x��7�[HԄ����z��,�5�O<q���
�~o����C杆���J�{m{R����|$]�d��R����8Q\3"i��������_��a�q�8�Ӆ���݅(�!ђt���9��X��ꊃ'��d�6�ry�f�v�1X9����F!ɭފVd��\�\�;�`�G5[��LTV�py4���mG�R�
L6PwH�W�Ҡd���`9Q�#'�y`�Zzs^i�9�s�B=��]918C�4��<��3��ÖV��DB�$�g��^!(�#���\�U����Eh�Ų|�����~�k��=V--��(]��t���tf�m!�ӵ�>/���7
k��@�!"T�{a��V�~����}%�|��w�v�L��N'��V@���V�aA��1��z��˂�k~�BV�jO5FY!o*�x�*�&B�^���K����o�P?�
��������+��z����SRI��V�y @2���>k��A�?����s�?hS�C~��n�,r�iب���9��X� �Dp�q�rQ��r���[���[Ḻ�O�h�aj\�4ӆ���\a�ìJ��� e�2Ш/��oӟ�ƶ'���\�lm�c��RE?긹�\�[�޵��YN�wݯ���N���H�%��G5{�.�ꮠ>��:A,�i���YȲe���I�E1�F@�&�����\�H=�L�C�6� �_A�T�J:��sg�qW��VUBˈvD���+��H_U����]2��7f�z�op�<
�^saKV	�-H��v����z��\�0����dh%OP ����0���tJ�I<מ�B:"˽�ET�&��w慘�����[�z�q����[�
#������7ݚ^�0W]�lr�%��^.Z�?L>w��%�|�)鐔��~�IQotM�b�u������&�ۊ��[����|J��^�S���f�-S�jQ�H�tmP�˖̌�j�Z@{��ͻ3L�'���D#ʬQ�V�ߛ�-ҍ���'�=9Q���0���i�W{4��,oQE41��OsP�J�:��Қ�ª�@ھ����Mu��쒵�_��:�U| R�[�մ��Az ]Ѥ��7�4o�S�b)�(���}todH��|���&
�_K<{2�!��$H�����j�+Zp	�W@ ��$��=˫�ե�?A�{Tp�@�S3��a�ά�<+�Z��皑����������Ē�,��4�¬p��?Fbh H�rje��~�����܆d%n݅2�=,�4>�.mY$t�����MԱq�	k���\���Nb6�B^x��)�ܝ��bd'��}�MOz\����'h����ɔZ�AXQ@�Ĩ�[_o5��WPp&��C(�E}�A`�(��g*�=�up���5D�>@v��|����l�#�]5k���g��[w��h�'����Q�����s(#Y��Ȁ�C<�3Pk�i,��p�Ў����:Ş'�Wk_����9���ylw.�o�[]�8V�������ېϒ��î��9~��:��B�(�o:���/�q�y����sݵz�a��n>��zˈ�%���Ӊ��W�W�>�zVŴ���(|�^gG��+���%#5��}��a��N����T%�|�%ç���Љ{�=�Y����w�S�
��:$���E�k9S$5ܟ<�Tw��˷��=y���[����4�̅t�O �$1H�Q��{��[��O��M^�ͫ�NK'b�8QL���Fx��=oK�*�~}sz�#f�.a�ɍ�J��	a��b�H�`Ȏ魹I�AG;��8���l0{��賗�!�6�6��Q��N��4غM�E�IdaZ��jX��I�a�>/�=���7sߛ�^�盎�^�99��3���ּ�ZD�ˌe�}`�_�dr���R���Z��~bqi	m�X��Ӥ�Z�O�2��_�����z�H�Ct��(1R���wM�$Ŭ�v���J�c��1��a�Zi)Ur��*ӥ!�u5�qi��!1ז���=�e�-xK��I�1�o������_3��r��A�����I�7R���|	���؎݁C|{��Ub�8ѿ�}Ƀ�aw���: ��ҨM�O�:�Ђ�C>�6?���_}(��61�Rxy}�����np�̓א	&{�sn2T���Ѿ8���X��p�2ߒ�\&�%nJ��m�S5�|w�ۂ7N��@���Tؤ�î�:�'�Q���ԡ��<��׏N�)�E������S�"����1���X�{�����JO����T��i��CwX5Qb����ۼyO�:�|��
��5�m&8kO��d ɟU]B��8PIV���{34׺~��W�u[�3����݊�<�E�O~��8rNZ@0*�٩m%��g�s�08�ĝ2��%Ӏ4`V��~wr8�/k�Z��({���)�y��n�(^��Y�����a::��ό��JF���#�����P���}��47��Q�������p�.��i��<=fy�$�B����;��M��������\llR���'O��Zv祃�(��!{ȮW�<�%˲Q���*�Z��c��k��
j���\v��xB.C\��+����+��\�/�=��Fb��J�Ez��Fo�
���� �gs��|OH�����\�9�W��pǠ��BU�@�	&K���i����H����k�lP�`�r���ʍ{$�T�=���?M� h�4�i��=�֡X�Zv�u�aE��s��|͊�0Y��ME	kӍN�ЎV7T՚qN�C���=���%��Qș?+���ߝ�PL�)���0�ObKF��^H-EQDL�ys��J~?��0����D\o��c��}��<�	�K�U5������N�{�SW��sϖ~0)K�u����\C��:��\;��T�y�zވ UV���D��o�RA�P���!O�F�L��Ys������T@?�/G�������
Z),DMi��։��P�Q��ێ�i�쮠�c����>��������u�0�S{`�J#����J�?�PU,�������M~ʜX�ud4V���ƚ������_�����P�l�]h�,#@ת��7�q��5uf|w��č��|�ɜ���T��N��oj�H����E�N\v�Xic�A^�|`�53
�G	d�� L�%���B�pO��υ\I�1��e���`D�D�;�S$�5�:q��c2N�H:��%DX�	�b��ճ�k� {����t�\Ho�otf���8��`��e��l`�;n�	��J��5�9�4�q��}�=����y+@C��h,%[��7�W�Ο/>ާ���Js�g��9��!��?Q|�$��}$�8|$�if`�ȟ����j=TqV��s��˫�Xω̻:c�~��0�̽�"�l�=l__��g�H7������]�'}��FJ��kZ���+�^���� ���N~�ʖ�o����H/fP}G����6�J�֙���g����9Y58I�M�D%�.~5�+�2��K>{q��@�q;�0i6��-�j;����n���0��|&����#HF)5D�5���>��l�kм�YN��
Z,��d�%s�uZ�f��|���BWx1��� ����;�mC'Vpd�{VX��:�< @N��P�����"���0iz֫0^ȶ:���w>7
��a��Ed� �.Q��6��{���#��:�8,����`��ɌP*�j%>|���J���2?����^>��9�1�f�n0�I��z���Z/.��<�i\�b9F�xaf��B��GF��=探-�6�y��s[��([���~��8�m����Y��. [c�huIZ�ĚpͫH1��n"�����tĮ�-�J���v[R�vV9�6m���˺�v��9G$�+��[��~��Y2��^�Q3�>� �|3��i�CZۇ�vEf�Z�}��(ޝ<v�@�I��<����9K�}I�Q� ˙��|k�*=��U@PGQ��1#�4B3�6h�{�z�eqb.�u�q�z��i82�,�z*��;��@KhR~�wQ�&�d�ZY�P�ׅ�`
�����c�ե;�/R����j���W��o�ip�EPӣ��H |��z:��s̬�N�z���}�O�Wؓ�����heMo�.[�ǅ�${ ox�ǭx_����,Q$�-��5n��h+�5�.�����Ju�A���l�bW�xƘy�F���j�4Hg�P�Z���O��=Y%�"e� �����fwu�ӒSg[LK�8�Z��ׯ�"8��rJZ��&r��:j�@�č�Dg�>,4*�]�UǢ�.��Y�O��'d����!�\� �ǚ��!��ҟp��S����4|�<��B����DǛ�Jľ�}���2~�YwL$�,Ц4����^L�a��LV��ĸ1t��{�:�'�=Y\̱��w�V��y+h� �(W'."��j�tN�%���2��D:���������&����l 9��N?Q��q����"v=Z�Y]�H���M#kL#�:��?'џ�@u@S�*'�3 )z������y.Qݭǡil�l���;���;5�|�"+먱I��G����g����j	T(̛���S��q`F�9f�T��|K��0m�2���g$<?�d���O��\ue��D\��~��r�(�;�䢛=ҹv�sg�Ү���-��E��_�l|�!Fj_�^|	����s3>����ME��WWuc�Nty
�/���d�x�jƓ�DZf�b�R���]��]��H*�U��~bT�\z��k��s��*ޫuΞ�k������<{�K龘�Ԛ�V��?�[zU��^���}�l��j�ild��T����n�6wH��Y�O����gRo��O���	��D�ҥ�n��CO����		!�U�'q�yAɥ�	�/d�(�r���Kkį�oԥ�ٍӽ�܎;�.:h�O��p7�&���^gG��PS;���ݦ�a|jI��\��E����	�=/5�P�����*T�7��!�&a���f�ʴ�Hd�`�B*�+v���W�˩!�� �Q�9����r0��	��f���	��֒}��:<�6k�A=y��&�i@�v�nx�鿳.elqR+%�d��:`�D��~�p���E��7�(}ЋF��1C�^D�z����yN�4\5��	?��>ҩǨ��/5��g|��Fd�5�0�E��%�"�v���"֑rs�Lƕ)r2�7�n�Gr�vuVCRpT�qo���-U��������{�~�PT���A�ə`����C�{�A�X6�n���jpy�gq'��T����n������H���c_<p	C??�X����M�W;�!Q&���:9��A�D����"/¡ڧ]AMQ�7aŸ�o(���@
kz�g%��S11��x��� �)M���<t=��Xg�[�	N��&�vd��.�H[�3�0�R�S�{$�eY q���y �V���?|�����!��
&Jy� {���t<�kK��k����$Kzs�
��<#�І�����EP[_E�2i�|�J���c0�_�`�5B� ;���V��87ށ��Q����Ї�����SZ�G�k���R4�K�l�#�A.Br����0L���c�EK�NW����{JP}Bgl�T�[7�e�(t	z�̊�/�L�!��7�Bh
"Y�Q�>ޱ*��X�x��P��Ȣ�d�m1Yh�� ��338���WZ��S���� Uv�
�� V��<�l�;�^���� apk�x�,�8+�MT�" �|s��V���凹<(�Z��*����*>}Dٮb�4��65F��_����Ƌ��p0��D��Z������1� y_��ِ�*5�p�4�V؍Όg���2��}e���ʙ� (�\@�W�>6#�|�b^��*f<e�g���s�bպl��HX�EUEXG��?�3�
��nG�R=��"��׈��h��K�:�+��{X�ګ���I�Aòz��I�!�ARd�� hZ�Q"�_k�S9�k�2�����Im'���?����� � C�&f�+�Jvf��'O�l�s�)P��1s8��� ��}���{�L����~F3�Un��k[B�7���k�����~Y~Q���މ-8 f�B�@\ӡ�5펃�z�v�1���Y��m�>�{TƖ
@�����,gX�s�dtNJ���ٴ��p�DY� _�v��AJDn� .����Y��n�����3����@_�x����G��k��x�{%�~���ީ��i��;�r�SAՏ�"Y���N����C��v�!�N�l��+{�h3!a�W���Jb�]Zs��||�E.'C:�4��㷥�G�b ���.���+�{Iց��j�GU�_��Mv��}�=�Ya�>��.XP�bz�%��c*d��?i��eL�̐H+jJ�O����o��C�T��2n�Qrh��}���G���]Y�6?��D���dGD�W2�p�m��[٤��9q���-[%Y�C��:q6s�%}�Ç4q_��x{pX�MI�C{ML�H�,�M�w��~u�k@	�*�pI�סּ'���2<�C�L��^-^�B��N,VٕM-ݗ��|hS�����^鹡�����J�����AF~��Hn����|s�G����S��v��)7L�����1���`V�"JDn�=��q! C.5�7H�t���������gب��a�"�Έ+��
�:�YF�Ū�F�P{��`-v{�@�d��\����^� D�ɦ��e����B( $�q�G�ެ�W��	˂�F½�!�2��-}܂-`�'��U��n�J[�<�u���#_��5L;Ni]��[��~Ԑ��t �/��2= ���#��@Ѻ���!"�Kl�6�q��d|�wW-;���w$��|�~�nSn0���Ҙ�;v���2
��A�Q�M</�U����ٕj��lS��n�=6L�ħ���7�zR-�&�����*ǥ?�����xu{������:���:��/�`,�N$q+��;��Vs>�%��D�3؊�n��gR޹��ԋZ�7o#b}�4LY�-Ϛ�Gj�9ML�z��c�Ldە�-����i�:�����n��[�7�+��?;�����aD�9
��Dt���W����<p�(㥍(��ʕ�K�ea��BG�B-d�����m1t�]�z_p+nw�=��U-:���i�w����Nu��k�� R��'d���0�T�{��BR޲����-~UΙ<G��)mc�!����Xlf���P��W��g=���
i�T���<�A���0#b��[��'Pd�+HQ�ސ�GL��JR���M�ӱ]�[y�ǘ�PPLH5�xO��S��'c��漦U�B�&��Qοm��]
d����2�F1�.�������_R�C��Kզ�k=��<| ����*�v�W������!����-|���Ҙ������,�u�X;?�l����F�c Y��o��Ԧ�G��w��A�#���<�D|u���BQ�@S�AN0/̺MSP�g�r�I�Gp����=���<1R�՛PwTp��;!l(:F�e��AeՔm����v��N2�4U�ˬȨ�̟����TN~E�ѝO� ��N��8L���V��kN��o�Z$N����!��(?�� q�çF
�x����Cr����쩿��h���d��Jj�áKT��2vw��ڦ��6�~*eB�4_L�E{#��i�~U�wF��<lBz�s�K����|L����C����0�ދ����:@F�Xx*R�l-�"j���R{H�bi��8|9�/�)�M���Y�9��)���4v�:�vs/Z�h��N�a��3z�Ԝg�Q�P���-f�-ĸ���쥓����*U@�YI2��ZsV��/9y�l�뒳F^�/�^*�}p���#e�d�s�f`��w��]�\5��ęG�v�W )�͐S��T�w$�	�`���8�/>�wQK��{6n�a� �\kXS�]�45[�����+iJ�~P���w�t�s�v���0	*��.E�m�pE�1@�.<B��ߝ�5�
�E�p�ς}
K�Pg����&�+$�YKt}����֙�V�{@ qtA�گ4 u{M��R��]� �:�
�f��LOX W@�y�z�U�<�sN�i�qU�m��I?7.��ܳ�UQEhǅ2�܉(!C�nKɝ8VfZ;#��U� ��'Ý���bbJt^7�I�ї^��U��ܱ_l�GH���Y�m�aj,:�B�ף�g[݇��#���^�R���#!0|��]P�� �%����3�%7�A�,�3dj�j���0�_�����/2���.��WS�,�J]�-ك�ո}ܰZ���b�=*5ʀ�cD����S���$=V�q�쎗Ƈ�HR��c"�R%����Ȭ�;�
-�Qab�~~(�HN�7�g7�"k��K�=rY�Es�%l�;W�	>���e2X��m7��g�wǾ݁q�s���l���,Θ�)�L��l-�/���6u�'H�͉մFa9 �6%��hV�:��4%��ߓVɸ��p4m�{g% ն��j�Tc��� 	v[�~`!B� N���Z�>3��6L0�C/�L�~� �r�=j0`�/.�7�ծŬ��F� /�l�^moH��0�_�W�.�yo#ڦ���b$�#�~�-$���D�?$K����j�V�j� �� T4���8arS�5��xܦ�<\�vN3�`O��E��;?� &O�'�:D9��@�e�n��ki�X���H�'/��~e�)��"�ӫ`Q�6@C��w!<��S��ۙ �	f�sg�6ѡx?�~��Ћ�19����}�{��5���VA%�Ʃ���ʭ���B��H&�.��s�&�X�0�Ϫ9po?��ǆ:]���/�PWR���@�XA�kL0�L�T��J3��n�+6��,��\��	����(�2x�X@��ȟMl�`����c� m{�]k�k%JQ: ? ���l�!M�����/+0�/MZ���fȤ|��w4 ���ٶo㺲��Ԗ=H7���ÅF��hZ�������tܮ�1�Eu����i	����W�ȶ	7��k7@�N�%���k]\ �q����?�qZ���PC�k�610�NRk��O��ǹ>���k=��v�c�A����M�s��?�N"dp���i����t�}�g��t��aW��?�N�}���BU3�U����7�����ǘM�|}&��,a�,�.b �$��\�2n�X��~^���6_�cw���	1��+�D#�p|u[]Z���jl����¤e�u�?\�*�� 7Y��5���2!����;�}���N*eMï�I��)�=�#�%�%Z�A�_<l�Bg3���o�Gkd�,����:��Ј;A7� �P�H��5d}�u��7����Q2[�mq4R�!�����ec~�%~CW��r`����V�Sw1,��H%���,~��
� �+K�ӕ ġ-��|����*��U"�*hT�D/c�"+�yP��1��i����@���wf�i���V�~�졅6s3���I{h�u�m�Rg���i�Q<D���7�&!'m�ݿ�K�E�:)�Kb ED���&��k�د]�Фc���9ZD)p�%���FU!�2���9�ǭd�]� �T[�Ԕi�
�_]|���FH�8;ȳ���F�9�%��LC�����l`YRYv�s�;�g�`sJ�����&��o<L�����g�7A�]Ƣ-��麢��$�%�����皘�@�T�T5�jZ;��b�!��p��τ<R�Nf�x<V�dp�aPr��j���kQK?�T�L���J/���ﶒM>��+���E���͵���]V�X{��g%�iK�/�J����z�B9EH@����2`�����\mW�7�:������[C�c���ΟZ��q�����p_+a���ש�$�a�$�Ri�M1�Q��]S!#?��v��4��k��1�v��	�G�ףrU�:�)���F�dFK���m�Y�n�i�\P9�jι����AD-�H�e{ &�	W	�<Z�q*���L<N�ֿ\q���GS��B3�w5�N�n�c���%�{,8*T�h���+#�]`gŗ��g/G�q����h��?���υ*y$�C6�0&?ӅԲ���A�ݗ��!�G�$�@�G�'��J4` }�a��2D��H����M�>��5�&���^ģ�����o����� F�i �y��_D(*z]��y��L��="9_�qA0ѱ��u/�z�_���$g�T���Fi��XS���R�O\��C�C�c#�*x�ǣA(^���`y��*@|O�4W�v�T]�:�ova��Y������)ԥ�4�I۶m�d�%�����#���N��6�KI�S�3��ʯ91>$�I�*Jx�CF֒l+>M��fw�E-W�o�.���\j府���vF+5J������������S�"߽��l=�A�u:/X����|�l��K|m����t�Pd@@_�l}�S��,\��o�ѣRZ����W*��hYN�p(�o%Ym%�ן�^F�\��<lP��ꪵ�ۀ�w�����|80^yT4��E��8�J��و���|�(�;ʘ�6�ė�U�td�Se�R���'cHo�w(f�<x"�η�.)29Ux�p���a扼9or�7��.�f���~��EE��;4�V�u�^�oˊ��4��=�};��9aq$s?�B��5����I}��T�{���ti���{7�K��M��{�
���Y�+������u�8%�ɶ(똀[�T���)��z��5����e��^��}����?�@�/�*��d�=�y���˟@\_nuKjI�,pj�
�-�g�h�� ���GҮ|d[3�.u�A�i�VW�%1X(���3��
��aIMlz�� ��W��܎Hs�Rv���4!�	��>yz�6�ʤfsܒZ��d��v(p�>� ���k9tfE&1e����ZXk�0�O���W�G3�Ƭ(�=��5+�i-g%en��ڇ�^U+�9s�w����r����JiB|(�S�xOS����oKǛԆ��S@-�vX�05Ht�g�Yx�/�����S�"�L�MR�=U�Tx����[��@�g0�b�*��ii�0�W�� ���my[R0�Jv�ƌ��ap­�Y4�k^�1Z�-�RP��GhV���'ot�-.�-�b8�?\ǓG�J�v�2Hs)��?��H��y�����jD��J�e>���@	� ��v�6Z�Dh�71K6�5�ǐ��I<5K�fP�[����X�� ��rU5Xa7P��.��GF�$2�Z~V�V0F�'���6�vGM#$.:��,�V{��lx(��r���N�Pr�
�hi[��w�32L�~<HG���j�}/�,���$-xb=I��A&Q��w�S R���tH#�C�cΔ���Y��oq��h)/,W#F<L�8\�e92|Rk2W;�]^��
Sk�sU�Ad�i��S�늩*]3����1/j�X/�j�]����	���h�آ�"�f������+$��tkl9.��C�Qb}Á�qZ���$2�I�1����!Mq��m�0p����G�i�xƁCVΌ����jW�oϳ�L��=�j~�}�5��R"4��>~������.Yγ�D��^!�e@��b��PR�u����K��4�+P�hf;��k�0P���T".[a6gO$��1�8�f,i�	����� Yjym�f/*�����g�,�1X�} 7�W���s�D_�(���VV9�u��K��u�.̐Q<O{������|�~��t� 3SsO�}���2F��S" �������M�P��8gLvO�1����d���ǲ#�僴�H"� C�W�mt�{*�G�LČ�g�k��ˀ�/.!��5r���Mp���/xr�w����2,M�t�h�
�8\t|����dt��u��i^��l�ܪ����t�c{�����u��b�
w��;*ja�H�4��پR`�V^�s�*7/�ш�f�3��P�g$Wf���'��'�A�R�5�i����f����=ޜ��͛>����^���%���"'G�N��.�w{lbܞ�N�g�=��h�����5}�G�4�e���|il��N��~CcdUZ�.�7kb��oh�SPS⿺]�_����,��^N{��5h���@0�0	�i~m�b�`�=Ѹ���B�з���H��~�u�]��ܸ�Y��[K1��Yh<�z�]��3��|�\ܾ9V{��X��	�h�=f_Wx'��z-�j�O��ԸK���e���6�?�"�����%�U=�=�Lgӡ��p4�1g�.�Թ_���J>��J��ûGe���Ľ��V������iv��|�v�ƌ*���>s��i/���T����?c�$�p<�.`��ҷ\
`i1M�����T��Qо��NS��*��J���zy�8P�rC�N ���%�5�����ᶙ���"H1Z��M�*��΃.Ǜ��S�[��d�R�<�Z&��񍺫1�R�@D����VO} ��N&5��8
G�i��5���TX`~4%[�4�p8i�'|�q?���rk�z�}U	�O�D���Zm	�J$i������T4��$�&�� �u���^���,��|�Ă����X��ԩ�j�>��Q�|�(��C� `Nw��D|,[��Gp� ^r�y�j����X�Lt<�l{]cWe9��blʦ�=���$l8UW߄�ĝ����ی����͌ ��� L!5
Ƹ��$��3�3�d׉�+x�e�zO)�VV1{�υ//>�����/'���(E�p���o?y?��rFE�MA���X4�Zo��t*��c���I���G�k���RI3��W�}��+�t�j9�k����`���p�XŁ�?@�an*f��@�����i�-kFm	�|g��5n���>DqC7q��X]7�mr�!���z3����i0j��걪|�=߻���N�vHG,�,���&��ǄXc�����������<�I���gk�W�=[�:�/!o֭���tXH���M^݊ƣ�S׺�� P.uy��o����(˝E	�m���ܿ;�\I�FZ141���9J�Is�gb֩E���N�m�n���,+���o�z�B�f��1�4�p���O'����|m��^�p_�/��o�#k�W��)^y�H�2��7=�+K�r=�A�mu��A��>F'��a2���:�������7��>d�ul|ou�X��qj�qʩNs�@2�/�q��P����!��rX[�o�r�_�
��`�a��wa��ؓ������M0;����֐Mn"��b��-�4�\��8�����P��$8ɻC"�V��HC5Ǉ��p4X$A6c�P��N�qVl�؞�^��ޡ�[����#3�1m���(�(��?y���B��A��
;�=��g��CC��8���3�g�?f�:����bvv
Tc�Zޠ:�xd��',�����+�@� �1z��A	D���Y����/2�C�3��2i'*����� r�0l(�q��("��l ��`s�J*��0r��l:�A���y�6���%�U� �g�M?�"J�]�O��<o���#�Ҿ��:�1���U6�ź��'+'{Ř�Od���C�/#x�.�!�d���+C�eڠ��Z���3�`�O�("'k&���� ��)�SD�f��1���2_�|W�,�$p��;�l+S�O+����@Vr��&T�礦.Y��*	�s�GSa����~�q@�Y��ҁ��;4�޾b�jH�(�ug�_�nwG�� �@��F��zp����,��	oLp�-��a�u`���ZwNO�w�U+�b���sX_�&�����8�"�9[/�E�����m�kÈcC�{��tr�#ݓq|I�?x�'�?�C�WG�+����J^zYl��� �S9��s�䁦�y�ჺ$���|q�8\)EH��U���z�O��%�0l�.'���Gv�$�d'm����O�=¦G0��ʥ��s3.b=��?Y�s1?��T�t��q���1�1�怟����y
��8=�ǳ����Q`5�Ϫ6%m&3������h����L!`_�\��R�\�>?���/�6�t#{ �*� LpO�?u�I�诺L�MJn�:�H��o��)��������O����%G��@��x����*f��3)�M���!n_va1/7���������4݋v���4ۆ�R��q筺f�m% �425d�<�+%y||���7K]2�;��������Uk��yo��Ľ��ڌ�5�Pt���-�$T`sh��[��Ŗ��}�d��Z:�j@�Xh[��Cf5�]�֠��aN��Mgb��b�ŦO^h�)�d��O$��j�2ėY��|�]�"[�-�|������㛮��Yq�3� Q�)�;&k)���ʨ�����-��dnQ�A^O�k��Z
���ª��G��o�M�������e3��p�;�N:����m�]"`��y�"'��m����kF�F��s��J==F��f�<T��$��h��\*�[�Ƴ���1�
��8;��/����E��<#��|5k%Վ��� 0��k��
6�lh��3�e�� GG���7BG�1��&v���q���g�#�SP.��Yfԧ���J��e���~U�;�	�ʹ53>d���M�
�O�!��<ьؿ�.��T1r�QȀ���,��	.i?�e��ޠ�IRB����Mt�sM4�  �j1�C����y����=�p;�^��MB1�rYU�I(��E�'��dn�x�I�����:�Z��8�88u]v2�В�~�jn�E����g<�9��u��'õ�eh�!.�uX����.̎�8����00�#�*�ˤzn.'��jG�ci6u!��~�;O���{��I�s�"���p4]��/��Q����Mj}�w1�LE\�g$a�+j��]o���CI{:[E/��	�~)j�?a��-�:���wP��S����~
���=�Fqj������m��n�տ�z]�C��*�0qH^�־p����"sYG��U�tU\���5��?�8Q�Fd�
9�P-"tR�,91u�!��a�= �o*����|vO5vڒY���,G�w�����t������7������]l>���@ ��SyY�o�_���e!���!��K|9dZ����d�S��)Yȱ��o��T�{�x� [U��F��[����N.J*��3jc��2�V�7�z�9}^�c,�[m�fZJ��Cs\µ�p(��<%ǅ3 o$jj�}�����?lX]��|׃Y���<K�ﷵ����g	>wU�ǥq��%�?7 ��qo�fP<����)�U��f�E��ۓ5S����]hV�9M��~l��Z�0�вj�eZ�{TwЙj����KI	�8���_f6=�����$�h9yq��$�1�z����8��0�}�<i�İ�G&�� �;����p�)�X�fJ�(��"�d'
���J����H~ƉLv�ף��SP귰�8ъ�\)�}-I��a^$�>�Q�g�44��6��3S�W���	���z%���_�=����Y��gvǱ���,�����ơ	}�����&�H����%�9����Ќ��$Z�-!ȋ�����E��?YR����ʙu�a�x\��Z6�%�˙���8'�|I�$���ٴS3�l�;݊���?~t�$I2K���] -y�N"���\��@qH�B��Eֵhܝu�e]&m��v u�%j�&�VwݝXzL ׬��;(�8M��=U#��?����)ˎ{��,��X9���Ay�%�U�*�a����"�欽Ƃ�/x�e���*,VNP��c75M�X�n�%�'t�/���ek��0�m�V�T�L~�h���b��[� �u)��
Y�I$ty!:�����Γ/G}�S��G���Ҡ�|<�t��0\1�:�,��(���E^yr,�(T��_b��\2A�v�Gz}�KN�w��L��:���$�?��ޘ�Y�H����EkC��s��>��B�A\�h�bVf(��^��bCR<�Q¯L�N����ɬ2��=�{h�e��W�X�̕+:n�g���fI7R�Y�)kr�2���	 �ׇD�訋��f��z�r���`z�qh^��3e��-���g:C8��;���D���A}�x���L�=�ɮx��0���e�䲯[����T��`�ǫѢr%��65M�)U�_1�;(HVV�݆	�\��c8&�Ή����O�ߑ� i��m�o1.��Р���"}��k�Y�!UHr��{S�y9_�"���kW��0�晵_T���9�&�U�?��LF���
l�<��ٝ�[�9��]�k̴4,J�Q��ͮ��]$��7f֦!����0R����0z�%��E��ĭ���WW�����2�4������D���>���8>�EU��r ��"�$��8�V~���6v�G�O+`�IQ@cr�=\IL3F�Y%�6#���:Uvs�B���������A�!m��g����jvX�;�a[6�鑺X#�V�V�����8K���;A�p��$��J���h	��^!�UK�kP��t�4ψiI�%�>X�Əo�kGI�ߪqb���]��L����%�yy\e�^ܡ�"o�'���r��v�����Xȅ���!�� T����|���M�9��x� �Z�L�ʒ���M���Ӓ���o�%� ��A�	k?������Co��ԭF���kGn@�T��{�#Ɵ��ݧ���Є[ׄ0�2.
[6�7j�fc�J�9!�9\�A�Y��g��	�H�Tɋ�}����"����Xfc3�<ʔp�t��ך�4R�79J|�-1]{O��δ�����B*��`�{������o���;�|$�@��1�k/p��yGue��h䕤=� +?�5;*MFR�(7	I���L�Z)M���U�~�b�8��07Cf�9��{s�¨dB��m�A��ݔԙ�h�v��5cm��F���&��f�s�T�dv�M!��������`�:���uBX9�q���6���sz����V�l.\�������9РaJ���{iӸ�x|�!��+����3��s؛׬�a��R�M�2��3_j��Q3&���ݣ�����Mֳ���3� ����_��#��M)�)��i�����.���t7� 9�~[ (�e��?��U�ob��J-�A�"(�Fwg��$��ٟsM7����o�`8�%m\�2_D`�b���$R�5�� {o�'��K	�ݧ��ܪ@k"9����)˽��ĩR���T�� �L��`��ŐJ=�CAVmk�T�_�"pfK?i�e>��� n!%�>��?7^˞��ͨ�a;�����X����f��<�d�C�q�q������j���t[�Lƨ��ʓP�(3��G�[H}l�P�ۘh�u����+ 1�N2���ol7j���d�?�b�����uy�|N�^sa��ksȀ	fto��Ϫ�3��񅗵���3n�q��3�xXKXމ��i�C���U�I�'���&
n�ޅ���a�0ܝպ��f�I�W߆<=�h��S<����"f��X����BM��5�prM��<�]�I��ZŲ�J)Um�x�3<�0�V(��Wp�e���W�^ډ��ǀB9�l�#�(?�梾 f�`�o{Q�fV5R"/�^`?�I�S��vO_H:�L�O����|y�17L�7q歃y9���ԺTT�����{`:j1eFtm���	r֛Ǳ�G���$����ۨ��i:,w�����#ڠ�lrH�(�Ņ�P�̄�Z^���A�}���d�Q~�_;S|�hPD�8�[���WD�>Lf��0v���-o)�{�[�"�3W��*�0��c
�|�`����|7�a���]�"�z�%Oڜ�d�Wa\�g�	����se������,Y�Q@��;�uXJܿᩮ]z����� H�?��P�3�(!NN���e'�zA�B�z��|��Mš[p�	�ZcҼ��,k� ����H���]������6`��1T����ڠ��FkC��YLg�զB:��^Y'C�+��..]/͈�
��GCz�}�ӵ�JK{���'�FA�;��6���Y]��J�p�K�`[����6�p�U��\��Kyb�>M'4��H_pA�',���lw6���#a(�+�vG�^�~)[�Wr]8~��Z���d��o��9l[�s�Z~h=%qA���¸��]#g�ѬQ�w�w��=)�a�Kԇ��(���΋��l�ϣ���bb�����U"�
FH�^���.�R�إ�cޱ�(�X�l>Y�JCd���~��-�eꪃ�G�	PH�EK�-����Z̊��~jtXRn�e��
[�=�X�78�<��ؙ�ڪ*���C��Z�)à@._���wP�����0m�r���KPݗ���~jJӶ����V��xh]��T3p?@l©E����҆�(&)�PВ���Y�S�\N��7%yw-:s(�P~.oXDǶ��o��	���|	2^�4		�4�)&���^�g��Q��6~o{��]J-"B����:w'������b�Z�=8���ٙ'��g��7.�U��TW+���k�%��~JU��������/��v}n-?s�Zz Ã:}�T��fn�e�s�yK]f=�m��܋��t����܄@[�0�����%7�GK�^@���Z>��V`��/}�&x+��:����%��ք�����N��Ŗ��@\�r�rVB���c_l5'�����3�o�&kn�܎��A��ʶ�k�[�����[��b�#mě�uW�YM��šy�/䏩���1��~��C)�7�M�_���Ph�w:��d��!��e8���IS���$�}�o.��xHh�����C�c�S�j���jm|�/�E�m"Y�r2E���
߹�.*����g��&u����Y�YD"\�q���t��(�1c�r[����u,�v�
A��r(��Y&��`��YAEl��b?I䳷C��?�q.2ɜ7�.0�2�MP��.e��/�+z�Q62*�h�c��R?�Y$��KoI��A�cB�<v������s�0rd���4����o%37�uc���(��E�Ln:䖧4��E�JB�����ȣ���(� ���czMij4�Ow|�(k�ps܏0]�s��4��H����s"����(�H�fH�V\68���=9� 85yɑ|!G�Y(�.w�P[R�C_�N���(4��];-�����L�-�9�}EN��p���
SJ,@��Z!��@�3�_oG����4e&b�L�-� ֟n!�A��M���0Ws�da�7��_`/H�`	R	��4�=��+�=�y>��o�q̅Ľ����0k���h��-D��2�xl��,s��M�z�1l��O�"7:�9�غ�����p���N�t@Jz� X���������Ԥ�x�C�щ��0/��{㞪W���G��*�z�HVu��9ܪBC���-o�N����ٷ�~�s�$~"2�N={�m�V\��G����(v
�5 �� *�.��a�b����)TP��4� �GQ�Ȱ��t��
}�C� 7�Q�!\:��g�w�X&N�ZG�R�n���i��Qh��:~�e'o�\10�P��Z�}��[
����i��pG5ճ݇3���q���{�8����/�7��c�)+�?/���Cl�ĺ�!\2'g,�*N���ܣ
��0������>��YRv� 6�V���P���Bo%�rI�Y�u�GBաrD� 3��4��q�
�)�����ն2�{b�^2�4����=j[-<Qh��ǿ�b����V+��`N#j���#IRr��� Ɓ{�|�֥s���R�J�P�U,����'�)����sBcc�:T�2d�nCǽJ���ұ}�!GP��w�gm�=�1F��a�+�奮du�P�����%�������+��9��s�L�e�U�V���������a��|/��W��m5x(�dE��u� ������ϼ9M�T~�9n��
rn���/���]����q�zMq���&������o��zҀ�<#� ���正p�l�5Y�F�/,ʭ��OE<��_�{�r1*�j�#�& �{��ͅx��z؉$LhP{�-)麊Ǐ����(�$`��3nG��8���Sy؊����Vp�]{L.ѽ��ˆ��+P2���-G
旲�����3�K)�[QɜU�L-�|��!W�{;� ��g�Ta_���/�!P���������S��H���L���.F� 
�/%H>��
m����S1����W�#j�'�EXb�zV)�b��|Jw��8����]�֙\��-۞�:~LS�1m�¢�ї�S�^è��T�	�1T�q[��wų�?A�ˢ��BΛ�L~�#A��id��2�6;�$Qy�Zr��E~����Xի}���\��4�B#��徘��x��'\sA�t�h�<��:!��(�t�#���#m�o~�m�v\��a��V�iuSA�Q�9<��y���Em������["K���'���C��>���L�H��B&.��lw� ��Ĭ�1A�+̈$���jO�/��m��ܲsk\�n�꩓���PI��0���3�����x?X��)�.�_z�������c��2'~�p,��\V[�3��!��ﴦ���û�bӏ���k`�F���\����<c��\��tYix;���*�#��{�8?_���nb:>��P���F�[_�D{Um-	}�\&�$��Ý"f����P�J�{E��H6Xd�;���+B�z�/���!z��o-�_�5���k#��Z&��=G
ua}$����]����N�'��6'"�E��r.��,��'�dN�R3�,�$�}k\�֘AGX�&cM��M�ף����ɉYo�����)1�D��1�y �c�+dP5-~��1���W��]]JE�5����-��94�f$@'Yc��?]�ɻm�RH� �E%�l1�K���?�hU^X���Ua)L����)}36*����67Iy�g���o�)*E�5��!_��#�϶0BS�i��]��y)����z��Z�EV�y�������
5�L2Nb]˔��zʸ�J~��(�L�@2�>�Z�����dt��5NT�K��P��I���h�I�U�N��`̈́���&6�����n>�*������0���_�B��)���7=#h͂ə��ŵ��3��4�6��ɂ�d�4���qvC�Tt0���4�wi��Mg�2zydrEx���	�+�r�I�>Ys��/�Q#�
~Bq�)� �x��bu��.�ɤ}~\�݅�lG�;#�M��q��y9�s,�3?��t���]�Þ^�j�V��!#G�^we堿D&R�����؎�t�[�n!)"����0�\21�Vj��BO��Ic��m&PE�&������ތ������.��wb���F���q�kK�:���)�� �� '�Bvy'�x�<���jC���M!{}�N�����F��� �I����NF����i]�o���ű��Q��=턔�)���<��
[���G�]�!�R����1��w�\s3���Q� �}�9y�i0��4r-����KyjlK���d���,�,�L���x��C��L��	�3.t�y�w_]iy�h#�q5w+�=[ɖ�v๭�Om��&�f���ſm�3$�@�<�̲�['��T��WsM�L����%��e����E��[�7>�
�L_A�|xb����1��^���p]�1>�\��P��c�� ���I@cB�����1�����E�JC�Ŧ�^]"� oʌŕ�����N���ϕ�ȉ��M�P[eK�.8�&�p�"�M5�^�:�N@�ܣy
�"��l���i%-0���
�*5�3�{h4ݣ:�#,�ø_�呓��K���;��9#rVDX��y���3�F��3UX�%i��𰡪�`�Z�O��Y{�Jlq ��B�����c|Rg	�n�ײ?�gjY���K�Yִ.a^\5m{��WM�V����O5�Je�Yˁ%�ȉd���o�;H܌!�3��ڢR��S��^� �ޗ/�6R�n����e��G!j(B'�H��]=�ޓ��E��8�vh�zٷe7۔h��#��O���J���-��#M:L������[�i[J��d�5a઱82�7_����/=->W������3�*�й������(��~F���åZ��0{cF�܅?��՘[�xz�j0�F����ۆDyuT�еd��G��r��O��#ؼ9^6�pߙ�6���K-k�v�[���W3AAk�BxV1��<���:C%BF��%�л��2��X��>-����2A��<�d�<����㸜��S� ���;�����=�$.�՗.��A�G��%�Op[�{�M�Ib�Z��� <Ɋj��+v�01T٪nwE�n
�ȱW��7��ѷ>�G$遘���"X�r�ٽ_���@���� g�Y��t�J�{�����i
���t�v3���d��8�aZ�D\�ؽ�JS�{��,�熟7Q �N\gG�XA�fU���~V`��$��͆��?�/�r�P��	�\ 0�Z���G\�P�s7���$����߳mo�8..9Ac=�f��,���Aá
>=U�ÛE��'w�qO�'���@L嶔j&c�(3q�b u���)���p�����%E7��\]3��D7mXgp1@�VT��k$�f|�?3;u�j�p� a	T�I�D��8C��������W�T�=8��r��f�;�+ f��>s�����h3v���K=��c�0
ܲ����w.�Ą+���uZ�U��7�H�2n��eF��"�wvڼ{/5�7:41��èX������}������2r*aGȲ}���ng�}~ԬO���H�Ā�s?���c�ߣ�.T҃�3�C񁤪S4���	������Q���q�F��F�����E������0j����6�������9ui�{xu�����-2�UH����q�:���_�v2��NC�^�}�|4��֤�g<��������{�n����(A�� @��� W"���Cvk]ӎ�Q?�b �3��d�QP�ƴ��D�!��dƑ�}�e���'��.�.*�B�?mT�##%�e��Z�HHF0�x'NI�7�m��\��Y*��@��Џ���i0Ƒӌ�KA������f^4@���Iƻ
j!�Ӈk���1ǹ~��17��i�dK.�*-cG�'哉!��8�t�`��fuP%Ў�.�剭�I��q7�\�fr���=�gW����ZZ̮�*z���@�c�%�E��+\tZ�Ѓs͑�5w���N��G��97Ii˅�O���C���I���3 uP{m��7��+�EK|�]�l�Sf�'���z��4��;sL��Y�O��ai&�g��p��Y���#%Ѷ�\���WR�i1�k�P�:��U!eM���7]$�c��C[x�:�R�ߣ�<��hqބ~B��j�����q�'^ى�����7�5�>�7s�� ��6��urb/5ܳ)���i�muUV�3������ܝ�V �~r��/#̴��J82I�b� Ny�X�
�!Q�����z�볯!�я�G�j�K��65R�Lq���:8$���#a٪m����$Ч����?[���)@���.;%?EGk�~��~iQOE��|����`tc�OC/Hm���·�u�*'��@-m!"�@$!�g�$���Ь��+�<�OR*Kv���H~��v�+.`9T�v�5�tU���o,�Nܪhʔ�UA�&K�M(��m�b������j�l�Vv����e�T���Y�f����⢟E�3���W�����"n�(N��4v�І�Wf0V�G�b߽�^6�éw8PyI�u��L�=r��y�������o��Q\hI���q���r�ɦ~���~H(8lW�6|Y`�
%C�|'���ꋒX��IȃX8rۦ�]�qw:/fY�m��lu��0����[�$��� R�~��S[6�x����L��`\�Ni�w�P��dGs�%����!�rY�ŋ2����8����A���
h��O����2��/1WyM�lx
%���jf�¯�
�$�f�?Zi�Mz��W3������
ӟ>6�!/�/9��9�ce�Uꄕ����d8 ���Ed�r �!&��4��+�)��cˇwY�[ۍf}tR�!������,ͅ�=�т��P��P���?�]XG-~����yU�
|�Tߦ��^��r��s`R1�]��I"%s�������t��Hh����1�����&y�q�7ݘ�&�.����Ɗ�� �)aA2<�@!9�as"P��5�t������о�n~�W�VP%����|�E�4�����nxG"ҊK��]���=��	hҵ�Ln��@:��(�@����,�Q�-E���'0M�$�ė��_��nn�"#�̉4�	Xob���6�K�	N��X��'P�J-����_��\��a���dM��5��3Vk8�lb�n��|��?߯�q��^��`�$���zV��aٰ�a���ڶ�?�̟�Ynv�b~�rEB��a��I��؈'�p�B����Wk`c͎�,��ϥc5 v9�O��A�����$��d,U�\�c�/_<V*�e�=�i�jY���f1�geE�ß�D�M�,*��KjB��l���{���{I	��1�֚5�Nm̓�7q����M8��0���3]�#�<��[�!�")��G�ҳC�|�r�IT��G�7 3
,e�*.B���FR�o�Ӟo(������V�X�<�; ��[��>�� ���d���O�6�E��]/��OX���������d�	P��v, c!)ֲ�wѶ:en=;������X�����h�3C�7��
w�о@|��x�]UYAp��	9�MA@���M��:��ꑞB�(~�;TDDd�e��[T.�����)����#�ȣ(K��|'�xv%�j�0���qs��U�1?1l��_xg� �R��aK~���� �t!�zUmd6�o6��6���DB���ĲR3T�F�"�F>�^��~��H���!� �f�uNb��g����� N�ڶd\��}3i�T>F*ŕ*U��}�y���(��^i�%���e17���$�@���7�2��g|ڵ�i�sZ�����i]��7$J�O�Yi^F�q��R���H��D3g�KT�y�O��֘�FZ�3�x<�#|��QȠ��l�#�&}i�O������K`�j�������KE��6�A�ؐ%YQ�� ��a��Ԅ����]��E��tw
F���������(�ݚ9���J�DvY��W�Z�;6�� 3nџb������xc:����J�I�_�S�;r݆ݔr�P�[�b�ӹ���� ��Bf=r��+����Ш�N*���tW�W�<�E�Ө�9�QT��b	-�a�qf���C�G� >(3}U�����=7���J]������ޕ���f��s�fp�ʓڛ�Ak��j��������5��?��U>��$9�r�ygf��w�\8ҧ�����{��g5�E%JXl�|��K��0Ŗ^z8���r��!)�B�C�DTɒ�>�{�Zi{��T΁�*�rj0�3V� "\� ��Ÿ-T���X��.f��㲻!��0e%��p2�A��X�]�:W������w�E���!U$G2s���|��^�UU�b�$�b�-��8,��_#�O�}�K̷�p^M��/O�9�J��?ߞ�I��1���dW����"�b�c|��+������w�ц4�M/�_B!dh0ߛ��:�˕N>�,�/	�S�;�6�����Ef�hxE�P$����r%R�;�Α%�L����H�==A�k��Nk��n��j���cy�> l{���ʵ׆]1���^�h�Y�Lv	�� iQ��/��3�b�2�u��u��ɠ����J����Q�9ԩ��Ҕ�(3�����5	Q�X����a�ίP�%X�SL��~ �L��)�w�k�A��'��W���iu�8ǳ�'=⌁�:��K8]�4����fm�<�>�8@�R�g6��$� <� �D{l�S5O~՗��m��u�SE��[y :�k�w����G�p쬩Aܺ_}��%�R�sY�<&D�m'�N��f6vDK
/�痌�����pmW��^�}j�@����920 H&��L�)PF�����������xՖ��_�B7��wX�@؟�6�Y����e�_�����Ѡ��o�O݉��:��K�&{�|p��:�z����OÝ,�N;��5r�v��%���WiZ�S$+H�%�ۚ=\4�l�B2u��m tbD+�<aj��kg8i�ˇ�A�T�5c�C ES��ս��b
�c�?�g�J��X'��[���񓮝Q�"�}:�H� ����-e�Fz�ToJ�H��d�H%�1��px�&8Z�E�m���8��*�\d�=;��k�F_��~��T�4|�4�<�8��zя�&�i`F��d�c��Ɵk��=7鲕�+��}�[���-�Z�t>>�u;�a����}Dfc~��w�j7X�pd���1R�;ܜ���>�0��e~2�V�ã��mJQc�~EKCꄈ(��)���D� h���t���u��Z�jg���ҕY`s�#�N�]{N�	�49r�Z�t^��3�ZfJ+@]�`�'��1�( @3�Ųg��;�����>Q�fS�v�a��#ϸ�����G?�mC4�ޙN���œ[��j�ag�#�@�L���	�M.�E�P��Z�z�����'���\5�R�rP i�x�J��il�d�<��MiƳ�'�~e��2phU� f��`4g1��#
�rĥ�^A�\ƻ%,���ҡ���7mސ�E�Gm~�||��E�r)��o��P��������G���3�G e���Q#��Qe.6dԳ�)���NmH��yl�@��YD���z�P�tH!�7OP#(��Qe��N���M��_>H=Z_�g�cU��J�[�@00�5�Mn��]�z{����\%�L{w��nD�����_P�M��� O�05�8M�8� 1�8�����}�,x���M���ӷ���$w����*u9R@�Nev�����2|�ܥ�[,Tg�5�=5'ɖ��t�H�9�̄�@�m�R��{�X��Z��
�m\�N��!(��!:������3��7�NJP���j΢��O��K� }�Hn��5��.�1ف���HL��{��.7-���Ш ���|��a1M�d�㲗�K��s�9Q�rVIb���G��/<��������]�Hx9v��E��X�8��R��,������f�I��q�6fP����/8�o�ʴI��n.c$��\�vӟȿ�ojņ��J�����<�~�^����ʗ�%�mS�n*���{��_���ꆁ�zQ�`�SW�;_k��} 9��ĭ�")h���U3�Q,}枻۩G�)����S��"�G(�UJ�f�J���:��=�̏��G.�w"�?qC߶����vF��O1� m��
#+�.&u�\I�n����ӵ|͋TJ���v�`i� ����/�墝��Edl�i��rr���w��퇚s������ZqI�/�{�r@�j�!$��ʘT*�Ԯ��� �7��Rq��JRRu�a��_;�	���2�,�����@�^�"
���I��b�~��]fjE\g�GU��G�[� y����h��_�T� �B��q�����݊-B�)��BV�S��G!8>�QN�(�̘��q�����t���92�ޜW�N�"6����G���=(�7�	��=2�������{L�ΦT5��e�Fx�s_U	�K�[նO�)���Ժ�}�{�U
�̪�-��Z�Z���5@V��Z^������:G��Cq� �vg�B�ށ��^9m��<I�3�uV�(�ɢ>�4�z����q�m��鎤�>"|\E�_˜���'��;�l�A����8��'�V(��qP]ta݉�pȇd���~%�*���r�%C�z�*`�Jk�
ϒ]v_�y{AO��@}��><t�2nKx���E��Z{�.��������M$#��egš����(���!/����)������C��Vç#l5�c�/�� ��i"e�d&�׾����Ǭ���dA���kǫh���1�P�X��?��p|hż #b�B����s��M����hSZ�˺B׋��Ê7MQH�6<K���F�O�Q �2"nN0|k�Y�
�݉�����8��V�E����r#��\����B�)A@<���� |�_�F6OY�v�f������Cz{�Ks�\��AK6���֑���)+7�8SoL|�aZ��,f[1!U�FÈb�^{�䨤	:���m�óK�V���ț��1��{MW��f�M���\��}ί���X��	�Ӫ�l�vS�5f4��Z��5XRSD$��񦰏HΏ)N�h�#�HT������se�����	����p���,E�;R�d��W0���w��p\v6��L�TU��p��d��
�Fw<	S� ��ƁwÖ�aNw	(��6�hzc�&��"#�K}��6��`�[��׌�va��y2d{O�3� �9�>�#o��ro�4�$j�a'�I.&��fg���U�ո���fM��\8������`��l�	R�t��B��'�[�Җas��F��5�G8��"*9�f�?�Z�ב
5���h�NŔ\��v��C�{y8��OqxI���G�0�\!<�<C�hKa����;�\6�nG�{�N�X�sȇI1����Q�-�.��s�1�sR
u�X���ɷZc�?j��+��Q�oK\9�&��p��<���s=_��0��kҿ�В��4k��<+m|ޱ��T�l-�iD��~Λ��c�h���6�?��y$�ܮ�O�g�Q�?Y�d(֩5Om{T��	�����t䍁MG@t��^Dy��2�52�ݦsqO4$Ǎ}F'��xj���v@�捩�%���*ᙬ䈂��d��|m#r�r�J���*�����ڶņX���'PF@�ϫ�*��7O;C˂s�k���k���׼��,���}:����RTH�(vD{�a'���R�bJQw-l".����X_�'*PY�e�e��h$�46�����	KP�R����*�D7ĺЖZ��ɂ�|�hG�_��ʲ[�<_��{NL��# ��;�7�n.����g�b�B���*p�@T��h�Ҫ�)_��oˡD7*�i������m�>��KF{3�:{�3�p���d�6���UC�޶�K>��M���)+�����#���ڢ��2���o���QFZ?�;qM?�F�� \p��n�	S���@i �<Y�q>�:�Q��j��OphAVT�^Ѫ�}���{��b��tY�u��r�i����JBf�6m�8�h�|@`�>��Y��4(��˴��Lo�](��E�Qx��U냡�)j����U�k{��^�4&7	2C�;`?{�����ߪ�3K��L�,V�_��"Q"<]WV)2$�`�!������{DIƹ+�������1%p�xp�e'��˨��8-��~�����} F���a�-�b�ce`]+0����"�"O�,@O Eػ�#^L9���U��Xd&��Bىe�����;���X&4$�e�q+��r����
 O(>Mh�`h��Kq-Xpثg�8>��PͲ����J���o�+����#w9�K�ļ�&`��r�V�j�Fu�R�n2)`����{�!ĵ�f�o!4������5��r���d�a-�
2�>�e�Ԫ�/=�/ʆ� J}<���[BAƹY^ �"|!�U&"�@���s�;�O�1Zg�ݡ1e��ğ�� ?����L��H��h�����@B�����|���Uu�W�myb�+��@��#���-�Dγ#�@3A?��f xR"]b.A�����Z�U�����ٓz1^��-��ס�T�K�2g�����0z���l���}�2o��JG�|�5튔^v��I��+�D�݉ ���dFt�'!��GI�?�tY~��组>\���2F?h�(� Ȝ_M��>V���̸��	*��:�~3Q�^$ ����4�NI����9�7_��s0�4�w�3�2�G����[\�83�c��`��	�h��'^����I-�;�@5��;/�Q8��5�x�����	z���2�4�U&Њ����>p�K��;`8hn1���V ��e͒7��2�!
�!�HN���K���?F,iC��1�~*q ��_2��L�BS�"��&�%X��B���<�T(�Ţ�W&��E- D%��r�J'�B�D@�7��(���5�_�Tu�,��IΙ��?��4����K^�����/��-�ਞW�Z���g�TT{LA&����	���9c�n���Tc�o���{�-	bpLf�[�ґ6�gD������)ޚ�vT�a'��]�TZ�Ee���ʗ:��_�h/��6S�d�'��Ձ�>,MrnA9z����:��%#yq5>��p�ڧ�S�o�#��}�ڈHxU'd�:(t�o����5#c�j����9�{���C�K8l�:��E$|n���>��q������ޡ<����X	 �2�M`�r����j�+q5��^sKsm�ZG�?)Y�Ȭ�����A��H����X�7!:QukHU�j�9�u'��Ago�����_�0���.t�3��$^��.����L�r:�� u�}9�2��x2T^�,wR�������_bMY���E�z+�EtٶV����۝Iw�Yf�+�Ev	~盾�����:�E�ȸ��Hp���M���
w	��ŷ,!�peF6��"Y^��s0Q6R�!�V�*L|U���xlY5RA�X?�R.z���~�{��-OY��n@�%��n��rN��-
��r����H��2�kU0k:����@�ރ��JkT��@���Ff�rv=]�����Z=�ڣ⸢���7�M/ҏc�"b��%$7T�-�L7�*]�"9h��j�x�:��m��,̓�?��=n��e���h�=c�^G��p_K.�bXZ@��E19����8�:4�/:�C�W9���Up|�F�7)`uq����+��B˴?�S=���`Wܕ	��b V��R-+JzJaT�^l#ޅdn
ލ)s@��?����7����PʺA:�:ݬ��[��FmW	����q�}�X��\4����$C���lֆW�t�GC�ʰ��%N?É�����L£$�٣�"'2���퓑N�X�=���̄-Ɂ�5r��0�n��K_f���D
�ԑ�2�_�8Efs#�
Eנ��E�>������@$t2[����?4�nJ�2�X0��s���͗^]O4�`L�^u.b�½�Ѽ.z��q����o��@�?aS�gg9��"N� n�?6���Ŀ/P[���t��{H�F�	��8ǔ���N�ik�`�*g,���F_b<�����҃@�`zxI$�d���(�!0)�2���)������;�r0U� ��K���K�j 3ʝ|pf�P��R���:S����d�~>AΫ�xF��:�n[%���zs�u�Ƚ3�G�ӆ���.ц�4��H݇�4F�as
g��S Wq0��ړ>(w5��͐�;�X�s�����e�6f���d���� ��Z7$1MM����NY�w�*c�Qbt�^���y�򪛗�e� Nׄ8aL_��M�.O�T7���ASe��qVxV����xt�/��2�H����۽oV�x�������>�5��.L�~���0<)+e����k�u����f?,��U[EΫ������s"��I����=��[
3&+{��/>I���$^>�/�Q뭇�r��tإL���hy��i�3�ݝ��'X/v^�Uws���Sl�ݞ~�c�B��� [���$��TH�����'7F�ׂ-l �7������.��J����@�
gU㌀��3q(}I��?�Ga�*��ߗ_a!E��w�´��B��Ѓ��v�B~5R�b7R�*-�=��HRf3J���uڀE��ӣ����0���!�����N��(�5�`Y�䧋B��vs�>θ�&@r�*;w�oB�Xq��M�3��p�N����t~5'���{�W���C�k-|��.��u~fTNW�qo��d<�9�!x5<~����t���*s�T���� R���g#yB��b�=��t�3�ˈXzՍ�r�lyض�1���L�c�]��	��݃`�~"A�'O����h8�!E*�!��+��ls%�l�
�����2��fĪӤT(;Yr�h1��S�Z�u�-!�JQ��LȾ��\�d~���aD\�9����e]�s���A�ƻ�\�$,�Q=6��f��M���@�i �]�-���f:B���ћWv�y_K{���Y�k��ӑ׮ShJc\ނ\?~�н�T2A�k���!"~�b��q}h�9�H�S����b�f���I�fj��� xF��lb���N7%�b�#"�FP���_��¶���*�� �+��a�7�˺?����U�����
ƾ�:��p� ��Ɖ[����ԙ}ؿ ʲ��^ǆ���� S���g���#/���9�9*���l͍�_07]�8�SQ�� �E	���nm␡	a�4iο�<����z��Ml��S���a�&�8b8�$�:�5 >������&�/�AnǜHB6��Y��r�L���ͤ�N������0��_����U܁C-f��d4����!25�T��r�^A=.e~
�%���j��f	\$�<1�"F��u���{g�!E�E�V�9(�/�֞%�7�ZŹe�\�!]�u�xn�JYQ�������0�h�ο�=���i����6V��+�]�V��u^(��J��f"ܑ��ې�NmU2ih�hLka��zktE��j���*�D颟!���.�4hz�&&K?7��"n /��M1z����V36&�9�A�C�7`ַM
��.}s�!2����6�ɩ�L��ƿ���E��/�XFP:��'<usiZh�l
�x/��ń���H�}���I�t���4�;���(�#�{a	L)@�Աx�?Y*8W2d[�J��9�-���m�m�WY.��bqs��ϒ���������pS �j��'�)�@��'���	.s�~Q�Tz��Vc����5*�+2B�v�*��19�48%I�m[��q9�ɁL2+�4�	AmG����Su�����yK�y#�u�8��YCP�+Hʎ}8��Z��A��y�$�J�,�ܳ�\�|/� H4�++���H��~�u�bL��x+6w��� �(��al�����c�.�����j�ς�w�4Q\��R�5C�����B�Vp�ڿ��$�����L����ZyDz]s�)��]� �]Z�����Zp�u�B��D<@���"��!�!�!͘��!�m'L(�>��ig<c=J,����_�p���0���ա��<�Vۅ��y�|J���0���p�k��Zoa��Y�)���=и�`J�$C.����Vh��H7/�^g��	p���8���n/?-��'F 5\�K�=IC��Z��n�K@U�]R�C���U3>�,��Rk�)X�!�=?���Sa���=uc	�'�uB������e�'�~�[h��ᥥ�9 ݣvu7�v����SH��1nÏ��<�P�ט+�[f?���y6�I֡��J��V�`�M�BifR�������	(�ƾhy#�hGg���UV��|�̱%NSp�1�2Cy0��gRJ7:M��c���h�ȼQK��*��AZ�x4�2d���k�d��Т���������}��Y�`\�E�{!೗�`/P,(���;����Z��A�r�:�F+?VUz���G��g�F����l^7tI�"p�Ө�G�
�T�@F���ћb
�1��P{�gG� @�ba^#�m�fǨ�R�%oXn�%/����Տ������ە�>�ʗ��X��є΢JE�2��a���Ww�I#8��Cvbtػ�C��.���@�l����Z����_P�e�%�]��kE�2�M��W��r)�LE�hɍ�@J�����ى��p��\"NB�X.��?�.�`�ȅC��"!ٿ'N��ux;�
q�4QD�[>��;��v7��V]������H���63��̦�g�A�s]z����	6p�	��b�</�<9'dW�����5�pu8K�n�U�8j�%P4�K���̈5����ex����^i�ҩ�#��rn��%�$����f`z���c�_$@��jŕ�׌U&���������P��tX�$�V�h�7��I�n
v|�A����b��:&��~���=��@��0a��i��
׺�p�:==ka%h;�[c��ړR��Oޫ0%ڈὅ�e*��P���Z?�|���v�w�3k��<��L�YJ�����%�l�*��;2�~F��&i��=V���}��+��Ԥ'�܂�)���/1����&�� C�~?��
��F�HCN�﨔%r\���mP ?vb#���m�d�r����S�µ���MMb�Ֆ������?f|h�t�O���X�3!O�2�D0-���.n�~���|.t�H���uG~��w�>p,4\��W�\�ua�b�x��'w:I��a�T��|��8fY*d�T��9m�И��E��$O�>�r� ��8SӢ� +g"l���8�Zi���*Ҭ��;-��o�""�^��se���3�+L��M��"��'�s��?POB䡝j��;΃�F�����6@��YLm�]�S#��k+N>�oQ���/��Ϣf����R�hIp��� �����0�/�� �ʱ�*k��e;�������^w�Dk��q�>e��Y^i3Q�I�\�U���C�E�|�ۂ�tуn�"+�t�v������[��`Yܚk�^����F���/��g����B��:�x�y�6�H�L���\Ln��FxS��O�| �D����vU�����:����q���N��T����V���n#	����H�/�x����[������'5Ջ�`���{�
e�˶�� �?�|1Z�9r��$d��҂'�WHh�'��<E�v,|��Lj4�S��_[C��vN�|�8�z�5��+!�ꛜ4�c����=r� �W�[��I�'�s	�]�3����/<ɻV�@��cy<����ј�%A��Y<\���Ȕ���,�î�OKEO>�_���M��ɡ} �c-��h4h�{ĵ�D�"�
J�#�>������~2��U���{��
9?܈��¯��-,՝O*V�����+���SC��8�M]��54�ei�7.'3%���$��"1��/�O�^xd��`=��oe����T�˻{6/>��蜋�&
};:o���]p��ʉ���a��X�
�\*��4�_kj�\������G]G+~�#HF�gr��Z����$��-<D���� �<���άa,2�ڙ����W�9%�_���UGu�nUA<$�Bn�	��;=Ҫ\���1!2��{r)Aq]=�W���������Z���Z�-Ye�G�6+7��΋N�c� ځ���89�/����;��ޞ�7k��y^8\��ۮU>5���d˪�fN��su�Sٺ{���X���>��u�&�\�c���8ݓR�> �$�V�'څS��
�b+2EME<��S,�f������x���Sn�N�+�f���0���n�0x���7�ԃ""�gH�٧�tu��J�:ù�ȁ8�FG��n|�͟Kr,�r��d�EϘ6�sߝ䀋O$�r5�ʗ\XF��7�����V�O�w�#����BW�}n���J�R���(����Cٮ4M��7�����&��?�7�� QV�����]URXҴB�~ѣĀ�c��AP���!��t�5(�<1^�t�k�Ć�e�/�W���+"4%L�th�ޔ��HT<mp�Y�w��5���2ԥ��N!34_�oY��8��
��Ku=
L̈́�deU��.��¦�3��`���-cЈ��O�h��,/��3�X���N��y�j���ū�Z=e��3҃��j��Ѥ�- �r �o�<��~hB �7��i�&O�����z�o<s�|���y;UCo˙Ҡ�)���R7�GX̕��k�(c%��.Ǩ���S�l9� ���L ���FS�n���ijG�oa��ݒ\ne�".��2��-�5�����a.H�p�3HԐ��3��*��j�umėf,���)%�5Q͡��H��?ĸnv���m̐�x�.�x�H����a]��< ���{��"��E��>㶓BRg�?M�|�%�[�	�Y��]_��P4���'᪥ ��#8�cS�9�U���*.�~9I��%���� T�'g��؃#��#��	�!m��Z����Z�	@�y����.��<�*ʟ_����|?/ ���4-�V;�Mu�sB���7��t�nr����8]���l�͍ʎ�KI�Lq_��z+}�!�_p��Y�:7�R�9��9�Za*WVkYq�~�7v<��ȱ9E���%k#�ۃ���?�R&�W��y��x3���zɚ���yit(2�)E@9�_%/oO�V�K�AX�a�0I"���b���ʄbu �a*� �uB�����z�ٖv^������.z���?�*W�!	-DǙw�����Ǌ� ���.2F��J�:�����d.�� 6o���z��P�*��
&��-��$;3.5�3O�>��&0Ee�j$Nw90� ��)\hj�K�9�6!��M.�*sJvt҅�!��`�RYFl��U"��
$�sg��궦䕆9��l6��)�?���w#&ՙ=��Baݮ(��Ϋ7�/�sD���A���fX�[0y��W0��9J2��VF]6]�+I�g���4�t� dώʴ�B>g�7��2�&�"�N�Kr��_������g�k��Ϩq���Sݷ?�3�@���`��4��M���.$֜�3>x�:���޵�JԾ��-����F?9�� ��S�2�^u��m<�a���`Rru��"t��O���ʡ.vD���s�1y�,ӾP��n(�{��)-v�d���{x�E3T�4�+kO����wÑ���a�� �H@R�#�����%�
�Fo���O�����:fgc���m�M�Q���ĕ����p3{��;@
�]������к�����})'T0O�k*��Y�2�.�9cL-O�O��W3�e��Uh<3�D��7�k������{|�Բ#.�{K?7W�Lo��,朲�ZE��\x���E�lֹ�5#a7{�~���2�6q`>�f�l(���(#�R����؍h�!��94�iJ^����֡a����3{�nu�H�����=����U趆��W�<Cx�����kq���b΅c�A�jv���B�
H�z�;���.4f<�A�����daL4��|]Po5[¦��Bo2n[ȋ:�b��^���h|��9�Q֛�p��v����m4x|+gͯ���W�Z�p>5Z����6bs�s�`u��'-F	�"�e)��ƍ��;�-k��=U!�X�Z�|�}��R����/Q,��U{׹������y{L��.bʻ��G0�ƨ�}���\�I�uw�b�{~��3�%��{N���©f��?2����y�$5���V�@�]��z$s�TFY��nC��ԛ	�+�Zp�%�3-L�%�v���|-�h0V�]��o�hnĜR(b|(]9A��БI�KI�F:.n�vch�I�f>5\I�؂�Lvą?����L����w���F,��p�ݥRo��6B���+�D=�d�U�"���Ú�t���_�A������t��)P�Y�}�fUo�rp�Gˍ�ML���͏#�J^ʋ���Ee�& ��v�l���_P��-lc ����N�`O�r��w�0;D�eW�5�Ӄ:{.%^��nTR\��RO���ze�m�&��V�6��1"��龎FR<�.3���/�$9a�SCO�1l�e�!�"Xѣ��%W,s����活�o9�?50u dPɞ�����0�{��'4��;�Y�#5~}Y�k��E&9ru��)��J�� ��Aӑ|zCR� ����EbK��
�e��i\��&y��$�Z���CYzr���;�����d��F�B<�0���_X%Ɣ:�G��f�~9�Iض�����z�q��O���tshw{�͟�>��� ��3��o�� ����#Ga6La=v�CW}��G�t��K�zR�1J���j�_{i��>����F��ڂa�?��G2h��������aե�JNs�	��ړ�3~��8�x��1�*���c��¸�e�����YH��k�]���)^��Ȼ�7��F/o�E���g�����*��U���;�4_�E�!�:�c��
���r��
|�]�CE�⑁�z������BLO[ W'�~މ��y�h��둗�w��@U��ܛ����h�^�������Au���@NH���//��(	J��s�H�P|����RkX���:�,�M�0�a[�E,��g�̑ k5�:�<�M��.i�D{�+�j�h�P�S��Ul�4Q��������MP�at^�ǟ�t���[��{�L<J�����(&����v�j
VN?���\PD/Y�W|;�%�=��v=cC-��#��=?`j���~t�t�%��T�`�"V|�s�&�0г��
>���L�7���f(}��-XŶ�M�*�A}Hz�nZ4I�+is!�x��� x��f�@[�g8<T�@�(����(��G�>�Ӊ�+�c��Q��0���P���h��ϭ�G����=�z)��F�c|�#Y��.N�_���{w�ah�Qi��"���!?��\��TL�?�)�����Ŕ�xK��w�GOf0�M�͌�4�5�' �.g�n�F�YdQJ��¡خ��ml!��w+-�<==	�.L5�@�i.�`�rgFT��0�"XxHNq�pґ�o�瘺x�L�����0�����Ʊ�b��}�^�?�F��5�p�����ڮ���Qo���D%���=?����y�X]yioNXoVٓ	dh$����1��bҐ��#V��a�@�[^���i�f׊�e��Q�,�>C#��}V�� SHC�7�]8ˋ�[D*�	^�ZrG��@�T�q]�����f���s��k&�E}0	��w4�B�Ts�K�p�O��̣�(õ��貰N	k���7���$Nm�=8:�"i�'h@C�:����:fa�m��O]$u�!A@��Z��|{��4��I���D]O֭7��\�h8| ҭ���nI	{8t�����Z�]��EE�0T��9b{�&�*^i��"���$����5�l���[�@�x<67�S\�{Q�g�P�B7���6"�L`��m��"u�>&y����7����&�~��9Jo��@��B���I�SU����M��,�(9�>�~̥!�V6R�Q/n����P�x+��B��MzN$~P}_�5���lz�U"Z�	�?q/�������K�Q�H�-���x�"��`�������AB��7���!�L���#�s����u��Wj5kl�'9�l�Eb $˞�����BoC��]��!�h�˶��|��5�;U���HJ��-����_�95��(s�j�g^����bֿ�Z����"�i��_�)}GF�P۶�]�eRz��N��.�-�H���рf'U���q@�Z�L&aT��g���b(�+Z�����4��"eMH��!-}�F��@��sa�$�o]~
�e����??�#À�X�'1�������:oB	�� _����zT(�vA�S�[ ��x�$Zv���5ED8��:EĒ%r�����Վ+F!�n�O���B[5!�+���V���=����ʻ�!��̒%N��^��]���mgKD[�,���4�?Y8��9��!��*��\��Fk�X�mϣ�^H�xrKPK"e�^�ΊK��AӖ���P���g�I%�����B����TL!�r"i��fހ(Ҟ|0��9�B�� �k��]q|���N�IG+d/��Ť�=9�甚��:R��2��x8���'�������ɣ]��j5��)p4o�X�F,���<�~`�^ڎ���?����x;���^��4�7z��oՒvF�!3-v��]��:A�sc�~RK
m�8�7��ṷ{~�����.މr���Y���֥�-gQT�ĩ�p%0�����V42	��l.�]���z�"�6<%憎"��앃K��q�Tt�R��~p�������_u֞�3v00�	8����9<�%����z�}k�W9�9�\\�i	��/��u=�:e��K��o6�.��Oߢ �Xk��6Ј�j�`�t���T*)�i��1:�����r�WQ��-T���x���ex�d+4a]������H*�g"6��E�.�*X��> ��Ã2��E���G	L6��/��1um�/��yP��He�"q!��]0x
����u{�Dt�c�F���C!���@N5�4���4��ga��i��f��K���͚�&��(R�PH���}a10g�H��Z9|f��<Wt�
�l�����%�\��u>/���V���20��+G���a4��7[���d�k����í��
[mOc`����a�sǳEG�4�w@�����ȭ�p�p1"y�=)������(oҼ&(�`$>��B>�D�'2�WqA�c�&C-k��j�J��gKR����(5���3A�a�)��Z����$��GZ���f���9.b_(��8���k3���E�Λ�~��F��;MD8�<#���bɣ�;�B��-&�n2��S<�޺ORro{�8��❪�7���TWsx3?˻k���)���cj�W�q�t��n%��an-��E9=�G�#�L\}$p�hO�i ���s־s��V\z�2�o���m��s�>7q��=�?�.^H�G�B������||��-�!�� cEJ	_f5Q( u�je�NdJ�=�&^���$��/,s�PU��d�4�*������ls� _�Rm���8v�3��чt.���n��o��h��x��F���#�ށ��D���f�<����Xf��G��JFk��3����+��2���6���&C[��x9�PP��sQ��2�8�L����CU@���5m�IX:� Ծ_����@����}Z�$ޱu��N�A��Ng^l�bW:a���h*n������F���=���M�ҐM����ȚD�0��c 7eХ�XR��������6:9?�؁��Ly|7� �]r
I;�r��+����5/C�+3G�9��8���j^NĢ=�u�z�ˣ2�b�#Z�އ��w��$fH�{jd��ͱ�����\*i�k�d-�Xv_�Dy=�N�0�L��n���,���o��u���Z�2�ty�n�U���[�w-���ʩ�Mt�#��o��4�>�o���B�ٟ'����>��	�3x=Q��w����b�sf��Lp8�oq��I)���
}����M�~BᏩ9�!iV��nK��}A�|�,�(��c/�����c�1�k�rszJ��z�����^�����#0��p��{�%��?��6܎;4='S5qX3K�9�֔6r����D���7��io��4q�~&�5�%}7��m
V@W�os�����D��k���+?M�h�r����'��G ��{�	�/�Ǽ�Iw��:�'�x���&7X��I���G��L�}��'��T��5�������������ȺY�zP���9�t��jH�~L&�_�*+Me%`�h�=�L��"y�vҚ���擳�[|�"=���L�������`{}��
�R��VU̍#d�����I76s��"��c��8~ؼQ���;qZxCqI0tHq�g�F}��q�ʹ���P������L���.�4�%>�*2�	 Cr���}7"vo���G��|c%`T�>�%�G���T�l+����E��qǍB1]C	���H�Z���Y P���q7�4�8WzM�c�9�i1�T qp�))����uzճL8��F�j��2.�/E.����2��E�t8�C�H�Dd��зY��"��+�T�IT7d�a �I�`���K�Nn�&N,Q2g�;.J����,���Jx>*oH9�dj�����`Ӛ��`.�W9���޲gG�����=�>�^/�GӘ?q�ì'����)��D0�h�l9'�����Q�򰄼��H��*�p(|��劁��>����g�+��q�x�*A/�\��;$\�QxGk��x�pZ[��>� �"Vʵê	<�%��2Y'�v�N~���.�ECѠ����I#��n�1>�~�f� �]�g�<�UC@����|���|)�׳��<x��}w%�%}e ���3�*�����i�R�K[�#�o&�Zt5�],��r%���i�!�vW C������e<�0N�ل+���K��[�+��s�tK�<���7��e�Q(���|\���i+ �=���!	�uuS�Z�e~���J�H�7su��Df�<�X�e_Wvf�鳾Y4kl���٤�?���Ӯ��>e��ze��Y8��T��C3Hh���q�1�����?�q���c�ǒ�j��ey���������"��yRV{G]L���&g�U����ys�&�fd���u�"׭8G��۠bV�,�_��p�h�3%C�8_�k�}Y��
1�l�-֍r���c|��Š/X�z�L#��,ǿ�}��0�����:>�E��H�R����:S��wɘ&ly�)��U�R'��2��"U<���Xms��#��(��\���m�'�}
xr�%�����7�X��� K�P�-�hpO̯�GW�4;#�s&�{�6 �Ѧ^l�O�􆐡��C}m*й��~�nj{�I_��s¼�]kF%��L��÷��:�&߻��D�ƿ��M	�W�_���A�4�����Yܳ�D�?�:�&kS�l�G�t׏
�h��s+%�:%������o�����P��8����V�'^���}�!����M��& �<A����҇�^���&c�-�E�m�"kh�4t!����� �t4/����V��&{+} �@]"�,q�+L���KM�
PF&�zL�(��-w�SdǺq,HYfC_c�e�����E_�A�#Z_l>bv�ǉ5�0�}���)�bީ\�^1?��a�s?��(�;?�Ƴq�E�,&+5�<��a<���wrV�t6L��3����I�|`�E��x����$�2ǽ�r
O���gɍ$�.7��TEJbv�P�.�g�ƦV�!re:C�A�m���� MC�G��{y���u��aϫw�fX��$��@��\.D¦���3jr<�b§]54��ʀu�v�AVpz5��k��2K�#���*���׍)���0�lj}�J�'2��C�\�-�^�ML�aM�ܩ�=����k>õ��3:��GЩ}�5��LF�\�<k���f��k�k;�;����M�
X��8?�xp	��l��"����a:�E�-Կ��30��8w�B��.wQL�3���E�M�RqM�o�3�A�%]_��������$�����V��j"p�6�0=�*�f�vk)�ǐ���pn�$���Ly|��16v�C&w�\,�!���%���d� Z�=6.��?�f��Ɛ%O���-��]K���1OCi������F��7��K����5�
���o��ݲY 4��B}��Gj\F�N�+Tm��J��CG%10	?�.j�7�K^J}���<i!J�ND0��D�5��l�8�R�����Y�,���J�'�0F�D���(�r�B�����'!�ƙ)���ө�}��T?�5|�O.�=�pgqT_8aXn�.Dc$N�+���"f ����������"`-YEf�n�Ѧ��koD�ok� ��LU���LU�C������kXԚ����;�g��d�\��C��2=>��.(*�>�u�!Ø�����ۗ���4�y��_͉g�lU�y�hZ��V�	��Y⦤��F��Ծ�݌Se{i!t?I����@�`/�a��@rW���+朅� ����Rz&���B�P�D�ٞ �S&0d�jU{r�q�~�}06�����hTO�/Ǆ�d�ov�2u�_\���
+[Y��j_W;v�vI�Tq��]~�8c�c7�B���C8U�*��V6�l���c�f�u#��ײn(p
�V��L��rx�hǼ�=Z��.X޷��j鉸���:�J�>��2����X7o3�b&���$�-�õ(/�s�*�E�_z8f
c褂�1�l�ӛ�bK.zH�����\=g�������J����ʭw�/���My��N���^Wój����kf�S#���|;�3����YN �X�*4�tHRR�GQ�k���ө�ܓV��_����˞��UT.��gI 븞'P��+f�t���:b���3���o�x�|m[޳��(}��l�8J8�!&n��<J�7|k+��^=������f '��8H�C�������N��1���`N���*�1&ʜtg�J�v}Tp.�`�i���+�,�6�uzC�����!���w�T���{X�U:�v�u��Y�lĉ��:Ѽ��(�Z�<�>�ו��*O�<M��b�@Wcj��n���ٹ���М����o���n�e?37<�b�$b�߁f�,K�4�� �3��R��
c�L>�<�@�`S�#�����SQt	������->]эEn�H*�tN�wN�gk��(��OFg��Wm��&�K�G-������3�m��G��v�w��D���ɽ�n߹�����Un28�*��!GۃU����H]�؍+zN%<��$�g�.�.��i���u����=?(8'�l��8�d�����l��j��mْ%���n��?J��}�l|X�i�,��J�.��Pa�������a�uy�j2܈�X-�_��͌
b]b8V������2�Ɂ$����Hi�����>�*��t�c�SjLb��8�cƤc��?�h#��C <d�ߘ�)k�WZ%��l��9�3���kDդfb�W����>���1�pn���~�ߏo��I��s��<��m5ϒr�"��ī�˳
ͣ��.��IM�b���j��[<�H��є!
PPّ�ߏJ���f�Rl��P�[dl�٤ˣ��?(�t-%�W]r��n��vN�C'X���"m����6�ӝ3�|vѶ�m��#�b�h�`:��/��"������	1(�aH&WF�h�t{�z�.Ol'��h0x���I��0���� �R�-4� �c<<�
+�LІK�+���I��#Űm�e�Op
🎝��U|���Ǡ�5J��>��2���*������9����p���0$�]	�^���o�˅QG���kElw|�' ���.�Y���b�ͩ�NN[��(�7g���vVs�o4XT���4>!!ʓ�=xE��6Z��$�_���j���?�>x�#��J0�z1Ɂ� iG��l9I>�\����T�@XU�X�廋M2S ��. ΚRa�`����q*���;��z"�Hl<�'ڹ��xS۽��%�0�wߦ�h 0�Q�(��VT�	��z�BA��1)���̞���r�ipWE���q��5�E�#:A��i�z���;N�z��u�+Zn6Z�}x2lv+nJ/��0i?#���\�Ů�v,� 7=��tl*jIz>�n�5b�ƻ5�ȑ��Eγ7xZ��@a�;�m�#G10�1��l��^���I5`� ���t�g��@�J�߳!����4'����tx�|4g@m1�{=qEd�6�y�uf<Ws��0]�ҶZ�$�p������NS� �g�����|u��ٜ5?%��7:�}屆�m���� �~�4#��T���y�{b�6����49!����^�e�dQ�(��Xі� +����v�6��Z�a�Ï|[ ��q����m��ll*
�u�Zm�y�SV�
�\Jް�AdS�:)�~͖C�ޔ��(y���]['��{�Hۖ�l��/���"?F�E�=��[<��EXe�B�}<�4��¸H}��G���:�������*�e<l���/Jj�������������(td���V��
㺡�딺%��e�y�1�1�@�{Z����&�	��v�jO@�st��&���a�� �Qx�M]u���k,�S. ��D�Zº��� A�����Duk��UA�(�!���v�ZZ9ҍ���١Ң�`tu�����pBo�X:�ҝ5 ~?:������(l����h^���!	ՙ.���{������b�嗗H�9)1���SB�n�R@�w��n��0xNk'~"-OL�ݚ;�a�(�MJ�\F$��RO:+�ט�t�\T=�����
t~�W~
�s/�� 82����Q�=n���C��6"][_�?�F�_�7�{�T�٘Ib��"�b��۾_11�i�y�����G�W�tF���}K�8�A���������l�5��#����&M��j�*i��6}���E�?^j H�t�ǐXI���!���e�{�e ������l��e��6�_LuM���p�1�i�O�;����	���>�b�~�Nh�u�Jg�L���+��*�
X�K��s6w0 ���F�A�e˫�7Oǝ�}�BI�QY��@���!�ɽa�p��6K�{�}���N�xO�K��\�k,�C���Z��{�@O&}D�a'�8�I���!���j !~�<:@H��2VF%!O��[}k䥋c'3�F��̯�&�u�_��3��nT,Vyk��XV�����:42��Q,�]	���0�r݀N0�6��z~r�uv�ĕ�N�� ��c��4�MǢ%��=c��S�u��Zm�[�B�gja�}ЏI��)IZ�s���3��Z�^�>�ƣ˰˔��
���s��N���,�P<�1��4� �u)�?�T�"{�҃��0��f��5�϶̤����e���E��lt�[)���_�x�zT�SA=��	�$%1MK0����g�s�5�i����b~V�������J-�Rd�f��$T���r��Y��βxnE�^�R·�9qÎ���;��*�#B�u�sp�|:2��K/s�郴�6�ޥ�3J�B�u,���(�Ph~R
��mXw�_F�(�X�4%΋��2��30&_��f�G<w�MΠ�4'�$e���ɯ�o]�ʤz���N�
���7c���x&���� @��I����꒳2��^��1������9��>-��}������R���6-���bÀ�}rA� �s >+gocD��8���ېђl�TX���@�\����z8�Eט��Z�c�>)�^k.8-�}��O\T�Iv�魰��)s�#��ꦸZ�'V����qL?/Q���@_ގ����M�,r���]��������t�f[M���Fy���u6�S�x"���û")%[h}I`u)��H��w���!�[�u$
��w�H�ۈbvG���\=��U��溗�}`�-�:.5UJ	Gi��d��)�Jԋ��qMs��j�ܢ8^j�6�H2�����~��R���-lpxYB [��~�����T��5\�̓��Wz�& �3�i?;�~#���D����#�u��ȕ�ܩr�T��&�?�*��9*�V��g�ڐ�*{)��_q�z�T�J,o�ϑPx�bD�w+��'�\?�w�j��Hwe�QB���nM�L���$3	�
���q�K���>4�_p`��8yk�-��zf�xv�	 B֗�o�?lp��ڞ*-�o��Z�J8"�-��
��coP&�������Y�NY��{/[���0�R	S ���)�HL��eg/�l^�0�1����C�^	�2̊�yk��"!�����3tfEDad���e�Z��K> ��n�}��x��q�N5�:T���c��j��y��������o��$�ل��r��agnQ}d}����9ԭ����QXt�Y��rĎP�_*���G����#�|=�J�|�?��R�Yŧ�۰�nN�d�"�&��e6o��P�)�z�����ñ]+i�ft�7� ����z������dݴ}�����'�ӐF�$�f�1*z��c��d���#<b*�ٷԝz�o��Mx6k�yHΕ�0��9�t]�����ݙf�u��0י���cNK}�jM>�$�}� +�vq&zu���D):P�p1�m�1==,ͤ�e4
/l@�����I��w��ߟ�M��'^v�<�_��NP-#���.�bqTLT��eA�Lc�1 �1O"WO;c�OhV�s�>7���b�<�"�g�����a�*Y���)^�\�ʋ��5�/ɾ��e<�yLL��޹���{I�:;E��|�N��l����/���̋�ɖdf���+� ����&��Ƴ�.u��e�����Y�ez�kiE�l7Ez��*10��@�,ŀ��'��Y��~�I� M�`]m������&t ���Wa�������8���p%G�6p3  Q�"��ɤo\���ѱ-̤���8�i���>ar�����ޣ��6���o7��5�y0�@��	Q��dȱ�GZ��Ơ�\�8���\ �j9�`ے�sn_Ax�X�gڇq�Sa��g&7rZ�5J���Ӷj��g��t>^� ���D�.n.`� T���ղ�([� ��K�sƔG0g�P	!7�^�&�Ǉ7b@�ZQ lފ4Q�K����:��21���Mf��� �iq��*��_�P9���ʿV�g�3��U �z4EFh�q�r]�{qKV�ɐ�R�Y/�;G.7�T��߻�$�|�d1!�jAq�#w��lY{��T��W�	.�̣����S�ՁB����
�R�C�It��P�G�-nj#>�F��pAL����*8_�	��:Q�p��ıx&��bc?�y�������y?�fk�τ�Q���Q��!����O��R�N�şߝ<0[�b}ѧM���|B��i	����D+�k�(���z4bl*��^�����=�\$
03��X� Gf��f�@u�վ�m��5��/h*�5ϝdv�MF`���N���j�RM/l�e��VSː�F��v?5w ΝM�XjC"g�S��H\"Z�R��}��"�mZ�O.�+YEs����9�#)4�2���5#|_X���"ꕘݝ�����٪��{��w�ڷ��It�+��j�?���͟�4����x�[���5{y�v�H!g��ϖ��1;����W�¸�_-0���n8��텭<]�T��<vφ�;��i���e���^.��m�-�D���ط�Z��J�Wk�Y�����M���d����%��'���0dM����ݢC�ɡ������!A�/VS;�Ʋ
�!:�,^�-GԵ׾[%.��:j,K+�ò�b�2�1x���c{\����FE� �h�sk���)'N��A���=q5m;��5p�Ռ��J�"9��� Ixu���%�NX�ڬ�i8��[:�_Z�
):��kdw] M4j��X���A���L�0�Ph��<��4B��n��l�Z�'m�h���c�r�6����\��T�e����+�#ZF�4��S��l�UW����H3���$�#���f�^��^�. Q&��!8#�$/KW.\��E,���8��]�̄ui<7v����i���6���Ú�-�����%�r�"�\*.�D�M���F\�"���2f���#�:%�W�}?�����`)tYM3��C+�V���Cw{��p��<LV ��{Ys�=018_N���=��(78+=����Զ�� /�C[����x���V��µ�9�7.ߨ?�6���['l��l[�G�T��Y��V�GN���W�1��a	�|��Ӧ�>��#:7��\�bوF��M���Wp�Zʕ�Y��%(٧l���i�¥�
���Cy�0�phc؛j|X'�4)|Y�Y�Y��S�&�!<i�t�ʧ3v-5����YJ�����t��+�6�6��Mf{������B���q�t_��Wv�W+�����"*��7����r-�a̍�60���u*�~���c�8��9��ė�� =
���ps �g�g2��<���6����WL5�&-��˻��E|ڴ*���v�)��,�<%�h�L�`x�=J���Њ���oQ��`�D�}��HuJ~l��r3N.{�3��c�)�:ˏǐΎ��k/�R�b�uRS\*��V%� ��_��Ԝ�4���K�l��v,�����W�i�[-4�fK����E�HyY���HaN��	U���D�y� (�����AR3�d������b(�/yR��u�� zO���u(ٻ�)xu����I����A�$dK	9������	/ON6<���4��ے|��j
��a ���!�F��-�ъ���̣f�������_���U�X��9��͌(�:Hk�T��h��/�ڎ�8��pKߐ+$�#a*��ě�Ed�l��ieeS,s怓+��g�J��n9-u���o&�TOt�z�A����TaX��+I1���Of��i$�e%��,��|nL���x��l7x:C�Pb�p\1,%�����?L��j0���d9����s�z�vg�_k�=1�Gf��stU֒U�����T���U����UiB�Ɵe@8��ɯ�N\1���*P�DfT��R��w/j��M���aHyw�}�uVd+Z_�q�&iJ �__���6�U��an�T�u4���E>';T�J�G�ְlW�xC��e���U��fiJ���$U��c2G����D[��aR|	uы��b���#��$���&~VFݷ�7���E�<��#!��B�{�|* ��CJT�"Q�NZ� �=�!c��{���q����vf�w�R$m���I�'5Ӗ?L�/	B�����Z����ȝ5I�3���ĭ�1f���l-��<���%���{/B����W�����-��"��RT���i�;�'�~O{�Uƌ<V,�70�J�ȼ1���`�k�4�+�x2(0�R�������O(��ׇ�������+�Wh�U=�g�����
&��#"_)�c�l���\����EO�nO�GC��*��4H���Z�_BE��bM���qG`R��a��r�n1]s�#^js��F;��P��|��#�w2r癑��-\1��Js�����,�.��\b��$1љT�=�L����@�+�̨oU�r��]�yj�*ܦ�$��=�R�j7/|} �aV~�(B������!��U�����0ɲ��l�0�O��Zi��ňͮ D�/:�|UL�#x\�~
&QF+�"�g3��Ϻ���@���h��Ţ��Z���?9��)�f6��^r5�#��PY��MK*3d�:��w`�'�����j`�pLa���ƅ��\�&��� ��ϟi�~ⷃA>�}�G]������g�8��G�Ir��i�t��VR��lR�#�)SW3ht����	4&�Г��tV#k'J3����<�r5}V��'�Z��i��oxnG��9 -^��X���$�#AR/�P� �XH@N�$�ԏ�bHq�hj
�jdwU���{|�vq�~KN��D�4ztj��Τ8Dii�Y�AnR�z=�y�϶�JtU��ű�^���HJ2��mF��֦�����E�A�6|�ހ��/.�Balir�ܩ���$��Dǐ� ��V��2{Ͷ�Ae}�TU���&#���ޫ1��0�������@�H\ʷ��]W#ଡ଼�;��-�z]&k�w^ډk�_�N8�ĥj��B�_rT��y�ZU+zM��5�|��~�G^���E�Ϡ�Z�s�@�q��Jci)��?$�c��s��t���nD>?�Q�^q�چ�F��?C�C@Hw�H���#@�P�aZ�p>x���<���_�[k�,+܁>�!^@-�FCi��U(g-;�h\g���>O7<�V��u�u�DF��r�#�\O6��1��&�L��T��s:!;�ay�ns�����X�ˣ�N���*RP�,l5j8��z7=A��.|�'�2?�P�&!�C���_g�NcI��S�
O�g�~!���4@�������{L����	D�!_��++�`{�-p]n�O��T�ޅp�R�J���pz��'�S�'�p�^�8�!j�[hB�03�%PG�].��|Kb�'���7�������x6%�^�s������5
*k:�(t'B5&fhϷ���N�#�:��XA�)�8�`������`���*�X���0�> 6pȎ�.�+yd��j�����8�g�ӫ�utu��8�h(=���b*+�Ŀ�rh�-vz�VH�U�V���o�	���\�!������&���j��#��V��(�L������j�V E�^f�wN���SQ�[}yݎ�`~��A�֪�Wg]�	U��h��\U��Gm�_� ��܌�	�P���4��[/�X��RЌ��UȘ{�H^ W��
����&]
k�C�3hȳ�sP[lf��a�b&o-�,��o$cV�f���K�O�е��c�^ɰC�R�%y�<�͈ŉ��pt��������~�T�l�8�V�\r�P�@��+�܅����Q��k߻��:�X~��{����Z�r�&�Ê�P��(�Ób0�@�H���}�y�.�_3i�ʆ@�j����@0�/?&��f��6d�@)���DkltFC�;�b��q,SG�譽��"����R�Y��T�T8b���a ���e'��㥏���cR��0+]y����!����P��?`�&W�s������u�_4�w�]V��e�c��j@
Q~h>��3N±��p�L'S|�3E�-B���e(1��1�ׅ	����L]�0��S8�!7>����Ie�?�Mlu	�߆$�t���)�,�ɉ+/�Z�h���Р�l�����re??��~��<v��:��W�) ��. �rZ+M��� k���X��u��l���GK�oO��ʣ,o9
�\d�ݨt���DtjL[��u|�d�� M��&���=s�]j?��@�}Ƭ��f��w�.@�f����N�6�_A����e^$0{�Pw��Vh�usq���VBQ��In�b�ʵl�x�G�с���\Q�����F�X��Fxр�ЊH{����S�Ed-�<Vi���Z�B�{�����87��}���ѿ���nꡄs��%�p�4{N��G�������5acцs{Vv��+�V O�S�J��F����D͛�W|����m��K�}�	y�<�
81�b����� 	�[馰�y�;I��1��4N�� ��86o�{�Q����������]�#b�p/p�?I������i���S�ۙH�}��h=P���ҫ�/�]l��>�7w�
�0��m�K�ɶ��k!(5&��n�ddj��i��M��;>���ሣ��'X</�4�3P<�X����q��,�w)k��W^��Q�gBZt��e��(0{I`�C��t0���Z{�IY�Z"+��^�e��w�u����g|�PN�3x�kni���8��3Y�fZb�-׾����9;��
���3�"`�a-�P^�6-��T���fq�v�O�^k:9�VRhz��<3@&~w��cW�_��^6���&,�r�UU�����O�1�
�>�jM	����6���K@�60Y��å~"Y��� 2��g�*~��ɋKߩ�9X]��N-�;{���r����H�K��ἥ��C�k�\�`>��S��x¹�;���xp�ߋ�g�H�K�����5�T����5��`�h��̅��6
D��y�����9�O/bQ��/�8Ql�����D�u�4bg/�21\�cB��m�c�  \�'��vh��GV�O���@�b�~����"��(���oP�]������24�0��"�ʁ�ԥ����L�ލ��� �N�ϟ	V-�mp��D��7��g_��s�
,�?�$�F�Sm�M��4�ғ��CO�� �\G����X�ީ���\��6�cǻX�ݰ��K=t�@���[B��.M��4l�?&�����4��"?���og�,�{s&λ�5���x���&���g$��.�eDb����%B�h%zۻ`c!�7YΌ�̻�9���s���};��^���:6J��vx�H�a�o�>�7�TtUg�����kR&v���4}x_�V�'Ro&PZ��:���VU�2;7IHAx3u��������ޝ.+]L��*/u6��H
�"��M*z�|���j���t���K��CWUs���U����G��׆0�Soa��^Ǒ���G�0��8;j0��u_�Xg����=���0���no���%���DE�}�&ݙ���Q��O������MJ
��b���-ғ7U���ˏ��Ԓkg����3S\���4.c���!��q�����@�>�Q�$�?:$�?j9����2�X��B��j��U�R*�������s�����;
�O��d�T�I;��u��4�1�i���n5��8�+���`��H�N�����$,`�;gY3*N��fN��0F�M�`8P~S;\��[���D��~;4�[i[�`Д�8��_ RB���Kόodܗ�1��5a�۽�{ogVF.��jf�Tw�X|a�Eɇ�	0N��Q���}�ŰN�"Gu[�mz	��C'�׺0^/iި'�:��DR���к��c",�
�wj�|-<���[ �Sg�������
f{_Y��\�Y�	
��z����S#�|v�t^��k�K.`�N~�C'J��H��� B����P�[^���(,rҭ	d��U0Duix}AY.�T��{k��:o>Z�ć��K�eɖh	�b��_ZC0���X9Jƻ�!]'�A��� U�62��N�����s��e��� �U�]��&���fA���!�m�xe�Ȕٌv�L>���y�.Z<.�����-��_k�,�F8;�eˌ,�؇��j�x6"���Jۊ1Fn^Gn�� e�Ⱥc�_-=P~ٕ����z�Lgn���(�m�oe��������l�w{�iSV抎��ņT�Tpk`�7İ@��6X�/D4UVS	�xd�'��U|l�*F���gF�N��C5����~��d,4�*�QL�h`E�l5�u��-�A�@n�Q߱rh,f1zwvq>�Hs�M��S�U�����x��%
�0Y�~�����ct˅�D�q�\�iN&J5�lz���M��l�)�H�՝&w�����3�Z��=�)R�n�B ���&
���#JT��z<~�0qLY�Q9Ϧv�k"�P<HXB��M7&��B$������;��x8Pn��L���'�G�r���C��𲏑��3�e�����3���Y}f�$u�)6��TZ�$�o^��YѾ�o�spo���?m9xu�E���6@bohS�V�0����Sm϶�"� ���P��d8�p��<1^T��2U����6�|-����[^4��^݉�bz��y)�>w��ah�S����W�1R�ϴ�&� 	�M*di�Ҋ��$!*.�:�_���p*���������3�e�;������vP��w��7���bA���p�j&ǰSO����K�� 1̊�;8�u�qRU��6��a�M�_�9P��0�q�����y���(Q>���F��5���K_��s�U`R���:�N���	�l�������&Ѻ�cP��% �������E��{�KLq��_�|�[q�����턐�D��/tҿo��,I��y:��������QŬ�~�&�Q,C�!�q^�&�a6������������(!)P�?.�^Y���V����z�>>p���ϑ<�}��+�{0�~n����~�@�(�Gh��~&��4�K�P�8�B�4T�I�����2j��h�۵`�H\�,�[���3��� b�A���$z�#�vsO�7� �8�]uW�������YKB��?��V1��l!��'۟�})���R��u�uV�U�]�<���!r�đf�,`j��tO!�qC�K�j �.��S��͢;�02��y�Z9��Y�w0���@�
I�òG�2-��	i�ڮ��S��;��w�ə��Ξ�&�#��ԃ��Kz�X����76P�爭%�c��������/L+C�#*�0�]�`�$�}���k���2B�|��ƥ�f�u���gM����}s��>��ЫD`^���8&�9�JE��C$�W����d���ʪ{Т��k�vg�O���~b���\�M����@l�1H�P��dU�t�[A,�Q<�%�0>�W�j	�BQAZ�x��;H�ߎ�!-W�>4���#�ĬaT<	�yK���zB�%�}���Z"}-y��rN���[BҮKf��P�^̘+àt�X��-�!�B��n��0S
��N�3����E��(��?_�)�{6���i���>�W����D�ɬ��D��mc��fd��AS�z8a���n������dTᅿ+�������$�G �N�Es2��Q"�<;�;i`'>r���j�*ۢ��!Ro=��X��_�b]�@;Sp��T�����U`���Q��I��uM�L�9�0A;=�9W3���O;�*�����k*�EB�	��l8i����i�B��Qsx~�e��{��D�Cx��3 Z`��ݸ���2}�׺]~��V'�����Ka�KK�_C������
m?�b G�u��Hu�FL`��ŝ*=�A3���v��fhV� ��uaj�U;�H���ԧD�a�@��$��u�'��7ɽ��/P���V`�-�B�Ne�=N�Ec�椑F����l�w�R�
��*�-��i!��Ŧ_����4�>�>��[ݩ�u���Ƃь@1��bE��Y$�7y�;B��KHɄ���fR/��,�~=�YE�7p�GQIYne�u�P�|^]��V�
�������?;�%���C��vn�K1PdL���E�^����?���/K��&��@�	^�ES������5��x����4��� �f��#	����j���K�@"�~���s� �vD!�-�kS��U_��?.;�&	�K�X�d�j-r3�\��]U͗Uam޹�`��~.�����Z��:��	��7r���	�>���}w�;��i/�_��-0�yo)���.�q/�s���-r��p����<gu:9�c�G�����Q�Wo��������=���2@����p���J��~;7�Y�K�Zyܙ�Y\QB����݇&]\;���)SZ]d$v�V츾�}ȟ�bf8x(qScu�Q�?A���K��?]�Mr�Cz�������%�k�gBL�l��9�E�����)r=����/A@ct������)۲�4� �O0
�oQ�~��O��e�畛w��x]��/��MQ�?G+��r��5�i��3���h6.�,-A@֓Ak��|�+��1�x���գ�D*�gᾱ�����Fmp|�dН����Ej�W��Q
B�TC�?T�aA����XGEoM��Ifo��.|z,+8��N�D�w�b ���H\>\ �Yp#`@kC�V�{#�B��y�fY,:����b������͆�B��kR#}rK6yQA�_�Oz��Iѷ�Y���Բ�E:p��c���wf�@�����NW�����!0w&�y��_D�%(�F�*�$�6i)�3 ��R.P��	��+NގT�,]*+�%��6.@	���&l�4q�bcBeX�g�����_2e�O� �t�y�RZh�i�6�zu��=����owo�C w~:hg*��3�`��kg�z�p�:Ⱥ-��LT���/@�X���Bs�m���`Ϥ����
�P���i�l[0,Zlv��C�,����'k��y����}�<V�7���$<'�羴����~KX�;��3H���M,!��������T�(`�}ڨ̂w�����2�w����I��F������p�a�_�ۿ���a3X� �ʢ��D�*t��J��%��g�1��P*u����� ���I�(f��!&S62�m]Sh�����ɧ+
S\z¤�1̓zfJ��u��_�PO1��UҨ���*Uȉ�x�`/���/��js��lT��8��7�����q(��&z���	��]�d�:.v�q�;����uM�K[G6�Bv�%3�)���.c��-|��Q��<���VggMQJ�T�_�}?�V���ݠ:���K%\��9H,�!p�.A�=�w"*�s�G9H�<DuB���A:3���׾W���0"�E��.��)U�TF��^.�U� !C�2���'�}Li����h̏��s���Ց����^��^�z��0�3�(�Y^d�8ږ��Rm�2�D:2w%�~'�>���篒H�}]r���,���~�3P��V�bB�s�ׯ�z��~��Êr�wc����z��Mt��)�(~�<`��2-jA6�٢��j㫈���f��!�l"�5�1H��YoU�0'l�	p�J���XH�"�@���ťک[���z��A��e�����ᜂ�p�ڬ��$m>�n��$9��œg���k��i��^Ce�p��_��8euU���Au(fqOw�����]=�#�6�$
���є��H���x�N�.�\�a�F����9ա��D ���8��y��J)��dd�iيf��@�W1l�Z��!�l��?q����9�$RbR��%�^P�F�/�e��O�ι��"��-�um�-y����@���p.��u� �s=o��m��G#<���a�f�|�P����x����R־7���<g��
Qh�y�����!vw^�Oq���<D���Eh�:���*���2�t�'��)���U�2�<��lʖ�>2IUe	���MK6�Xe�pܻd׷�$	j��V��w��!G�CW�P�]8$��p_	�� �%��C���ʽ�Hym���2��e��OS������f`; #dz���,
��5<~��̷)�`j	`��A��R~[P��$�A��7�5�^ȥAuxX;�A1hvW,�bw���fhL�/c��B�k�]NG��+6�A7��0~2Q�-��F�%<|� ��y8�F�l ��}��Z3�s��<�̵�������;)�Z���*f�U��H�O�}�t�����Ix�T/\IR�k�����}�/��Pc���ڐ14+4	ź$�H��Ua�?'���WW`���fEƲRU�[vh������jxz[&��nS8�t�����v��B�̅r�߷u�ԡҰ�{ $1��/�y����SO�hu,dcd�$��"�\d��X�LR���O�}�2�/��2��9O�����61c>Wi���v����fu�M�tޥf�tޏ�6��oa����B����d��s~Y0L�@�v����U~Y�_Ul}��$����©�ф�DY�q�On�V�X���gU���Ш�����.�����,�/$����GIng[�d�Ԇ�:9�9=5���|e�(qdq�5���5��l9�t#�����$�V�#���kN}"��M7~4)�	��.�v+�
2!�z!{����\*�:0����Uv�6NJ;F?�nn[�>wcS-͘0�t��\6t��4��M�]���Mt�& ы]BG� ���e#�_�A/��$�l09@�J��/8H�"��f�L���ϴ���a�R�3���AN��W9}�2��1IX�S�?��s�Uǁ���w�,H���1����0.{�����*ns���!��Y�\����ez6�?'%�Ȭ� ��H~��9�҃�kgv-,>�c��4>;s������� �����Ziob"F 5C��"	��o�6��D騅�xH�����?�Q�ڃĄ�������?j��<�L0a_��g����)�Z�?��Q��>|�jk�o?;�� �b�����K����tL^��p��R�n8�և�T<���iҺ�t����7,;ムg�,f?W=�1�E��f"??2$��ٶ�8C)l����]%���`]�R�v��ZD��J����,&o�oQnh���FZ،��@��(	��P��M�pō���SÂ$Y�s��1Q����K$z�Mc�o�4;=���>���qr�K��Qm����1u{�������ܖ��o�(�&^��l���R*�%	�(�r�*� P�gR��7{�y�]R������HX�
���wь'8���_`u�ψ���#�{�u"?[}�r>ˁ�p�ӜO]T�~��nn-���0˒���5�} �(�����S^\�׏��}-Xp�M���{}IK�4+>���7R��m�׽=U�P}xt_)�Z�W���b W��2\2�^�#m4�6�/����R��&���;�-���R��KR7���M�$i┚iq��)�:�W�PX�|Zq5(Ƙ�`^�}gcw9�J�X�d*q�K�&�\yA����RP%�rUr&���؄��'j	�Xn� o�Z����U�_j[Sн���d��&�g+��^�Kw������1��b(��a�yơ�wF��L�o��3��q~�05pV��V���P�ʆ��6��z(�@9�g�~�!�o#G����4� P� �3G��:+���u����T�b�zk�xg@��*4��y?���g���
bV� ��_��ޞ��"�`�X��ҽ?
ʕ����ˬ:�J=\@"�+R��'�W�pP����������}g�NwD��B���L�����C+y�M`�w����� �W�]٢�;_��A�o�.z����o.@x-��`��7��okd��a���0&D�C��v��dw���ν����K��	1M�/�+4� v��0���n$����������<\+�tN�Z�c���G�����
�G�~�����<3��$���J��F# iHq��C�� @�j��ݼlo���Y,	��I�>۽�L��\�4u�I�/�t���O��L��7]��{���xUB|Ԝ���/
]k�1�?��%�4z�E��N�ldY�J�1Ѫ�������_�1%#J)d˹0��,"����X�?��#ˀs�7�L؉�7v�8��5g2���	P��Ux�/�����ж�~sM��, ��G�bm ��������,8��ѯ�j�A���bዜ^�; �a�ˡ��z�Xѻz�?�ÃͶR��˽������������ͻ���ÎhŞP�)�_1�h.���d�[��D��a��:8�|mu�����UL�`�#.ٺ���ֺ�Z5+����Tm,�Sd1���u�()��+Te����?sS��X\ݎ��xV33�Z��ϥ��*7�;������%���: �յq�8u(�;zw6?��� �B�1��/�aZ�G��AqLQ�'^�\$j��S���g��2�If��M�{K"T���~�46���rv��ΡF(7v��mȬ�b,T���aӣ�+�$!Za	w?j#�@��C���g(k��}�Fgߛ�̒x\��"F炆��TD�v`��m�l;!�?�)�g^rќw�Wķg������m��V�u�����b��4=���_���C1x`�~Z��߅�ẃN�M*P��n};p܌����z�ːֺ���d�5�7m�19P�ڏ�΅Id3a�r���^`�K���M���"3酪z��(ʾp�v��)����!.��P�=�6�v@����2�w	�έ���̰����5�B�MPrs������Z{��=��C]�;�m����Y�d.$~+�Fc�3��T�]y�!�8x[,��̡��Yj����TeV�J��w��rH�@�N�+�<��2.h�%��/5u��ixXU�
_�[e�inö�Mm�w(hG����/)-�(�!��^E%�=Hې3�r|Ϊb�2R`xF ��s����ۋ��n���K7����2uZ���P�����z�s>Bu%b:���=����4�l��ʴ+�2�	L��	���IM��r��2�+��S�=M�p!>���v��G�;�d�Q]��H�<��Gw*����B@KL�Gr�>1��j��.�rJ�C��r�|HL {� {;h��!�~oA&P{/�Tjޙ6R�7c���ҹ�FI6����+��Ԛ"^�D������ ��* �1�Y��k�&����	M���I6B�U0W�^O7�o�I��?��rǓ��C���l_(9K�|O�]�y����g��14>_�A�˪g��وA�Ѵ� HF�-*�#�:6	�JD��1�8���w�U�z�B"�\����=gdm��Q/��yqn8�����7�0m�9\�=jA�j"*��c����9���%�!��G�a���~�W��y}o]����Ch�ɴ����7��Uߦ��Wn:��0�m7�<L<Q�>��׷��-���-�!4\��*��u�u�b/��r��է�<�ă�NNo"���y�8�H!~կ�q��0ն����Qwb|;��RF�6J�ɺ��E����	5�~&y �[V#�:�"&�³F:��y\���X4�YXsF��8�d�X�bs��Q�S��1��|��Y�!>��J��nL�]�tv����|X�h�f#>�-��v0���Fп1�}W<���Ղ`*feT�5�n������|���?`kZ^�i�+�3t(���H.×e�F�!Ύc)+�r`;:M��L��S�����`<�Ý �M�v�F�5��d���=9�{��#B�6�l���9�4#�HZ� ������w�
*&D�u�Р���,6՝�r��Xk0����Z��S�Ȃ�ɯ���'��@+�gB�h���r�Ϲ�i����.�ڹǱ�"WK��`��S�`�DGѵwl�^!ՋU�:W���$Ӫ�8�BSm)	ݤ�U:��}�0�"�K5'Q雂�ρ�J��C���L�B���p�$ӆj�:���~�D��3����#��)��m�ճ	zݵ��|~��	.���0˜�"mz�C��>�6ӪN��%x��N���������Xm�ja�ƧA\�Ԑ�>��4���G����N�Ҽ����r�ݐ�	Su�H|��a���U���oKa3�
�w>�Y��DEqs�g�u�����!����
�F�Y�%��>��4���j\���؁f`*Pr��|}6�ʡ	����E��G6��C)~���'+��<�[Y�q�#q!�:�,�j�G�T3���KČ�!9 פ,�x�G~�,��w�W/U}N�#e8P��F�	�+O]���1K��w��Wh�ӥZ�!��)XB/knQ���:�K��Ǉ0K�1��5�R���o�:�B
�tac�
���r�rK��iE��w���V!'0��P�+��
�t�)P�B�����u2Y��H|ԠD�0xCL�ʼŊ,1;�4�b��p����Չ(eT��l9o��~�N��c�9B�%�)�zE!A���G����y3��2��`���.��9�����s�����M�8����}��!X$�U��n� �6�FR�H8!���縀�F�-6َ��'g�x�gzSr�!!fx?�q��pEKqi�q6gωC��V�Y��_�ߐ�i�o��?���S�.�Q�a��Z^��Wv��� �̞MB_m�Y��ey��R���-��T��.����~��zϠ
�q����'���^7��i��L�f��N����Ό:�auT��=,�=�������/��=���� '�/ٱ&�#E�3CVea}+RH&H���)eĠ{�����T�ꊽ�%I�sA	vZ�>����ʏ�-:�퇟�kL�Zm-�/H"i]�Lp��^�nh�����;F��gO��[`�XJ�Q�Pw���7��t�k �8
�a�����w��ʡ�����B���"�1,"�q������Լ�=_�cP�[������2b�+�p�3�����^.�Ў�i�{�����II�K�����j��ؖߍ%'��i�6Q��5FY�m�!�˼Sji�T;��W�SDR�a!�%�t�?��Ϸh;c���v\�M���<��wkD#�w `9h�_�;]cOg���\Rf�~\0�9e,h��+MI͚ؓ�oVaL�5�R��4}���Tac�qe�e&B�����W��D��Y�	vp���;U	�3��2���B=A�Y��N,<�`�]5�б�)��ށ�t.n1{���xE�f����{��=����(��N���(�.���X�c����	 �8b��2�j��� iH���IfNj���nέw�����0�M!	�o|�L�ZMx�������\5� _�[.��r;jܼT��z�n�� ɓ��U�@�}�S"w(	C�s(<�r��i�N��}�C��/`?���9hfQ-=�l� E�$~���p:QC����fW�/��L���|'96_	o������ӃH��x�̂ݐL��`�����2�K`��"+�i�()S��h ��Ο&�x����ٻ�6Λ�K��~���VD�ʭȂAhY����g����4��]B�b�E"���w��4�h��s�d>�e��v���1B��A���=�\!q'I'z��K��F�{�方i�S�5�C6G`dv f�n��>[g�ߜ��c�h}\�W8�2Z���_y@#����An)��M�3���-wm�{E0��&��(�?%ra�5��}T�s���Q!�+�NB�#ꨒ,ID9���%He��{�b��F���ź�i��ZQ�D�é�� ���>P+&pJ��������c�>��>^M�<�[���*2�8�e2�i�q�j��O�}ǫ�O��Uu�N8�h�"_�p�BU�?F3��*y��F�չg�~�K���#�N�c�N��Y\�9,�{У~<�[Nn�a�9"c2σ� ��"��h;w�z��Y�-f$BӓPD^�	^]����ߪ%�"z�O4Nic��+Vl�E���"I���p�5��47����u�<�j�f�g�i"�5N#X�������o��2���G;�2\2����s,a�=僩��u3)v(yZ/%���&�]���t�Uҷ��74��S�"�hs䱖�Q�&��%ׂ�F��E��~�E*B��?Uh��+�q�b��w[��."��U�GZW��t��߁���ٮ/;���G����ﲡ�G�����OF��i�����<���c�����Ae_���wx{C�0`m_p_��K��pum���DT�~5i���9�]�/b�g�3*
B���x?)��u��'"��u�&/zly��Z� ����6@�3���J��H�c:0D��"j�/�n�/3��o��pC�c��K˯GB&��B���J��]�&�q`�5?o���[^ӿ�Y�'�Լ�@���g�MR����:�Cȡ�-�n�A�����T�^r�u�[��C���y*��{6���R�d���Ko� �:ꐻ9�x|X���:��s/N�h��\{I�C��>�д��Om���w�E��U
�'9*H;�hU`��&\�ƘOz�v�$KN�0�����QM��nHB$��H��Ӳ-�4�ڒ�'��u��������L��$�"�W�Z��ćԭ�E<��W4H0J�'i�#��2"m��+Һ���U�!�s����%le�%� Gt��E mf�9��@1�=G6��$�}��jԽ�#'�3���b|9;�g���9�[�M��}q<�;P������~�:����\@pb؅�2k��w��+-`�9��I�TYE�u��>��6�[�G:��IW����MR�=�4I�z�s�x ��\���.�g�������͋rK����\�fӸ���J;g)�e���]��L��4>?o�\kˆ�	0k%ړv�1�d}��������?�NI�͜K���@,�����l�1�� ���A1��o(V�g�_��<���&�VͲ�*cg-����.�G������\A��L���5�����OT��!/�LS<тk���>!ʭ�X�����+� ��KQ��ˆʹ'\E'��o>T�5=�+M#�&�R�������"�/X�X��Lv*ѐ}�orB�5�}#��)�LѾ�CE��xk�J�Krgg��Ӂ!"[��M�4�9���:�8�C��[��,� ���qrُC
�A���WG���
���� ����{Ah\�G���|�Zw� r����]��9=Yx%���l��es4M�|�����J�ʈ������B�@[��,���������li
��H�
����� ;.�����P�Q3{��:��׽[�x����½xd&~p��̺j����<mM��A~4,K#��Bԕ���kB\��Q��!�'q6��b7�e�C=e=af]C紨�N9����@c��\x��7�=:�{�5
%��D�*��*�#��?G�����?jL3DN�I��N�U���K���+�G׾���<�ӟ��^����#Rk#������˱a�l�+��&W=��Ԑ6ڕY�
*} �d�i�õX��;����L=ėO�²U:���!����x��~*}��@kL���Y"%�ăi�����'�+D�?��+=�4�kH!E�7T�q���3�R}C
j��f�[ر5�\�`&��s�`�������{���\{m(3�������pt����v���Zm����,�sz<|^�/$�U@/, #K��})��>?"ԌԍJ��ƍ�Oƣ;��F�y~�@�{;(���&�ogRi*�&�87�&���D���l����F��7Q�dTy6�O���>�h'i�KJ�^�68\�u;�O�5�5�����QnJ�u ���4�yL1 ��q7�B?��+��b�b���=3c�!߮�h\�p���_��ihz	:lh�n��~��S���'�2������,*T�T�kg�A��k=^ "d3�x��L���6��(���/���`�F�X2qj9M+��Xڗ��z:w����5v2�SK�o��s��k5�~,9Â��t`��S?w��}~�Z��3Wٚٸ"�����͇�uuc^V����b��GY���!=ŀޟ�"��c��q"!�Ğ�/"�'�	~2�%��������(�V�54A���x�kA�� ��"[�s��B RW���������%�/��٪��u�c���"�	Hmٙ >֎R�˜�M�m�(u��9�|�C�e��l�|,tf� G���L]�,�<k����Fl��Xau��k�|��M�A?;�{N֧ �χo�Њ%���t�pB��#et��*��0��?�7�)���,��_����{�l��A	�;�֎{+S�?��g$�R�Y���lgB���e7zP��O�M�!$+u�@�����ۇ�u>�?mɓ�/��f����%�����I�����l�rO�y��S(�<�����]{��ث�6�[%B��
�U;�x��-�`GD���,6F�PأeRU���Y�H��0,y���v��lw&��ǶP�Y���$��m4�%������w����5����}�2ݮu�6i���]ђ& Y/���T��_����N��6�t%|
>�U��f���l��=���ZFF���}���{H[�>���8'���v5�&+5{���7�W��P�tx�<;X�.��6MO�Yk�MI�kQf�~�n��#T�N/A���_��I�j�
'O�����h��9�A6&��t�U<�L�O���<�f�����?v"�#KQZ���Z�$^!�zNXtF�|��|ycs�تxq���:���y`VR<.7���}��Y���z�(���S�7|�pA��p�� -�/��p6Z�$�M��!�24�t*r��m@�.k�=R��d�T�<J����ؕi���R�D۳D>e��Զa����ƎR&:l�n&���eٱ �'<���2�g��'�A�菳��2MF�ï�k��'��3sd"��a_R�N��0P�� U�)���W�7��H�C���G"��&g�����'#҇p�h�S�G˒�MU�� �#�+��o�œ�*Ky'�+���X�2��w���+]/@	R�9�ϐS�o�E�$���	�@G��\�����)`/�3�l#ő�:`.�q`2�$y�ھ�B���B�����4�k��fY�t��o���qǒǠpw���BI��O�RJK�0ӟy���g���vRWPQP��<EW��Xi",k�ꗤ"��Y9�q��!}�95�Q�U+|�x~�7����N�j�v��j�lcu�Q�`���e��/�Ma^�%Z�;�P�fqDЦ��'
�DD���
A%�x���uK��mϧM��Ut:�Q��m���І�'J[k�ԅ�ݭT{�9#������hߟHHX�>�����H���,���Ş��6��	����zx��*(���ǡ�h��l?�@ȶZNYi�����O���Ju�!.��������5�v�`�g���L��g:�g�٠��yqA�VR���.��h+����#c*�R�������Az4�l}�걤���w���(��Ux��?�=P�AF<Y�/��@o�!8N٫HY
���zY����У3Z�A�%(�#W���7��1Y���;y�'�&����r&~�笟J!2��Tw�AEэ���#m��: ç=�VW=�����=쒹�<�^����'U ����N�#�SI���2m�Q%�/ �������L7����[c��$W���4t�|�喝�7!tS��rc��{���$�}�t޼dK���s��ZD0c�M3yg��)?$J(�(5C[�����vU�:
O�"������ܰ�����K��	J�qH����@MF%]xM��4�o��v���^ה�k覴Ì-Թ�ӝ�W�������B<�R�� fp�Y��MS������
����(�p8�%hbX���i�ڄ�|1��[p�dI��+qV>�z�b^I�acV���ш$M�f� ؟��OrR�lੳޫ2����#%{ �fd��9�y@|E]����g�����=|�uCi3$�����Z��y�!�z=�h������W*ɰ��J1r�{K�0`����!��4�nOR�����#�9�Mz��� ]$�ł��g��>���ڳ����W�U�>��5��2:J�3B�O�~�
���$�>MP��������g�q�w��8��i1�����+2�Zd
M�!}�d��;�#e�@� ��ԅ�Qy�����᧰��=��(��"�
��[J{���s��g�j1a�D~�#�n��w:�؆a�Ų��m'A�G�R�1��)��Lc�񗄕D�b���f$G��tT��� }f-�u�v�>��m{EUidxK`�ꄇx�9��I�۬8�¶K�E
��A���B阨@.?㼍�# 7���Nh0}Cuv�W��x�.�uL3ܩ��뀀E��0�'%�g�Wù�$���i�yF=Y�X|��"r�ŧu�(R�1q��V���@
��zp�G&�@�Hߛ��q𥐁�Y@B�"����r��&��o_���ω��It����E[�v�i�r��K��{���G�� �F��i;%H�X�G3�u � k�O6s,]�Ă�����|���t-���8)U�ŧ�h�4,L#A��_(k��dqY����j��I���#�ӱ�5�6�M�+��tu�d?��@�]�a��:�=�8��7�s5Cq��κ�S��84W��"�k�̹3n�igɼ��絰}��|����'i�EN7���Q��~g.;��J%FGD��x;A���*�\�9��*(M~��v*9������]����M�y��-*+��*�5�3�#YqO�<u-�Q'��jT�8�(�e-���.=�p�|��/'C�T�9W�걯i� ��x�m
�x�p�h*��O���PN�j�O�l��G�m���\XT���( �s����Qxg5c�_���u9�A��Q7`�+��m�7���/���A��a�lԭ��� E?;_rDa_w�sp~Cqĺ��Лr*��U2�&��r��b�j7�Y%��.�|�j"H�&_+�ޕ�� ���Y4�IO JfU}�*�f��X�e�Y�Ѝ*���Q\�~�0y��!����G�����N�m�G�)]j$���W�ty���1Éq�$�@e�2q�e�`(4Bd�)�ײ�4	�4O+�����.��Y������	n9�|X��h 9���Gvd��v6�ϋh=�2P�fr�K��@�ջ�s�`��46ae��%x��+$�V�i���3=b�BIu	��zz-�;�-�~V!	Ȫh= $SΘ�SY���
qC����u%]�w�����Ro�n��/:C6����"�Zp�DΌ�J�	��eƥ��Jrw�kפ�	�����~w��ӄ)T�d�ES����Ġ�Ƣ�|?�N��ҕ��U'��ɭ�SA�Y�AZ[T�i$�Ve�o-O�	�@h�T�i�dS��e�W�sCXj|��F���Y��Zcn	�^�q���2�) ��m���3��:_*�#�.w��Q&_��50���&� �ss>��>]%8�5��!W"c�K� S����o]��f7����oϐ�B|���)�jRsFGe§b}� C3�"%.���*���8��G���O����� �����Ԑ�"��C��X�baA�3�����F�y�(%"���܄���]tZ(�������S��Mdnbd���C���8̣�w��Y+
�߂�
	�����Ǐ�V�%���W��z^�.=P�^�TTC�7�\�d�)�=�j���	,���6K��Q��4K�fd_�btfY"�<�^���}���?v���,�kјkg�2���:zCw/�Ncj�q�������]�_ ��>�CRǟ�,��%<@�K'_:6��X�3Z8!H���]fQӕq0(&Η��w�?��~"Ɇק��Ѓn�~��F���|�y|:7P]6��4���_ ���-�JEj�_���	1A&vW�,k�#$�ą��9��e����C�lG*W��d_㫜�RJ��7E5f5s_�����V��q@�}3g���6}尟Np�7ΉNj�+���S=��
\X @���(&����H*O��4����V��Hem��'����j�'�m|K���0�c `�<��T=鬃Ě6*�;K���3[�n1Ĵ3���ʆ9�n���^D�{�����(z MW���P��8��>�^�j��[N�������f��[�D� �nW�y�$�l���-��K�$^�GM��Y�TB�B�"�EMQ�> ��h'�OU�26�Ā�<@�'Ō��{��l/+>�h���� Ѫ(��L�<�GLPKݠ4>�Γ���ʭ�S6AQ^�T�RA�=���Y�ub�z݂�q6�~��� �&�|Zc���)^��EG`ih����b�tO.<�Ip�ޖ�~;�@2�����cw��h_j�T��J���U�+�x��iu�"�@ψ�a���њع�����-7�2��P���
��,M�����Z-hxN�������sj�d �X(�T�� �J�������w�l�A`͹�G��[�,�qc�E+��蓒����`�}5������j�4�ZE��c¢�М��78Bo%z�x�M"B
^��6>Z0�E���ៅ� q��AY2Ɵ�L���q�uB����;�7��mM �U�$��JC���Pڕ_A�;Jj�_GĈ���,#*z<�b��fLI�XSn�
})̈́[�i� �$��{`����3����ސw'�+Zj���|����@_��5���.v	gH'�{�(�e����q����QN�	��g�i��� �ה�n=��!̬�#C=$'���̏����76ؘ�h���`JZ:kL�3.w���NZ��
� (D���F�v���������1 ȟܦ�¤�$n�5�YH�t�ݛ��ԁ+Z�bd:��&��!�CR��:�Z��2"���\����B7���i�U�������L*��^�P��Ҥ�͛�p�|E�@YK����J�]~�+�W&����S���n¬BT�#���rʥ���ub�G�W����M;���?�W�[������Y��i���yD���^�SmY�+�p���� �J�e���?*Rc&�� ��䛫���$���������\���/�툄;x���ȵoW[�"�]X�TH�:g�̩ukK�*���p�0D�"5f9�׼"_5!�f���&~+�e�!��M`5�����z8�L'�j=>���o-B¸o���n�OE2��)�e�ߨ
�!,���(�!�Zl ���Y6 ,�3'��#& 7i���
ն�)!��µ�鄷�O�RB��h'���?�I���ٛ�Ux�q�]Z��M\B�ȕ�U��2��Z)���>���:��2z���s���'����m:$Y](2Ï�a}�K���.��s[z�<
�!��	�F?1��v-��v�0v�CW��bsc�$��0<�,0��PV��:�^p4����bA¨b	� c�:��l��^S9�;��%IW(�Ha��Ti�|��b)�e������*_b��&�f}w���%��qC�o��b�#/����������T�	�����i=�]Z��8UVߌe�(_qT!oK@Y�õ�qH��)ޱƤ�ʰÅ>����3 ���)�
R��@�#�3����1�[r��?hlC��)bj�X(�R�C>CUܤr�]h� ����^�{�w�;����v@�U�|��]��g�~��&)9�jlT�Z��a$��X4�AD��M)�|��=�Qj��`�`��q��$쐎��c��՛������Jȡ*���$+����ba�{��̵�N��Ax�����b�,F��&:��ġ�8�B3'�KD���ǰ�C9W��{�6J)���!qIa�f���]�u�񏇓
�������@��2�ř��֓?�[i�t�7�T�獕����'E9�7uRZ�$�����*[�y��M�hR[Nn�� ��UX��o��l�Z���3DA��)X�3�D��C���8���Iɚ�f}���T͸��]Ri��Q��h��
�e}��w+�l�����
g?.Y6?� ��
J��&O=�j���\H���8x��T>J��R�N>�1LM����+vŁ��k`�0n�Օ�yq��-�=�<�����DG�l+��M����k�G���eT�����΅�ֿ[�T�材J4(|��p[��isy��3Џ7�#�������k��.YO�����#t�b1H��
b���q\7�A��^�wG�F�(mD_� z9��	���ށjd��;�.��*���S�Mہ0�|8�}�]���eX.�v�� P�{�$�opr��>��ĳ��0n[b�_mĲ�ث�h�ڽ�>�=�X��E�5ȅ/�8��*�����Ji�����V-^$���<��kt[�b�d&]q`��@�K��+�����F�36�ُ�� z����	�^mO[ ��E��y��}�����L�6rܡ�P���^+��t���OQ�G�:�'<*p�y����C٠)��iԼ}��<����)�i������J2 
e�o�fhJIgG��^F<A)���=�;D����	2|V"�o�X` *d?3H��إ�u��S��r�ǄE��F�,u4��ΈA�	5 �B��UK̑�,�ᇤ� \����:�?��s6U�D^u�M妱A��h�^@?�o2v� ��~sd��<���O)I뿂�:Ԙ�DxO���:������|��+�ѹ�z��O�!��}���N�9�(Gu���;���̻*�C��}�R���j�y`e�
`��d+fE��uI�j����B�jtDH��#8���̱]���W�u_?'P��$�R�>�g6��	��o���P���m�i&�m�:ǭ�ͫ�ȓ�퇪?� LJ�7yyZV|r�Tq�D���ɧ�����	��4��f%2<�z�1��}�g�:�lId������D�\:�X4U@�������B�u��;��c�C�O����o�c������FĘ����x߃-�=H�>2��u�� 4ۜ4�gR��1Q��H�[�<�;9l���5���GR�����a�6�Ƴ�8�.%��m��Xa�Q�j8ܲ��5$rq#�#��`��t��"$��+�e�}ʹp+:av���b	��V�$��F�UA_�`!� k�Q̤���JFT�nz�1ޅ����زힱIG��=��~�����H2�C�l
��-O���Ip�$�y�v,B&Y�z��Aѣ�ns6���Ze�%j��s�KT��O�Y��tv������� =�q.��t�:�]�����ճj&��96�'3Ab=�[�u��	d��b��+���hXT|�W�_DhN�eǖʖ>�}�LqL�G�P6���z�G������0�:�N�8V�m���z�&���^?+J�eŒAh��c�r򷞙H����3�Px'���W��7���M�!�[U_'���`�Z����	}H���~�}�JX��]�-݄���3�3�'� 3�w�j̨7^k����-e �e��Gp}\7 \�q�%�UrpD�jq��ƁL���4/������k;ƕ��
���U��dZ��,�����چ\�N:�u�BP_Z���1���{iY�zi��G:!<��Y�s~�:��C���#2'Q:���n��/��*��*�~�!@E���F�������;�v&��L��
�n����Lo���i���-o��ck���板n�c&���i���M���{F�X �L�o�Bt����-�R�r3�CHThw%�X���TN�t��u1��m�> `�����~����ֿL�(��!k���r5[�� F�ѩ��Q�]��F����~����Ӌs�D���N���&.�t�4�*'��#�k>�jՅo����)��pg,^�a��eއ�����o?]�%�,���k1�2�8 %���*@9P	_�����f��D8�eu��@]�b#�M���e���|�5�
�*�r[=��4�ʲ�w�
�".�t�S��"Ǻ�]��ґ�^�"���u�[��y>?&��3_��\Pb8HOqO����{kU\1����>r6\��rdX��,���m��2A�[..?��pa�a��1C�د@�y��
���>m���y@��ȝ��b��_d_&��4s��`+)QO{j�M�bJ9���bC������B()�^1%q�\,r�\�	��7j�O
���R%y�N�ri����(�yk��F��Q�����p�l7��=�i�	x17��Qa�i��i�Hh�ʴ�C3B�F�3�c�#`�9�yH�2Q�sl��S}e��͍���{H3A�T��3v�=��j����,�L�WӋs/��(�/�,�k�`$V4�N�:�2�E@�lH�v��b��w
T�띟��^8�1���B� Tb�ݿq����G���@RDɪ��rw��;���h���n�v�1�>XJB���q�tB�JsX�7U]�����vp�~w�#��2̭���Ԥ�=�o����a��� ���M�B��D��!�v�A36jGb�1R?d�IF!��L���M�4_�=>?Ai	Ƞ�g|��)2������#Pfq�R��a�w�� %$&%8i��s=P����T�E��V�Tԝ�ln,f�oϣY�Ky������6�����p�T?\���uGٽ��iб�K�5\(��8���a�JBs�bZߗ�Q��fxC!�_u��k��o8R�e��و�w�\c�	�F��k�w��fYZ^�w��k׿���W�q���Q�-UL+� E�~�[�������Ua{P�+�y���!s�� ����T;�Rϟ1�<��=.��)�$�N09�Ѥ� _XS�����0V�&�N�,���էF�4�s�.�Qx��=yMd)��CZ�Wm���Zh��_.���f�!x��&�wr���'40r���������ii��[��+�Y�5'�D��B�R�$�)�f�^��$Hau�2�{ʂ\��¼����s��<���ϳR��%.��Pp��;�����}Hi}+��05a*ܻ,po��ϊ�ۤj걈<�ȵ�tƮ_)\PU��.��ˋ�DC�h+�F�ǃ���{��f/�lJ����
u�u����!��Bd���CY���W"�M6�zъ]h��#&��S������&��4�ϝ�ao��v��87��;Ζ��?#��E
�W�K	@9k���}���PHd3Vt�$|Dã+���:1X���>�k����J𥙗%�u61')����ۛD�Z��g�����ԇ����f>l��k;7ӊ�3����##�;s��$�Ax���k+�8}���J����~���ب��	ߟSQ��?��{ؑ�wA��`����yՄ�!�g�؍i��;�n�/�`;%���4�C�-b#� �Il.J���Y��2�4ד'e�-��6��ZA��3yAt��(��u-��P���j�*�5��UR,UD)Y����gʠ^ˌ��  ���H~%3�r���#��ir�QJҫZ{�m�+iA����50�zj*���f����8 �l�<�
�W�C���`M3^��D����P�V0,�?�u:�Y�Ac�R��30X������_����6�|���+������o6ӻ��S?��0LƟ�1�6�Ʉ�� m[�v����V��ѩl-=@<	)��P��Jd+�_���n�j"=�ubh�����*	�ܜ�O��Kg6y�䍭����n��)�o�˱��HVZ"0��3���SMμ$Q��:]�f����b��!ŏ6����b�C-�PN���细v��43�!AzЫ�"�u��7�җ@�&2�R����j�Afc}��weU"����m��c�%u�WfbDP�uJ�ϴ���1b�o*1�>}�Ϛ��� l� >)
Ƨ���j����o_U������@nT����!{��v*�������ԟٔ�����ƿ����<:�Q�A�9mx���k�NJ���q�'����"$W{�ɨ��Pvɫ���Nܼn��C���S�7&
��~Քa����Z ى
3"VE�@�k�����*tM��PX
������#pT�D�oѿG�w��d�/"6#�Jl���q���\i#=%)����O�B��
+N}f[�>f^��'�6���8�%�=�z�ҩ�����)d��G"E�ʲz+W�N��[ ��f;�Y��֚���E�x�(J��_�#D��0F��7�G�b�,�LD�<sw��ރ�u~lj�rȩWթZ�;�8���?�_Wف�7�8��f9��JmO���k�P���Vd��DN�8ż�5	�B�3"�VR��XuD|edBNw"
�����5psmU �����H�ް���~(�X��;>� G�t�5�3�A�0��;�0y�;��M��4�G�%�k�:SP)$g�j<s��3�3��ȊEF���[;����2z�n���W	f���\qX��m[p�|m!�v�
'a�^��5;���)܅M4�|���=���9$CҳYwF�3���pY�TP=��$~f]�~���%
�%�����v. ��
��T��c���1�n�������R�mE��"ߡ!��8ͳa����.������)_^Va���ٟOo	�@�?� 	�U�Ս�J5!󉠰��������;�A[R1�8���F���pg�#,���M��rգJ���\��O��c�N*������ƣ��-z�?�@�}�ܹ祿�EА����
��S�?���'�{1�r���ڡ)�G�k�>4=h�>�C}�%vf��6��Ɏn��+My�=6rYn؍"|9$�qܴIÞ[Ƴ^6!�,�_���U�V�RO�G6�ph�����ӟȜ�t�1��U��B�m)g�t,�ǳ/��a#��O
�����Lm�Gfl\.C��vLr^�D��
w�R+�r=�6 -T!����BG�e���G�	B�o�
�~���s�/!����(�F��d�L����8Mׇݐ!t������	��gř�~��~
��6�t9�Y�m�:��X��L�"�`e���Սs��i�����n>,i8~N_���WATC�n'}L'0��F�[ӓD�n�É@7O�RBs�a8��g���;^Qpj�%5*9`zo�$�k�d�����R����}����Il�N�i�=S�ɱs�ʠL�w\f��H�i��]%�g+=�9<��D1����>����޹(���O³��M���
�����(b�!G�}`1n�R�<Y*����j��bC�?����Ӻ|�:��pV�7S1+C�;t�B���X�\���@���*��ۤ���A�3�}-m%�O^�s�)�:l{�ln�?G(_�5_ۄf��B�r4{�$���b���\��x�P�n