��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?Bk��nߨ\�j�J/C E�6$|dȂ��^�#|�r��ݼ�L�f̿�A�2"��^����a��;ȁ�{N���Hs��,>߯r��$��݅�}fEm7=QV}ŠB�:�NƳ`�!~:��7��u�g�V,Mg n�pi������Px�8��{�E'��y�<�Em�p�鏡P�oд��ǧo$��a�wKʮ�!�E!���t�����S�Uqʔ�}ET��O�}�YK�8�tY�`ZD''�/9�J0M���f�b�D֢��M�9����������-p~xvl2 0́À�G�f�0��ҬRL�:0�g̑�D������O�z���b�W�_*���3#�7�>�J++C��?w��L�m]y��R���M,�O����}xm(���?-\���zh�(����
:�u�(:�P> qӦa�/I{�V�-BMv�Oerr3|{�v��.�W�i�P�3�+�]��-�:a��_��R�7������筇�h9��R�b*�ծS�;x���֮�t%x��R���LYfq�ߢ�V�ض6M��Ȳ�5�����T �<� ���Iߑr9+~��o��tBMVͶ* �^��^�K ���!a|N쨷�.���e����`G幼1`�#G:l�ΰ6�83߼7���Ļ�-�O�7�#��+�f}���R_n�;��>��%��Xse�]"��h�LV0��;tq�Gn�\��uR��q?���P
�i\Q%���ޮ%"NZ�Qd�y�&`�jx��b	�vY۾�����R�1ř%�ϩ8LJ�ƺG�7����)T�o��ǆ�P�b?�}ɸ�W�p�M&!���>:S�KB�s� <6~�W(�(F��ݟ���n0k3u�]�i�2��&2�w���W�^)��:��lܨ����yip����Y%��� ϱ����ٙ�˶�P;k]��|ٔ�e|x�U"�4�N�Lx���C����=�􏃇��⭄	DJ-�6J~�_P�2|k�6��0��X�l�Qc�C3`oF��i!��)���..d"v�*�O����	"������g��$ى������[�L�U��,O[W*a��a�FI�![�I��h�ڠ��v��"T�z�vU���\��77��*���Ny�><P�k�_P����`�S��I�`(NI�����"~�M����cz~C����� /}�eǑ_bf�GU���m�`��D��8V"5es��Zsw|I���Č���OJ�{	ZG�635��kK��d� ����"��=m	�a��S�&702�ůBėE
�Z���v��?�Ny)�O������K�� �dVg[���e)�� ��#
��hx�I��=�L�&)S��yv۷�F����+��q�˃6i���G�g�G��TE�7kAJ��74���E�QL�m��{�m��!,�I�)��~C� o3Ћ2&�M�a�B� n򃋺͸�K��T�ZNR2�26�f�}�G$ o�e~V��y�ݱ�
�J���(���+t��,y��
?{�>7�
��ܫ���Ծk?�=^�.���b�e�HS@���]�����0��<a~M�݅]j�RZ21�hC�I�!@c�����Yh'5}�j8��X������I�<�e��LK�~�����Y����:~�;�Ƿ�l7�Pp�+c+3�4����Q�Y�+�N7#�Y�0�2Y1V�7���Ss�XK��ΡX��W����B�BK��0�s'纖�A\��߫,��#~�>��r�lks7'�� J�^�9RB�M�
p����;�L݈��Җ�@��9����F	��nm"��ipr3^�ͦC��ԏm��q��Y�_�A�phMm�Q�(G�hds��4��u�7���OKU,��@ߊ�%���0�b��Û޿8w�+�\Ow9%"�DӉש@u�C�(vF�����$r�m����`�Hf����o��3кؿ�֬o���x)�	iW�P%�hy�ۜC�ĉ����5c_���Ss��a=��@�E�|�=��?�cy/g���77�m�@L�#<R[�Y2������F�"Xey_G��BR6Ӏv�1�bb�L �桔0J�l�f�@��i�ǻRTA�U%��f;n�����"���SM�Mh�;��7�j#�N�<�k��Tشo������-&V���Fk}���d�ic7��=����d%BC�$�cO]tȹѿ��8�M�uj|VD�3���r�6��LU�2�?\��Ħ�Wӣ���nDWAc~|�7�<sJ_���l��c뾀�@�T�%�dG0��+!C���Gֆ ��kO\��2���Ϲ��y.sވ�Y��_5Pn�o��'��\���B�&tj@x�o�a0y�������A��a�a���Y����5Ŏ@m��^w�$1�x�q,*�0�|fz�G��c�'������-OC������3�D7�]n�8#9��Q�~�
��JI���U�/�f(�ݡ�1YQ�j҉�}Yk�0��m��)�$�<\��tp�)�ש�����wة!�
�9�C��)®�滑��%6���nqa�"�K�=�E����[��kB"~�i���#�k��b�:��JU zd�.��k�ca��[�8�V�,��Z��}�M��X�����7\���{>��$.5�����T�8���~<��4	 	d���;���̛�)<0�A�d��<x#���!A�*�������l��r���*�.T���<(ё.���E�vl��#��.���k-G�1	�a�����?А/�+$,�'��"/^M��
&���ٿ�6�U����6��H�gn��Q`�b�KO������S`��5^U�����<R�l�����0t���tS�N��}b�j��B�S��Ѡ�u���, ������~O�� 5�Q1̬:�����<>���+Q7�2b�i�Ÿ���?����D�uD�S�soF@USȥ"��-��^Fr[W�ۦ���+.!���Yqi�弳�H�#ܤ�k�F+�\��t	8�~k�m�����ۤ���'�IT��
(r��z���g���F�viM����G6��Pq4�8�0G�'B�\'vVBOZ���e�'?�<-���M��G�³���xm��7C��q>mO	o�Jq�/�����F��k��:P�rX��}��O(�f�c�F�%PWMr���̲�Du��v��yx��w�_Rf��aw��J������@���3�����2�_rTa��|[��67���Du�j��rB���6��J�7̹(�μ�-��A�(���vo�qD�&.@KW}C��Bl�Da{�xAޜK$�WGoFVBUU��iS�@����E�f��o��	�8�t����|�'�>uZ�Ym���������L�M���;�Q��BG�����u8��A�}��EӺ-�W�f�}�:S�nT�8�V�V��w�ܪ�f���R�����
-p��i�Sv�f�;��{j� 꼜Ƃw��vl�����A���R"�t��G�Z�,�(?��4���F��5�G��TT��ċ�q}���j*�Z�:�	�)كq���W��z*�Gt�$z嵉�ܢ��(�>pW\��-������]�
	�1�	�bP�*��fb���[�C��RE��׾�1���M���z��e���)�6�S-�����M�U���:uPc��wp`�'nޡw��4:F�r.&��v��:���ε��Ϲ!6����+s�3�ݍCW0�
�Dem N Zs�/�Y�b�������ޝVL��R(�H����*��B�׈;3 <9�Pe�q���7��NEѫ�[O���*�nl�CF��b��N�+�8�c1F�|L�
tش-�z�����R+6B�{���8w�C�/\�0�%�t|��äc����p5�!}� �`�k.�#qP�&D�d�\��8]y�����P��g�Fo���'H��3�(��������Z@�@�l]`���ghZք���*�f�'	"2D^MID����ߊ �,ӏ���Po���ң��lP!Pmu��!1�F,�f/�J�N�%�e\���x�`<S��A�];!<+��'	Y���]�+p�E��ňTߪMgͲ/T&=��*[
�hP�j�?9�S+Ymm���?G����G�o��i �� �'�?��YN&x/�
l1]{�=��]o���՚��];5����i���<�ż8�4��tyT�U�Y����6}f�3]�h��'�P�g����>7���L�����s��҉2�K��Z��[�i�n��,��@�NO��N���dv��D���c��ȉ������%3���W�vEY�Eb[t��d� �5�nU���dp�@�Cgӥ�Dy��S�k��c
�+o�D#��e����Q�>_>��5�!���S�8.�n��aG��`�hc��.F\0#�.B�}mFN(gf5�"�c���*N5�%�V)�-_yw�Aw�I�E�9������f7�*��5G`�5�A˦�@Z�]�"��~�fh�z:xY����fǲ;[L���h�V�ѱ���E��ae��F60��H��$��FrKL��.�z��8��`C�0�����F�&�d�V�bؚ};��ޣ����d+Ey���h�,���)u�op�B�*a�ὡ�mA9����m�!��68��L�XD�Z�����V��_Z��s@�2�J~f�Vq����V���D�Vp�z��Y���"�����0���lձFu�4��N�<�߃#��1��@�C�.`��2Œ�IN��J��W�0gE������=!e�u�����&�(�����wү����L�Oڑ����s�L�b�Z�8`u�e"�ܗ	���Y�Hǫ��VO�K��v,���S�&q�x@rY�n��'_�v� #(\�S�Jח��%b%�j\�7h�l.d�نhu
�|�e=���2H�<9c�&�����nԖ�	����)a�U1w<���n��1&�.���u�!%���y���+�W�ն%�����'�P2����R��0L���!F,�/a�"�����h5
% ����֌�4>:��^�0Pd��z"6�d$���O�?�y#�`rԭ��ބgf̪��{~�:#Y�K���i�R��:.U���6pZA��n'�8?N`LC��C�e�ԑ�;r�"sKxՀ㻿�OB���"��'EX6��+��dN^w����ɡ�Y ��[\^$�������� ��ϡSKBf�/ن
o�/�KN��%+#mlsG�ž�,���1|��縅�4d�T�Q�Q޼��5���}��Ú|�����a�@Rw��;�9�Zn+f�������8��p㠜\7��k�=�|��A!��Oi���y\%z���S?�ja�2�1t١�͕]cX�	���׈��.�V��8&����gh9��d8����C�YXU�e��{
���|��f;�2�|_Z��������t�<ѥ+�vT�vN�v�q�NSx�TzLRr��v�R�Uk�G~��\ޢZъA�8���By�1p눅\]����=C.�z0(�w�+��ـӰU��3.{is��܏QH2��e�LZ�uފ������=ç-�]Wo-
Z>:?��L�/�_�\��}(,���Lf	YU�i����8��k�bn�x4��4�Biv��J~@n=�Z�Gr%^��h(�N��tDb}8�_���B0������qdARX�v���q)	���ukp�X �|+��  ��t�����ܑ��$+Ax�#t
v�`�����lV���s�%���r �C��f�M��ہ��ue��{I!���+�P��}�P<���.���w���0��L!3
d�����Χrks��T�	M�.O`���d6X�6zr�$Ź؀���+�!�s⎊w�=��	2q��ft�ւ���y$-s/L�i�Q�hI$�ÿ��zC��zy���֤�n�L�}�M9Ɗ�/Jh�4������y<�#�\]<��Bb	4y�΄�n�WlRk��JX(���6!ķ7�}&P"?u��Yz�M��ր^]q˗5�.�ҩ@Lf���c"�:L|�ݕ���qn]f ���ŒJ9M����P��TCyr[�H��L�0�/�낡[5�=@6����[���@��CVS#�
����l�ZM�)��y"j%�3;��莡�y7����x�ʁi�CH��mǨ�e�)	.�L�� 4��ר�m�o��rjK��Hd�q�'l𨫾�)90l��=d�m��/��_²E>��[s�������ʎŜ�.��ݠy�:4���+a�p��e�snE��=^���J�.l�.��Ƈ�{�4���-��ZS�$�U���D�o��.�xZ�¶֪��>��ƅ3�t�6�4�7�d�+Cv�
c>�M{�yloe�Q���ۋ���*�d��� �����:�E�3�j�l��=��놹�"���L�IT�=X�ڑ�n���*�ל��x���6擐ww�v(J�t~�(2{U�O5�Y�҇�v�� ^B������
�����=��6+��z��Gog�#0�$C!m��9 8*�R|�]�G<!���ۓC�������dJw����8�� �=��/�y _yܧq���<��>��&�HT̰�&��ǔ^�����S|�yt!���1y���y�W!�ȟ'�oǇ*X2���GM�����j�-�ok�ˢ����BU�2�Ӓ�y���#.�"����ӆ�'S-%t�(��͍*^FZ�2~��:��7L!|"���.��s�f�������i�%��dY��0��boE�܈���(�gߒ�0�;�e�x���5[j������We1a��%�bq<h��ћiNup�H�36�5�;o�W, 9?���y�q�._��a�=����N~�]@0q���G�OG�(~�	ċO[J����g���?$���S�E��!�51qs��_���>=�3��{�q.x�r�!�Q�Mz<&s��_(�Ɗ���OnV����'A�}u^�]n��>�GH��I��_ɇǵ][��x�zP�T�l}o{g�]�A۞�ɤ��[oXT�̭#�!0�����'!�-m��󠭻���,��%�Nˢ�h\�
���k Ȍ��
���0ҍ-���
'��^�v��	�^7fZ�P���Cy�6��FT��a��D����T�XM�E����߲o�J���T��<�TC�q>:d��Ǒ��#������2�.���)�*����	Q	�opX� [��-C���)cYD9���Q���v4���r��`Jq$��b�^$D�34���9�{ſ/n�;s*�׎ V:?H�p�~��I)��Vز��QM�� ��@���� �5%A����o4Y���jI�Oe��n5Osd�*��:�B�뷿y���A��\x@�phb�gk��=ΘdU�cx�Мy(�6�����I���Yo��]��3���U�"��$A��iI s����b�M�dȋQ�������p]�@��~���DA�D��=j?�(���"����l!vǼ�2�M�O=T�[[-~�|�+I|r����z���%kB���F����,��;T��z�:>!�4=}�5�u�ˁR��|_vG.�Q1�mn�E)����3�@�H�L$Lj������P-��$|�;��P�o�.�x4�%���g���h�}�w��1��6^�n;L�\*ծ�*�,�"�����G�����z7�&LB[U�������tD�;���<��V$b��٭�4d	Y��\yyu|���ꌇ���iv����^���Zs�fH�L��ɸ�+�40��F�Q�Sq
�����jwNj
@c��n�A�Fd��n���bs�:�,�,�z���(��!����O��c��y��-�����J���ک7��� ��c�)i_ j�~��U�ȹ_0��S��F�_�AT4��q���WqL�������d	�)��aV-z7u� �ئ�����r���J
&T+a6 	EK�'(势�~RV0��
�g|_�a(u> pj(�C�'�����������[k�quu��{��ܑ{$@��nҿOA���P$�Y6��+��������%%NB���Bނj�2��+`�"Ӷ%��Y?.���"9,��v�]��&���[M�̓+���y~�u?�pS��H�f*5r����\�(��
uE�&�)�r�l��8!�*�F@R4�L��I����&���IEz/JC#ճ�VK��,}��"������9�&�Ԑ�C�=�\Kg
5�O�*�Pa9�$+*�sn�#Fo�\��me ˼z^�ǵ�u�/�0"�Ȋ.��) ����>7��E�;�
Z�Oc���fSrʣ&JC�h������Yb,��@�f0�Ē6��Z-���^u�X���������<6����l�&�'�Ι�S��9��PȽ�۝険G��v-��q�]Mݿͺ���'uR��鰏G��	� ���o�iP(A����]0��Q����{D���~.aO�/��c�
�
j��$���yb��jqU�hg%�[�t��죍1�G�ϼP�R�{�^̀V)(;������e����w�G��wr��%/R(������#W��b��?��A�5A7��<:��U@�`1����Z���{�80�,q��O��ٝ0f�C�B�X/��~�Z�~\+��Ӛv��z�z3��#����g*��XaH8�Jr�$QźcQ���G�V�L�J��
1��d�I��4�I�m��c�R�Ʀ�"ĹR�Z��cP�7��� D̝n�i��L-�ɥ�#D�V��*�ްrӝ�5��^�  ��:����Nqv�vK'��&�U[��E��:�_H��˛,����u��f���M�����k�;2�g�5�$Jڣ�FF8���C>`�VB�������.��<�1����ǹ���:�RtdU��g�)J9��9����69�_�%�c�,�j���ᙯVd����-\GL��n#3Y�m�[ �$�5�s�������j�47nX�.�"��'E�;.�`�h�BtF4�r�?��$!���{�~�XH�b)a}n$�5�<)|�-y!�
��m�/���hL}�B��4<�wOY�W���эQ3���;��ޒ�#+��[G]߆�%'�|d�����B�k�z��O�_��s�ni�B�4�k�
ևpw�_�atI�۬<ü�IQ��׳{�F�^�ku�=����6A���k���@����S>S	�~�IW|k�cnlo�˱A,P�+EX�f�� E�Ͻ���4�O�f:KLD�\2�&�����f�E r+W�X�%�"u�=4�݌��lv'�;�F�#�2����I����8��_:ݰ��IԹ�\RS�b��c�#	����o�o9�P��o.��e�D�//�$���!��#ܛL�Y�����q��o<5�EM���@9ˏ'<)��T�y|C��a{hV��
�\������ǲ��7(�=�zU��Cn%�Bh�5M1��6kcV9_������'n0�&g�C�qF8&w�\��U;7�`�.��/�P-��?�����J��E�^���u5�|cD~<�^�uN�[�͑�����PC�'��?+J�eOr��mlv/�gmpS/��˟���Ĳ�Ǔ��ɝӖ��S���n����XZ���8̏����K�X��%�vk��bֺNSƄ�V{�{M���;��l�C`��i�T��}ׇ�Jx��xu:e�A���4��9� "�	�Iؿ�KUA�:q]��X���=F�o6��r<��	?;4��(�r"k
si[��޹=�j��e.�/YMS�ʘp!�����z�,�CԸ;�Zk�m����ϫ��g�;Tr5�