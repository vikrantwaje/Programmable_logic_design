LIBRARY ieee;
USE ieee.std_logic_1164.all;

 ENTITY mux_2bit_3to1 IS
 PORT ( S, U, V, W: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 M: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
 );
 END mux_2bit_3to1;
 
 ARCHITECTURE Behavior OF mux_2bit_3to1 IS
 begin
 PROCESS(U,V,W,S)
BEGIN
--S_STATUS<=S;
CASE S IS
WHEN "00"=> M<=U;
WHEN "01"=> M<=V;
WHEN "10"=> M<=W;
WHEN "11"=> M<=W;
WHEN OTHERS=>M<=(OTHERS=>'0');
END CASE;
END PROCESS;
 END Behavior;
 
 LIBRARY ieee;
USE ieee.std_logic_1164.all;
  ENTITY char_7seg IS
 PORT ( C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 Display: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
 );
 END char_7seg;
 
 ARCHITECTURE Behavior OF char_7seg IS
 BEGIN
PROCESS(C)
BEGIN
CASE C IS
WHEN "00"=>DISPLAY<="0100001";
WHEN "01"=>DISPLAY<="0000110";
WHEN "10"=>DISPLAY<="1111001";
WHEN "11"=>DISPLAY<="1111111";
WHEN OTHERS=>DISPLAY<=(OTHERS=>'1');
END CASE;
END PROCESS;
 
 END Behavior;
 
 LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LAB1part5 IS
PORT ( SW: IN STD_LOGIC_VECTOR(9 DOWNTO 0);
LEDR : OUT  STD_LOGIC_VECTOR(9 DOWNTO 0);
HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) ;
HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) 
 

);
END ENTITY LAB1part5;

ARCHITECTURE Behavior OF LAB1part5 IS

COMPONENT mux_2bit_3to1
PORT ( S, U, V, W: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
M: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
);
END COMPONENT;

COMPONENT char_7seg
PORT
 ( 
 C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
 Display: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
 );
 END COMPONENT;
 
 SIGNAL M0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
 SIGNAL M2 : STD_LOGIC_VECTOR(1 DOWNTO 0);

 
 BEGIN
 LEDR(9 downto 8)<=SW(9 DOWNTO 8);
 U0: mux_2bit_3to1 PORT MAP (SW(9 DOWNTO 8), SW(5 DOWNTO 4) ,SW(1 DOWNTO 0),SW(3 DOWNTO 2), M0);
 U1: mux_2bit_3to1 PORT MAP (SW(9 DOWNTO 8),  SW(3 DOWNTO 2),SW(5 DOWNTO 4),SW(1 DOWNTO 0), M1);
 U2: mux_2bit_3to1 PORT MAP (SW(9 DOWNTO 8), SW(1 DOWNTO 0),SW(3 DOWNTO 2),SW(5 DOWNTO 4), M2);
 
 H0: char_7seg PORT MAP (M0, HEX0);
 H1: char_7seg PORT MAP (M1, HEX1);
 H2: char_7seg PORT MAP (M2, HEX2);



 
 END Behavior;
 
