��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#���˕�ɮ!~��'�࿬����G;�BV�e�(`FQn��X+��`������-�5���^�#���m��V�u�`�"��gY'��bP4�~�H�Eʡ��nv��������~t0f'��=��Ċ��:r�1�,�[p*�z�T](�����L���&��q�s�*9�\?��0K�Q��PW\��:�b�،�nH��pB�N�xX�u��'jPB|D�%$iT����ZkZ�o'k�%��͔�SO� ����q�=CƀC� �%���6�~�z�#'�h��V]Ɲ~X<���VGgh ?��ڣģ�L�]m�s�ٗ��/�T��r��t ���,�$����ƥ�[�!�*�?l�%��K�Y,��22y�2ͬ}ћQ)�VřF9��#�Xg�BK|~�ʴվE�%���#8�C�4Nn�ۈ�W�?\�8h�\��ow�#)�� �P��+#<��D5<�H��+v�c���p-�5985�Ebn�7��C���
{�;����"�+�U�fwd�Tw�w�<y�>4Ms�� �qh?�w"d�Kb�`)+���d��x������*M����(��1���oc�dw샴�@����]��2���E��:���̲�D[�����x���e%�^'���7��.��"�e��-�����sKm���̠�x�oO'`J��%Ţ��+�Xp�{d�0��Fr�#��2ҟ�|��,5�G��o����c�2�90�c�����}��/b�*�De�	["oO�_�1��Q/�+F��5��[�:�F���y}�k�;l�1�N2;��ݭ|u$k�"Y��a�T�9���<g�q��0�W3���M��4�ײI�
ϑ�� ��9����r��>p���Ls��D�jC� ��Z���v�]I�K+C�C�5��ѫy%����2��W��uB�����	����T;����+8!������ez�m-"�DVJ�-�._g��{y�1Ka¼#���?+��J�������o"��d�Z<R
�U�?ІK��uX�7p[�R�^0�o#����tHx������zQ�g*L(�r��V$�W4S%cV�PޫKeXk-/���L�j��Z!�|-*sPE=��tv���>A�6-L&k9�2;uQ¶Ԃ�'t3����$����r��-"e/(�1Opi���y�U^�	�G[���Vb��a�G�Q�����XB>z�4#��Zᷳ��:�Lj��k���|H�h��@}�+�ǰ1�@�,�M4�P��z���/t���Ƥ�o^�����T�BL�U�@�o���%+���̎5a��	J���!��gz�DZe����Ƈ�d�A��	[B����z��9tZ/%�'���dq4l{BѲdf���?��ժ�uB8��u"1W�y�|]��7��E�O͎Y�ط�� ���7 �Ȅe,�W~*_ߘ|C�Fx�8�ݫ��K���³�x9��xk��y	W��ނ-��&4!�n~Ӳ����뼓Ϥ��NX�䭼��Ҧ��~1q#�߽mt��R��h~�sF�
�����p~��&�Q�K8yyr�Eퟪ�e��A��4Z��l9^4��&�X������)	-a��
�����*�Co�S�f,�.R��D���.�=}P�s"ĉ$`Y�:g�MS~�C[�,�F�j��]ğn!Fz��������.{�x��oY����R�~ /W��f"阒��[�� `�Bd�qs�Z��"��MC�ʍ����E���N�BA`q-P\n< ����f�� ,z9��Te�8>nG�t=�_����X�*�����t��[�q1���͘��w���ep�(EJ��2���T�/HD���Aw�L�d���H�o�����_H��Jٛ��!S7_�Mr�@�]�S�@���&�C^b������`��V�E��+��x��D��!�n�%w�
p���y~T:k}@�5M����~wW���o���M�<D}�J����\`Qp��~� �k���G��K���e�hs����|�r���<���<C-_���lq�Mm��E�ӸҨ��_v������No�hԃ�櫱�a��h^�sb�aF�j��q��bۋO��'��U�S��8�0z
�W5tR^�	"A�����*FZA��ҙyc���ꅜ����r]Z%� �T�Q��ψ�5Fm1��֣��������YiK<�ad�'� ����So�~�#��{�>1�S�*��I��b���j/�DX��������+Z�H�x8�`h��ꈞ�.�1%�I��I�o�N g	I<�_"3+��m�}�B�Bc�a&47,�j�$-�@�[is�k�ZZw��%� �a��LoO5�jx��m=�.��%D`6R���J�qCHd��Rqu�L��_ (�f�΃<�%���+n�so8G���-��{�(M�+���͋'�>K���}2�L�#L�g�Ǫ��y�r7�|�h��<�^5��<S�>�r*O ��u�[�+��'^ �dC$~oc]I$r�T48���d��rV�]ӓ��C� ���=s�=I�mJ�1��Y��?�)��>��q۲�KAA�e���TΟ��])�9:U*��
$�R��pA�c�q��%�o��,~���i�<�q�� �mգ��*��l�吹�Y�ZR����Xh9�o��5� ��E��f��\����87�^]�~$nN�e�~�16)���E+�4*ʦ_o�>a`]�U�x���Ŷ̓��f�_�x�V��׋+ ��B�xb!Z�F~s���YFV�C�_�rF�R��X΅L��I���9�|o�G�juS~(9��6�/r��f�����L��Ov���$���c <�4:iB�֛�2横��g�e�D�~��*?gI|d�-��x�G`9Mt0w�B|dx3=��q��S�x+���>ߢ��V�[�ח���Y0�{m���f@xAq|�`�S�l��E����cE3�������ƚ7�aiEv����6�TH~|�QҬ�b^�*�AO��������Z}�J2<Q�%uF_�ޟQ�*�rO�0��q��U�'qq����#����G�t��W����y�'�n_?�eSm,�>��� �O�K�䟩�54��F<d4gYe*srLA�%���`9l��b��?����s])VP����0�`��![�P�j�W�
�m�a��c�h8���o@$�?$�wPzB��������W�@i�3�:��g,s�B��X�ϻ{-^"(ӯ��T4l=�@J��v�����33��6��@�~�P���*���&��B|��&žn���%������jPh|' Y� �<�)�M�^x����!���u�v�k�1�6=�����'��Y�� �!��AM1�|���Ur� �����[�^�w����a�@�1F������u�K
Jor���Z2�ۈ�w'#Գ�K�O3�.�Җ����K�x���d�N�C y<����������%�M��D�2�RH��������~ '�Xb��P��^w�`��v�7�:�&b�?!$���
�?W�q���8d��j�Ŋ� �X,�:�9�D��(��������4�C�n�+�+��\�bݐ�Tm��?$��cY�%�kM�]35���*X����	���0bVY��}��G_;�MD�)�v�