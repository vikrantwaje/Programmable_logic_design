��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#��a���p�� ���w�1$4� Pkd̰P�	�{bne�Fv��`V�b���9^Ln��U`�ܜ,�T��W�_2oRPx�A���P���\���4}�pQB��5`���ij�'�z��h����L�v��v
y&&*u/�n+|o�{��c;c<;,��I�ƦhU�H�YmOWB-D��`��:���M�W�P�\��W���W�sV��8h�0gDw�m���"1[Pqgm�iwj�5̚��փl����N�Ap�씂�q�_�������ɚ��%�;|�J�_k׳�PdѰ	g��C(!kD��� "1��.��@����AP�=|t[2J䒳�]3��3�OT|���I�7
�:�O�Y��K�xӦ�$A�LGf���?�Ê0y�����)!?~��c������:H/K�o-U�4�0�Ol3�9YG����ƪD�RTnT��k�@?�x��2�§Vʵ�u���f0HP	2'�T�F�fQNq�.�Y����L�'9=��u
�����5�N7$���:�"�hC���Q	 ���*���6*se���s��~G:��b�?�S9���{�nLD#�3�)��)!kK?�i-Gn�y��]ɐ[��9G����	�n�9����G5F[牔�=SC.+C��S�	�Iw�I��-s�x��
�,�)��B�s_��,��MIQd���y�<�Z�,�w";_ 9�**���~�_7McoF�'�/�$d�����?�7�y���x�*��o�Ouf���.�B�f��*��^��f,��T��tP4/��8%��8�&�.�mӇ��|Q���6u��С\oD��-���Z؉m;��IsUOb��Y/��X���$q��"yM�g�eM�w�(ص�;���
�� �Q�K��b'�r}M$;E�y�B��d�畇��t�- ����δ��;rarg���.�f�2Z���OS�������TaWL ]�8~8y�~�Th��6*�'.�R���#T�'�$h����LnC��x〃�
�~�F�x�"x�"�)7�}�/��J�՟ S-#Q������y���=:f}ֳS|�?E���Ժri��I���ľ�j.���+v��^��?\�%��T��M�l͕�W9Y2ڸTq��u�N���vm�Ч��.�9^����*.F�އ���SS��CR6�Ѹ�`׵ւl&+`��e�Y���;��O�r2��Gn|�(�V[#�e�<|�dq �*ƒb�so"�G���c0�5�wAl$��8��Ze�����GTy!Y��>��r�7���H���@cLY�,��[8�峏��i`���l������p��U{*�����+2�(�
���:g!:�oMd���Pw��P �Kp�q�,�E��P� ��	�oY3`KnS�ӿ�\�:S[Y�$���64�G�+&ؽ4
 �?��*��ꪙJ��(�U
���?=��Cߊ����[=zG�2-+
&�-�
��$��ƶ��KA����\o�-�y�~��r�pfl���I�
&W���l�����+����|@}�ְ�x������ea�fn�����0L�2����חwS���)b#��W�$�R�,9��oO���l%)����W��6�vh�=�}̪��/25Q��;����D�������2��B%U�����*���í�f5@J�
�\U����6��0B��Oe6l���7WK�4]t�B?�;o"��,֥�~M�ВKPQ�[��O��1�����R;�q���j��4���o'wk��x�G�� ќ����0>�I� �?�����MJʙE��Bu���yX�p�K�a�)��B��F3f�p9S a��=gT}��}f���'R6�l��h|k亃ñ���B�?,���9L-�aJ�X�Ԓ&��5d�s����/ �L?��1�[�zɹa�-������п�<��|�+�� [��Ą�/���c�o��l�B��rq���>��>���q���d�Ԩ���ﳊ�9�ج��yOUa�v�Į���2��܂RG�tĩ�z��'s��`��mo�9ϸ�Z1�A9�C���2�h���5�Cv���������Ʀ��B��1Z��aa��m�
�X�Q��eW=���g,?sE�	��(��C�pj&D�Z6A���uf�'nHSad0��� j�\���_1��ZcOi>���^��o��P;�����'���-|��1�/�7b����y�����R�����~��yLϝ{$���� g��Y�d#Y���3hw�GjLqD*����` |M:�h*�S,%K��n�yRw~�Sl�TH=�z�(��*����B�d��� �ʏ�B��a�տ��$<C��Wq��#��L
��XZD6�"�[P����BO�;��|4�3{ �s�M.�Ke1���{;�UI�oW��d������M���
�;G�;B�,�?��v���-3{=T>sh{�)����B�PƄ�5|J'�qK�xi�!�VR�gWz�v4�Q��'��7�d���	�E��2�țuD6�@w¹�z�:�/��'�)�M�"�v�]��������x�s�~�dK����b��N� 7�L�k�9���V���V��~`�}rV'�� �0��UZ�?PY�ݟ`�kݘJ��&�QݒV�WB�;���~�˼b����M�ek�?p�E[��k�З�w�����oN`�Q��L�1X����S��h��a����]�#�@ �?�����I��{:�� ���B!��64��,
>����y������Q;L���Y�Z�O�,5�,���&���3'�߸8P�Ȑ�Dܟ)_��=1�Ȏ��v�i_u$oqB O�쮺������.�������>8���G�gF1o�C�
Ա�G��A�3�p.d�<�#0�$�z�e?Iw��V�Ȱ�"��#i F��PTq�,]�Q[�O������m�E�aK�̣_#�����Y�쾴���}4�yw�W�q9�jv�k�B���ůNV�!�g��jsP���u迀�Z^[��A�XZN���	��("����>�/�f�l�ۦ3�#MfR[���%�H#��:�<o��f�t���pAA�,^�O`3J�w��<��?����yD�[2�{ ���*��@�:�$����TUd�pgEM�f�Rj��{�?Cݏ���kS�lzz������(�3����L��7�jб����ey?N������4�5{��v��N����oD�u}&0�C!����m�-�pG��1