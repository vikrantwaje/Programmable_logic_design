��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#���{��F�ї�,0,���$�a����i/U:w ^ِ�^h�eK�V[P*�w/���/�Mr�4Xː���]Aǐ1?��50" �	?RH@f.�i@-�4	�G��a����S2��
"g�*^�ج�y�K��<�]�����a�0�K�m%1Nn�^S`�)��w�S����K�'��=��M+���<[� �ࡪ�B�tS�1q����P���Ԕ������qŤ��4�E�����|:vZ��=ǅ�9��9џI��+�U X*U.��N��ۤ�l�a¹� �]�3uaܿ���-���������H������Dߊf�W:��ȯ�%c��]AI�(P�y�\�OSt�J �^+��.�-;U��#�}r�P�a"\e]����r�(˂֛V>������lob�������Scg���G�1�N���f�ߪ��vB)�뭚�.\҅��l���0��H=�ƪV�X��l���vL{srTC V��ϛ��1��C�0.�;Y�X�r䋿~�j^���;���	tz�p���v�OZaB+���,�����.I����_׸�a�3+�g�����:\b,К:���% B�/�u���C�V)n"�7fW@L�}��4;������&�c���]�S�9�2������Ow[��	:S���]ۥYn
ǞU����G��6��y�X^h*�y��o�\=X�^z�a���� ��o[�"��s�	�i�L�a�G�޼���7?B�Q��+�5*%ZA�=I����w$�~�<g�C�QO���̰�o��ay����Ur�M�靥�ʘ~�_[��N���&A:�	Y�()�޵8�>yK�`w��X&�UL%�N�E�s�K�w��T";!1���xuA�]�1�8إ,�6�����{�}�6!�A�I*}�r�����Y='
Fo�Y9\!pfic�Z4&h0u�Q��4g<�p� ��Z�<�1��jً�!�x$�ם�7��]%HB�U���KhK���`������9]%��ٜv�e
n{W���:��������]m��X�#��JJǱ6 ��K�\����p������fL6Q2�y�M������c�IK!��<��a�i_T#K< 
���o�9������>׿��Er O
�eּ)�4u����+�&/"V9�B��Y1����=8m�6dI�o��KI�v��K�M����'��>r��?�y�w�������U�q���e�D�:u2H-�m�*���!} LC������yTuX����R�����o߮�Y�B�2`T�����,;0��ț�E�X氛r�Xb,�J�O�����i��KL��d{� U��k>���4��~Fd�$$�b�k�^�D�����2'��rN@m�a�J���l���� ��V,�l78`_;(^`�ԯ�9�
��N�w�`���dC���¡P㹕S*��;1$�1�ApۙA��+)	P7�I�}�ג̞�om��,L�5��Dʑ��%t�͊��/�A�.��:�h��P�ek�_7�O��K��Cܪ�������v>W��D��b����.����0�R�����?�ncD�'�8I}���GB�+��YMɰ�������voWDNXEܟq���״�`�v޻��b����^�v�Uł�ؿ�p���%���[�jGt!G3V��1"hhF����kOڊW+N�v� �O����W]O'�z`(��(K�_�(�/e�}�T1#�uۆ�s�%u�{�)�Gx�m�a�4;���F�a)ô^
a��l��+���*�՝cv�6�i�#Ao�aa��?�jk�S[�Yy'��0�<���L[�&H�d�\s��0���\3�A�my�c�<��|$���m�-Շ�ue����0|TNᦎ1ZTj���!4�(�%�GNiq�tQd�y�T�	�Җ!�;GX}������AB+�G;�ⰺk a�� �{>7ݶ�:C�gXs�Lg��6��%o&Dtt�\���T���ڋC��_Wa��FK�C�֘�p�	����+qD���90��,2ZK����3�Ne0jxV���R1�-\|M�W��J���5Ugh0 ��o=�iۅg,�J�VwZ�/��&�L�Ȯ+OL]S����o����M��>6Ҭ;)H�酉?!�M�E�m�,.e���r9Ikb���	3�)B�w�܉P��
e50�>g�@Z_K4��4Y.�1:O�w)L����Jh���B��c�f��3|(���PC�0G�D�ζȿՈ�DO
N@���nτ��893j�Rw��5���0�3��w�u'n���v�"{���%�����V��uK}>��ܓ�r�D����};i��P	L;��|/�`.Fp+q.$Qذ�úY���F�Rb�Ơ�lf����/�'��P4?���Vn���3f�b�]l��u�tKL� U��<�~��]({�����!�Y�3�?~}�O�Q��^h`�y�mh�w�������f�>�����p5��|�ҽ���V�Ӝ`�[������j��ȯԑ�uX� u3����pl�J�I��KݻY���I=M�m������[�ɍݔ�-D�Rl�J�R�F�"����_�����
�fأN3Y�j��;`�1����`���l��F���ۑ�*__�[�|��1|�2��Y3P�6�Z����.��h�v0�$��wk�
�BF㚾׬�ѐ�o�P2�����q�Q�p<��~5�M�~��� -��K�ݎ,o�x�cp�����s!r�G%�oRնc[�/;�ks�(`���D���7����z��W��lN2�Y��L`޶�Bʟ�DD�Ku�rь�������?�;�������ɴCwx 5��az���U9�?��^X����!)�
�C��x���$9r�h�o�S��Dd�����Yu�p�m�s{��8E�7�:����<���X�=|(��� �_[F��l�KkfN\D�!�� <���9r]6���#��o-G�8�b�\��{sJl�)�s��15�t��º�H{�}�tFgL�g4����Ob��Cj���$��iM�u��4�����Y��b,4��E72�=�us�e��<$c��@X�(!D�^Y��.%B��6�.��3�[״xTy��`sU�r�C'W��)�T�(�eپPƂ�s�e��%��eL� S�����-/m�MT�\�? ��6'ܠ�OXQ�<-�h�	���7�aF�