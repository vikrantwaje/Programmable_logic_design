��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#��a���p� \�M�@m9>{�te1S��_�)>n��:�C�O�$�T�����Dz�/��DAc3 ��,�}-��lr��K*Z��Y&xX|���(*g�;e���φ4�5w��}8g�uj�Y�������9#�w8�u�˽�P`���iBBA�����g@;�H�s>��?y���h��p*I;�-�9�p=L�Ou�Uߒ��e*��ց���G;��-Zb���*|�<��6L^�X�j!��\�<���r�7Ԏ0��n�"'P�����|��� �d��0����\�?���y�WŽ��T����\��-V�W���b����� h�[ևҺF	�(V���7�Rd
�ݛ�T��������n�:��rhq	���}��XwS�����l�mt'mf���RjƑЪ5��(<��F�]�m���|�!�0���3Ny���T^�s�^���Q  )�וʻ<g�+�]�j��T��>�8����jf�_|L�G�u��x�J$��3��u�7����8�ka��iI�t��0z��'��7y�-�Y���W�S���-�5�Eخ�;H�z^�Xi�w�ME#����ZJ=��_!;�W��$���9�P��
�KG'���\��z�[e�@��͎�<�Zl��G���?䖫3ֽ�7�2�3h&՗��
�$��h�x5�О=*{��W;��[�?4�T�#c<�m+0��
cf�?��v�T[u`��A�h�=.ؙ���ı�ΰ0$�Z�h[���U��܇ȷˈ[��f6��])��$�����7����o�v�#�q��%`��u�E��=ɑ�΃K)��1�N9zt�{NpIV�[,/�܋cp�����X�&h�nʡ��>��L*�meV�-�١W��5G�����lN<���!��+-OfԪH�_׶��V��~�-��)Vb���A���ʸ*��Wո��W�ՀP^[�~��Bi� ';t�����8�]8]�Z�A�ʡ�B�7�éOU���c����E����T��B�vY�:�ʹ��	�WU.���6��ʁ���}ތr�G�*�$GP��d1H�@-	��������Al��粩��Ɛt�>�Hk����lO���2+9��
ڄ���1��\hK[z�������t.�M޼g�<�:�s�Q=�Oz�SW����et�l1X!�'u�~C��!�Ŷ�])����kofg�c{vQ��� ����+�S,=�x机�K"�2��E�Ǫ��KP�q�c�8�n��O��v�p���)vԴo~E�߸�� �?�+�a��H�ڿ���*4�w�K���<�xM!o�|)���H���3�Ḏ�џ��ζ���Y��w�8
u
_�u��FjV�=���d�����w�����m'�P%ھ�DG��v�*JH�L��K������9�w�?�T~���Q]��T�;K���ySt%B���ƞq�y;�i���u&#�܆�u��F�R�uq&�I����#��5[3uF�����F
�i�>_�s�{���?U���w�^�l(����T�Bx�K���с�I1����MM�c��T�H��A�����r#!�N��D�]�́�QA�����?
�,Df����'��q��>�1�����~{R���.}���C�����i�C�گ8{�ֺ���,��{ ��lس��X��8�jگ��8e�多�zd��7��'t�y��3�S ́�#,��Qk �΀�4ӏT���:�W��#X�i��D�;�RPB�èz�e�+3dB	z�ŗs$���QڦUCL�*bS%;bNB*E�hDpB*3nu4�y��^:i��>�m�:�ΑbE�	ͳt�5q�c�눒�ƶR7,��
>ʵ��T�2��ʇ9�u������kz������m�퀛�8��l�O���P��ΕH�HFU����MF-W��7�.#���.Q���8k��3�ߑ�	1)hQ��_�W�C�Hc.�0{�/bd�w?dp[M�׉9����
������EBD!^ĩ������3O%���SӵB� �%�24�ک�������o���S���a�dh��X��`���43?�w�I�"����O�h���2b���,� ���2�� i-׌s6�W;^�y���g!��Ґc�/�%@��	�Cm��F�|�&\8N�+���HUo�w�Z����� �h����qؐ
>�eu�u�!3;��/�>=v�@�OU���Z������ D�������:T���,�� R����}����b'�d	��d�����H��}O���|Z�ϿR;�=�YQ%M�	_��,�sF_+�^u^�������Iq�7�A*8l�5���n����%Ň���L�.��-���C�o>�ș'�aw�Q�I�Dx궲�]3*���h�u��+��]y?\��W��9s 6sr��ݚ��T]i�@���ބ�M+��W���<}^�)��|]c���~2��[ �4"WX�3se�:���0GN0gY�}��)�����$h�{�����Z�`>�|�j]�_��4ޤI6��n�����b4>�����&~u܂F%r+a-���Q�A5߁�!CMM(G/?�ϊؿ�l�'�.��9^VF}u����ҪmF?FƲ��H�AQ�'���^Ʒ��$���90LǙ]pQ� E5[��Cx���� 0��$s�ă��?@����~���~�?��v�4����a���ӽ,c�z!w���j�Sr2�!�3�p�+l�/>�n��@j����Zi�e��	`+��:uy����	Ec�!7�`'�)�j0��\�f6��##��<���Zp�n�YO�1���H6��+~�sL�Mh�͹����!���L �l�Ԍ���`��D$�&�����o뺩d������Cd��@`iY��3�oo�jN%��wƏ�I̬��o��f�����I����`��·1������=�����N"��}YW+ǽ��C�Ʈ$���{6����l���?	Y��_�r��p�o�jz����OJ#�ǆ������ve�f�=��bIv�0ɃZy�)4�V�i�s���0�/�,	.9��l4�rU�8�V�y���}E�*	��V34��XYRgs�-��`�ē��及�!w��x��\-����a�	�f��B�Z�G��*�Q/�@���wN�x�:�6Ju,����yO�,����`��."��BߤM_���� ��FF��<����t��ڣ�R�9e�cec��U����hy����Aw�e�^�q���3:�~�OM^��l�3A?z�/�F\��d���@Bw��*�ˣO:�&N�V��h�P�ȘA��� (�J�2�lR9�Yi�~Hz���(��}F_��ee�������N�IR�r�g|��[��r��W݊�j��
7�-�'@4���d��ѐgd��f��m�
���܊>�~���_��"�]�@8w�/V{?������Y|h�ǢӬ0\��|p%D�����'��Ж	s�e˝��u�q˴jn��E��O$�v�5f��_y`���Ai
|�^.�܎=��5�}�{�ip��R,S�������O��a�X
2)
K�"e8at�{ͳ����Q}q����:И�)�y#c�&�P5�~|7y6T�_�/�.�숄���S���q��byť���߮N&v%a�֦S7��.m|�%��<��	�e$�x�P.����g�3��嘆�t�"�u�[	DL� ��`�w��~�9��K*�;��\*Ҙ0��M�Q�Z��A4t�`���	b�0~�K:o�(�k6b�M��x�ڑ�V<��fFm��~1X���쉛�Q�I�u��L�]����f���}�_���_e~��ww�]�q�	X����I�	>nq&n(}��ͱn��Q_�ՆY_fA ���Ħp��F�"X�"6�;�p������?����pרUX�-yс�Vo�o ?���Y�'n�ԓ�3�Ak��_�Sf�K��c��ʼJ�?	(�����?ޡJ������
~}��0}5��J��!��e�R�s�j}��Y�,��
�"/K���{�bCk?�8� ���5���ra~;�,���B@S�
n���I�[�^��j��C�/�26a֭�Kn#����|é �
7�΄��s�����޷��ӈ��_�	�X�(~������!Jk�U���jo�{%IN}���Ce@ٶV�-�^s��e�$��w� }ӑ�����cj�3���� Û�z�(��ّH�d�� #�8n��ݍ����a��ϰ�bz0iW�*7����(�x[���`-�H.|$�H�zT�ڧT�JZ5DX��Sl����r��q�1���=�h
Q����>��D��j/��&�K������652`��E��y�Pw)��X�:}�V
2'd��uk�����4y�hT�g[׮-�{.M%���z54:�.
�����.�X�%%��%�~�j>[$'��3�Lkf�V1�h _��,��)�����q�P�m΋o0g���5fG0����e{��7h�w.�� ��\9Η;ҖX}L_ :��#����J(������1���xߥ�Y�1=�΃�3D�Nܹ�iP鵶�?K	�C��^Qz��8x�:������&�(�a��d��T�#����T`WRֵ4�P�E<�V«JtXv����o��o�v��&���`�� ��J�y��\���zT��b����P�*zF��]uzQ=�кX���g����GC�B�F�����>[�T����L�$UWA��*����b����R(���/_�ȏݻY��A��&G�۸2/�΋��3���mIPlך���i�\�np�:*�6h���7A:94_s�$CX9�Ϟ���ũ���%����Mz��.��%���V��uw�m�˶nIF�Z���;Z5��"v��Rn#"�MS�5��B�ןe	,���������d��'�m�o����gZ&Q�uFx*�뚇D"h�YE�;Q~�ED��?y�����J&(agD�ݰ	Q��X(��?�VL��ͺ�7��k�u�Y*o��֘{���i�٩�ٞ	X���09�{�!����UB>��N��T��kⳣ4�"�,w���=�Q|�BTz���A���s�����&�&h$�>�i��,�t��!˲r�?3�	_���œV6}8�
�O�{�kacC3uxq���jIn���l�����)��B��}��Z��E#?EVx��'�}���2\�it������$l����a�*d�[���S�_p֜�Q"��"��ʢC��l?SC�s����i�q��I����=�.�F�v�G�9�����i�C@+�9�wJw�&�q��s�7�>Ջ��Gy�7h��9>���j�����Q�T!)��Jw���tBm�8y�ȇ�s(t���/> "���lO�͚݋oȎ�r�y�?x�Ta6��i�u8=tՐw'�0��-�I�U�z�r[E�fL� ��t��:��̴�{��4qV9��gK������x�Ie���Q��9�O���mVEf�j��	��HzB�X6�v��+�Z���!e������K@e'��PF���2������5`gɆ����6�b��l�Ǝk@HN4�!Ia>�ؙ@c�B1ne9����Ob U����)���ޗ��|-�w���O������ [�]����0�e:(�Ȋp�#?��j�J5�?�K9�(̊���|,���W_��<k�9�Z�D�V��MSz�l����0ME�&fo�.Vى	{�d�)jr��Om˵}�m���������2f�{�Qn�C%M������A��mH���� 	�׉WuJb�9��_%����?��n����	�hDH�ψNKJ\�Vj�鬔Ճ�3�TZ�i�~�]x$�a�S�c�b/�4 �G�QFsW���m6%1񼀾!������S��> �?L����*c=q�,C	 % �Q̤r?oh�C�����=*}3�3�(�Bsݻ��1����Ã[�4��M�b.��G'��h�z���E�1� ���9�v<,��7{u2���wH��� �/QD,�G	���xhFk���� 
uQ�����g�z��G��;	4��]���#˵
а�"g��c�X3���<kD]{��k�G��9`?�.c����J��݌�
_�"�l�ot=ns*�`m��lUC~��͜��m=2�mEj�f/����]v�LӘSB��5D��?d���%Q���R��x2 :aa	��z4�T��S]�g�/��X���(���j��Pu���`@��f(Ғ� v��;�V��* \좣�k	�� �z8����PG�	��-i��2���9,*���@/����3��A
��]������N���7���2��$����W�\���`�k�r�D'݁�eCι�Ͻ��y�$0�)(S�w�h�	��Q�&����b����y>(J���m�	�_lG&F�Jb��yG�1���Gy/�Q=�iM�N�]��<�JF��	����[�DŲ���'�L�u�BDoW(v:<����;���i�	��*�h�IK�<�c�/�̀�T	mBQc7 ����2�[�Ӎ�[��bx{��mmm��?Ӵ�DJ{(��E������6��< �޶W0�j(�����ߘj�3�>�o��ռݣ4�Y�*�6���qL�Bu<�����������%��)�zm�!p����D� br�%�ܫkz 5�u%K��ǀi�S�J�r9�>8�������kk��5-�n�h�N�+�H ;� 86��|�u�_NE¡�m�e|���>8�7Z�2�	9�7��?~�P��W6��rl'儡| ��֮�������~��B3C��%��8�+��K�#� �a�K=�
��".�MBD ��,��q��(�kg
u����?vX���h�C/���"ɜ�ɋH#��=e�����V���_<=��d\�Z�k�@~J�� >m�����!��*���9| P:J	z�0��j����`(��?��t�+�6����j�� �xa�}'���If�d�G�!�.N�rL�ԙԯ's��=�`���X�����\o;ߧ[ʾ{&���T.efo�ѓn��ZCk_�mw	�ǖeN�*����Cj)i߾�7����;>��۷������q!D7+ ��1��kS��`�E�:L��B~<��o� �0�2����w#��[YK)�z�td�$т�q�#	��SKzZ�l�j�{�A��9��ye 8��*�y�Q:H!)�D*��4�6��%�O���Wo��V
���({�q�I%'8�V���Z�{�e��/�0vΥ�!�s�d�:V.��5Y�U̎�u�F����E K������W�7�
�C�ܺJ�R��_T�M�X��v�:��W2];��Jql(�K�mu�v�j��r4f5�V�jm�](7�#J�}� �\nm8���u�����u%����1 Z�/�3?f	�0�,_m��)Ђ�� F�%n�8�����Լi4��U7������e&��@i��]@$h֬��:�e�w�\qv%����Z���"����������r8��!����c�bϯ���R�p��3ܷ+�_=�Jn����^�����=�m��m�3��w��C�,�qݱ{O�T�)^���(���.�-���P:�F��?:�+_��x��֭*�&��K`�-9A����;�r_�F`t<���t��i���k��tw��H#9ց���0�����&d��B��G�Ű)���Gf֠�.-ӤO�V;p=�	>�^EoyS����v�!�V)�|�dnDB<�.�pt���M��΅�X�x.�H���>����2"6+���_�@<6�=*�2Z)[�$/v?��C�N]?��lHYV��t�_'������c����z)�O�ݶ�Ⱦ��`�b�>!D>T�Stة�-�y9��߆��`u���'^Y��c��I�����o���R*L��ژ�:s���o[N�"�A�m3X3�s^sgGt
k2�h<�L��b[��)�9 �`�� �͉.
�GCPN��1ߞq%w�p�un��
�J�\Z�

����}���8�kX?^���n?af����0�����w�������tR�O���u|��
~���Be���Jy�:�y�:2�<Ɉ��ͱڠ�:�=ǎ����M��_�lΛd�7U]�)G���I�,U&����W�ڽ:g�E+K���GEx�۸M��|q���<�]p�.*~@A�5̳-��\/������(f��Mq/�6�ͳ����O�SY0�EG��u���`����~b>�$��z��%i|[����C�����Q���zo^�LJ�� Ϙ#���
�s2�`+������<s�-�)�*Rի�Ҷ_��<Yjn������.%y�����[�&�
�IWY��vi�p5%<l�*	�-��`:5rT)w�n�r?s9���@��5&g������=>`�,O��0~*^ab�Q��=h�0�s6}O�5չ"����<y�{?���x�ԅ��w����i�Ll���ȷr�� -Sh璒M��Z�u��{�Gx*15T8�����E��]��M5����b56d����2a��h��@Q��
=<�%kQ��R3�p}S�0=~�VÁ��`�M�ZFn�|X��Q���DTWR���u��nr??��n�;K�6�&@�tˢy0Q;�%�F�>�Z����ʇ� ��$�*�"cq4����-V�� ��O�ph��^��K����^�j4􁦩�\�~������<Yo[!q@����3�2�J4� �׵Ʋ��퓬��=F�@�~���Բk�����ӣr��71�:�o	nD9קG�B' &L�΋��)�9�����yUU��z%~n�W��⋫+�&A�H��N����=�?�KhZ	J����?�����E�N�@P��Eo�W�z��hǫ����YA��o��O_n9�4Q��j���91���;;���֍���/	���r�_��H�e�zCd�7�xN;��&h~R�RC�C$���Q=��K������Ԝh>���3P���R ���_ve~�Yn^�t����+{��8�efX��}�V�#�=.ޟ��cw�zXAN]��P�30)Ԣ�z8������/<�&� ���U�~�R#�3x+��
_�VR�y���@?,�4/��*�De�\��j56�������A�������4�H�|/���4O��Z,prI�Ma��	/'���.;L���A0�&�W�AeC����k��A�|��ۯ�]�g�FT�(�`��>�zB�4?�_��\�x�=�h�>��P��V�ܐx�+�A���f�s��%�,{�{":^��a-�W�5��EvB���L��>-^k�3.E�S�26�I�����&)�H]���~�w�]�z�A`���'�=^�J�_�o�ײ��⑾��p� �8�l K�]���B�Np�Ӝ����]��Y��M+�r'���L����$7N�L�`��>ZĈYd���F
�F#���p~�%�}�����:�*їU�8�lb�8��NzX�67�X�$��g��zТ�[���pM
�Z��o&R�m>~�Anu�-p���gwX�>�S�~G���Vj��R���A���4��Z�����ϗ���,ӧ����Sk�댤0H��f�_�Z��f����c�{�
���%�y�J�@��t�ō��/)�?*�v`[�?�;�cJ�i�����$���B���N>
�M��V����̞���\�*�5��c���Mx�)��(P��ٱj>��#��:s,��n�wT����r/~�򵎢.���W'��� ���Ӌ�6+�/L���@O8�< �� �$?V��E%�k�w%��a��c.����;�����Ѯ$E�����+�=ds�)Dr?���Ss�K�V�`ⱸ\����C4�8{�),\�w���N̢	'⎁����v�p�:y�,sR<����zu����τ�'������r��#�ޓ�E4l�6�:n�̡�J�y��K)�~%=�ԙ�ɔ�!�̡�Q���M�$I�uL�Q�9Q8B���'D���S�����Z�X)��������V@�Ī��`K�?�ΒŖ��y�K�`�sh5#����2��#����=�״�Ԇ+_#ZC9P�����ɢ%��: RNws>���k)I���ߎ�
�o_�~���9�q�a������?�yB���S�R�Ӥ#�ϻ7ФԽ��T����X�K�Zk=�C���,���T�Gd}����I����#ѧ*}�7�A��Թ��w���<�Z𖓾�a�����ԅ����7�j�k����+�YH�?�) ��rv �,�?1u�Kp�E��VB���Gд_ޤ@A�)J-�����b\rT"��L:���	�����_n���#tZ�L�@��0���V;?�XZn������ccڵз���ִ�����!:n���˺�ѓ@jj2�C'��U���p�M���7[{Am�ź�*��_k��_<Up-�>��6�Eb���!東^�� �.�iĔS����q5ȑK`!�,Wc�d��B!D ��}v]�.I��F����Auup�"�����
���X6؃M�sѮF��1�}���5n*�V$�\��ۜ��`vt:�*��_Q����r7��'WS�<{?��d�i�U��ReBWHv�Ӟ���eu1�����?��
�
�f