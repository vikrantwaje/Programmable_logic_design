��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&�8(�; #�4#����%CR����ξ���tJ�$9[�(L�lϖW1�8e�O���9�Np��!hJ��j��þ��j驵�)��eBh�^�m��,��0!듍{��i4gXy�\z�)ݕs�b�����?��C���h��Ky�R��}������g�զ��B_��O���x��Z���s��(>��-${��H�+h������K΃mPͦ�H���\O��GE��I]_�-��`.���%bl��7q��E�b���D���'���e#f�B>�k�#4B�J��f�����2��
�8�-*�|�������~��&�yN��!Yн��0W�GE����>ӊ�-S7���"�*B��/S��s���B1���X���ʔz"W䙚a�ctZE��N��#G�����<�Y��!���	giY�%���/3���z�veGw��z5�'�W9�3���xH�Ysc�L�ɶ�w��p��|�o�+j}��W�l4�����!�d�����4$��N�.{~��>ӗ� 
7>��0��ǘ�u��aN�٢���|�e�DN�ܶJ ~j۲K� ��R�dg���PI�2�2T���ПY��,IW�Nl�ԱB�.���m7��Y	� �1Gb���д#ln�L�mܿ��ݫB7E�Ϧ!������UJ�8�fL��U��>���L�&�	aq��������sR�x�*�4�i݆�33�Ny<��{�R���k���>��n�{Fv���{l�����4�!�B����u���"�P��e����j�a����XF0mW௫�V��Aaz32�|+�J!���.i�U��/�]��>��<���Y��K���^�Ԕ��b3�����|)jBm�!��I� v�.�ӛE{��k��J��{��$�ϭ�%V���˓����L���|뎜E�*�?m�8"��~�|kP�' ��h[Nl���~�r���u���k����J���'Tj�^|����(v�����_�Q����ƹ�-��'dd*�������@#;؇�`w�����'�{Ѹa?�4js���E�Ւ
�67j[�S�M]O?�4��#�3���B��Ǒ��<��s�!��Q��ґ�A�#�������0�w���a����P{y���5f�� �8�3�0��\��պ������>�z:����EY�K��TI��w'}勶1Z^����N�������p�����D�o�H����aP��)�|�Ч��b@��Po�Z�=~Ʃ�5������aÂ��{������D1@��1����0�j��U��Õ��$�k���>���A��m�֬U�ߪ�@S�t^�P�/��.��z�Ŕn�j6JTR��U3ύ���sw;�)��E ��_847��U��ަ��FK�'a��%[s��=�����YLl)E�K+|W?m��+ę���o�ә�h�h2�x[���d���1M3�i�R�iʥmhyDVn�|z"����zT�]

�;����@��n+�����V�}[]+.�u��G����T�|�1�ֵFuRޓc���c�L.�$�ݸ����2�]"���qW�]�d�}FT���6����< td�B��je]��mw|Ώp?bI���\zo��i0�7�FH�?_�,K��(+�W����=�W�%�0�_#�(��;�Φ�������0��-�[���XP�?�+v!2�7����U�+a����q��e��!*����vl��0���W.�6A<B����>���Qj>7=-�TD;ڇ�-,�3���va����Z�XG��"͢V���]N�<an�T�g��%�U�@��|�sϳ�L�;ܶ|�����Ν�\B���ܟ�t�s%Q�R�^5�Y?����l;t��kG
M�\���t�B�F�e+B��
�M�j�2}5i[-�w5	���'���}�`e�<\�'�StՕ������],myk���>3l�\��0��s8Ę�̀�b���1`T�pf�t�Ak�F���L'��G(�: 1 �T*&#qs���{���L��%/m7���/�+(t�@�I�'��/����l(��k<3rH��2>�#U(�pvy3?�'����Dq
\� �Әmֱ����-�����Ǖ&'��h�I�@�P�nk��_Q8��Ƒ2`K�5������j�9�&9d�������گu��D��3<��r�*���;��� Ǒp.�(���
T��śj��!_�O�T���O�ay�I�^�'�܄4&^o�����}����=]�� ��ʍ�ҫ�)����cu�b��� �J���;fkPZ��lOK�v4�B�7�E���]��8��Y����6w%wڿ[�B��v�T��!w�cW�O.d��_�Ϊ�>I�Lu���֓�JhK��6�����W����7.��I�afp1\b*�W��2�.�U��(�����!��nڼ�8t�qJ�#�H0���ŋYɝ˩�SM��6�L``m�:E��p
�e��ժ��W�Fi��I��[,O����c�D����κ�th����Թ:�߼��ڈ2���[��T��Ǐi�0����I����0��6��!^�DD]��:�,���6̥�n�D:�Z5ݔ
j���+�
�"5`��'�Z�ķGy?�ڂ��<��s�ZCY+0,���>�f��L-��/��i�[=�뿩뙦�����;׼�;Z��3b��e����=P�n�+NC�jiq��pgؽVL�N�����V���x�vVU2F	�\�#�)$x#�<_���`[�� _�)�K9����o2����Q��*��%�u��,�i��`@8Ҍ�|��e�{�"�F�2��Ezm��ϱ�r%X�ഢX��L�aDs�����G��h̊?K�� �u�#q�X"rY��)�����0i��W��><�q�!��q<���5b�H�H
��M�r
o�i������N]��Y,;z�ّT�m��8oC#�)�6oP��������iV8�F7���t�Te��������Sl���R��I�������K�Ś�����,�ݦ�E|�"���rg*���������b����\�O��h�/�QM�
����u�x����I�\�- ޕv�nc��c���}��J!�s'Ve8=RY
jA��`�zg(�-/��I��︋ĥxV��3X����:�;���c:�?��q߾$O�+}�BN�{��`
��Q�X�,�&dy�󅏘��n@�14���ClK'e�k!?P���K�]���Cu��a2�2u���GWF�(x�Ҋ{S%SF/)��������<��ż����ue�4n��:j�{��D�B:�t�<� �Qk[���Ә�wZ|7�����p�}�jn�b�Oœ|uc�tL`G�y���}���@�@��Uи��bG�4N#�E��ȃ��$TgHuf��HP���B1�c�"�[!4�
O2�:�R���Սs��Bd��~?��׼�ƨ�q��#�|̎��j�~b�~���r�:�B���*E���I�u���NNO�~��H�-�	�D�E�x�sF~Z��2ƨ�v�}��-�-�17�Y��~��<��A/��y`��L�NR:җݦ�)�W�a��(���"T]����ٴ[m�����V:o�����U7��¿B'mY��ߔ"8��z<�$1����2 ����u�jg�MQ_���W]��,�59@���|�v�����v��+v�k��'��林>]�f"������Ψi�2QF��Ƀ�"��o���1㱤��S.���X�Q�y�D1�Ga0�|��e�g�����E�M�Uњ�'�Z㜻���,8K���N�e-:&=\+���� x��t��{��'��r�Fκ<t��HRiW���������u~�p���u�Z�7��z�Pw� �� ��R��щy(툣K-/���BsLZޕ�I��A�`�DJ��3�y~�`����;^��Q��2�½z�2T�bގ׆Z��f���Ό�3y��B9ɒ���u, �񷛩�F"T��s.�-���2	��rF����6 �ɹϢ;ں�B���>k�5���X�!Aߕٶ���	�A�Ҁ�9k���g���D�8^aU�!P-۠�j��Ek��,]��{���E��2��r/�bQ�:QN���ek�<4N,��L����tD*#M� �YڅE��Ѡ�KH6ĿF
���ne����e�:@5���b;�d�1�f&8\����v�OJUC��T_�i��B�c:�X)y�uv� �e�r �\�r���o@%7������b�����,x<�[�9���2/_H����~*n���	M,�\o�\t��|!��!��J���s|}�vJ'���.Rg*��{�m��%�퍯�OA䃛bH�M��,q"|�"�]�1W�?�P?�X����.�л)��0�a��p��k����<�:�d,
��%���J3�\sEy�$�����:�'f��,ׂ,]i�����b��Ǚ.!c	�¥ʔ�ο]���?J=_�O�|�&�NZSʒXS�4�n�bߓ�g1��e$IJP�s�<��-�t�(*�w��j�>~�]d$oO�t���0)�܈"Mw���,c<d�K�&�X�]�ؔt��J�@o��ǱĔ�UO�T�TeV���Ȇ�p|��&k�/^�ʈ<��(�,�jT\'��3�G��{M�����:
�c�s΍.w|*xyT=�s&�r��_�m���=ei~��5�X����Й���p��t��w��;O p�pxx4>g�J�ﺤ��J`F��b0�`��YFe�l/�7~�����wdES|��[�n�ip��1f�N��ȸ�}�_��6zK�H����fx�X�����&G�茳�l>�R?K/�D����M��HZd�Lۻ�?�;��ą0Zh��1h";M�^!��;��;�t���p2x[zӉ9V����p�S}�4i�i7k�cY���
�7��A �p>E�b��KR�SL�lS���Tόkc͢�����3���y		+�?��yx�zNV칊���F�X��',���mzgw\E�C�����@̧/<�V�?�C&p3��v���*Xz+T�ک��c�!���亮!f�G����Z$?;fU'܉*��f	���Y�Ij��1J4�KtnW�1�9�%X-����}X��SYýV��#9���;y�ͤ�e�9+h�Q#���6&9Ӫ��3bt��ʜ��-�X T�h�>�����L��D�×wv�^1��Ec�GNo��gV@`?� F[Q�9l��Y��sC����n�\`��65)����I�ͤS������� ��Vl�I}����o�5�70,�o�͋�����ډ ^���j�N6H8���H���o�qφS_���ʎ4�(����� ^��7�AiF|�ËRS��_/�A:�U���;d5*���G���T��j02/���(X��74m\wZ؜@�!�B�J�s�������P��yq�v1X�<��֢��/��/;=�-z�����L�B�̨��6�X��3Я<�IY+铰`����%�T���-OF���x���
�O��~�z��M�e7_ΐ̏0��R�m\NN�1�����|se֍��%�M�g���K����@�H�Zx�l_�'�=�|̮c���i�U}�	�'�5t;.�	ב'4.xo��0���a�}��V�S�*<x�3�p�?�l�905FۀY�>�Qg.�<t?3���-�e���%��ԓI���e��'�̋�9f�*��Xh�����^'�7���\�mͪ�����۩շ�:D�Ǹ�W�"��Z��G$�a�� r�g�j�:Owa��R�a���Y������Imz�J-]��O�2��������z�{l��5����~�0�����-�ac ��ntU�Y�����0�~� �O��)
�+��qEI��y�f�*Ja�a��-##3T�2�L��%���٣6<��╭���+�2�w��lI�Y���r����y�|��Ii��vKLf�z<P�B��J���GmD&�?7�4t��\���T��#|Rk&�s�\�br��f�x+��'`9������&)�0��	�P	�r�6���Z�9xdΏ�%*���&��^
3:���gr{؊Z�L�sPL M�;3��H����Jӈ4s��a��R�?�o������Q'��W[bL}�@���1�G�m�0C^W����J�
�9��ʭЊ�+�A ��э��� ���G;Z)�w��:l��c�{��[8pH�&V*}�(UI�w;�U��s���E[� ��͎��,��)�ayw���xsJ䐛6�2>W��\El�B9��E���[��,���L�R�P1*��ֶt���(1gW7���j��w�]d��M^�6{�ޱYn�S7�]�Ng���4��y��L��1�\�+q+�6Y�E3l���>�Ο7a�h$ �CC^�"���>k��% �i6���H����b=��+�w*�~v�t)�`�q�c������+63�_�5��3yɺZ��e���1k�Zdg���u���56z}�ے��_��`M�&����aɩo}u���r�B�6�K8X=�H�MtDݨ㼠9���ܬ�2Z��KdM����������ˊn�F�Lz�_��ߌ���X��bE����%.6�ٞ���宬"� ��B�>��t߂[��Q���s �Y94@��;T���X�E��D���֏OH4�㦅�ȸ�ye�D�P�p����K�~��^(��1:P>�-�ƈ���0�%�K��?Q�_I�K>��|��d_��VX;�3>w���ǸE�3�y�zH�7Ө2����T{$e� �t2@�sD^N�:�ӴM�B����7�Jaq��/:������|�
&�61�  � ���v�+���H���������g�8U�|8|W�9�|L��-6F�^H~��G!�7Jt��v������h5�� ٗ�2�eF�"���Ϝ��(ly�4J ڗ]+ 3��$��Sp���O囯��~j
�S���A�+m�D\<sV�%Ư�>t����@֣�Iw�,ZB��������4$��;|�֤;����AY��e��xh�QB�Ǿ?�J�w�=��ڠm�=��ܯ�oNQm:ʊe J�8�O��ɜ<�z��	��iY}�*g�Og���ͳ�+1������sB����� �9��$HMTnr�˫���μ���zt�"DR?D^d\$s�8P���/8�����5��yȁ+��^f���|����"��&85�Ci��tp���M1�v�/�k�4� ����,����Ɉ"�o�~#�no1(���PԙE7[(&#r����I,x�����GA#\00�RQ�Yo��(�9��V> ���sM�އ�5�d-P���Ҷd��l4-g]�3ecM��`M����������ǘ�_o̥+l���OOE�L����?��>�F'�r��X�b�e�͗ �<
4;�����ʡB
����F�p]�����#�U�A*��ᆂ~'h7�(��cqn t�(���
��*\�w���|�И�\���~�� Tw��k	���H��735D�	xF��aZ�zߺ��m)Fq}�"4:8��d�W��R��/� |0�-��L�G����d�|�>Ow�ub��G^>�GU�R%��s7������cq�"��'P&	��G'��������blTthj<�!i xs�KU^�K*Υ�V���uu�GaCi�V��
Q����<A�F@]�����1�9��G����Ww�Ab��w�=�y	E���"���;	������b��+CD�	��g+���Qགht�h�P����1�ǒ�4��sK�>oo�ӑ��_#n󔫤C��"!�=O�SWՃ����V|���f���9w�ʬ;�j��I�1D�~H�a�����4��}q��l���Xjޱ��$�d�(�ς���27���{�m��3�!��}x]����G7,��m:�I1����d���s��DO����G� ��2α?L��1+�1�̚q��̜
�א��QО[44�6���+RsU�A�n�υ)�wC��T�/,27���7���3���_O��X�=��D��n��V:�Lk�Wy:|���q�� MQ������r��9 ^"����CB�i�XޣCuV6[�W�4�oť Hɳ�\Jɶ̹c��'2⫚��[x�;���J�>Yo���T��麄Ā����(T��k��ړ�gɲ����l�����]Е|O�/J{H���'�Dt�t���»��Cכ����c�H�Pg�a<���O�#6\�Cu]fӜ,��O���m�/t{�a��a��L���H��4ꇮ�zR�T$)<����(bb�����P��>��6�4ą�4}�������^��b�z��>�ѡ��=�φ�k1{��⃖e�ɼк�od_���B��l�skS'�OO�;۰�I�KGy#^�|Ԫp�a�S�q��<SIV�X��ne�T�&�bzX�
��5UX��,�v�/�z%�_�(��I����W"�H
����6���(c8[N�BF���lj�ә��+��*��l
�����[��a���M��r�sv�ދDǷ���cW����ĸ�3����17�kEg�%�	��ޛ�)��_c�ՎY3���	��WԽ��qK�=Q���	D�:�Y��x�0aC_���ن^��<���|�����GKs��cx9�%��g�].l�;Q�u��ʧ�km��a�vX�+I��S(�5���Ժ�{�C%���l-Q�7��=�y!����w�����Ӭ����]���a�
s�DO�ӛ�]�����X*�\�3��@Z-�m�����<�=d!�0��+����pV�K[6d3���(�u'�0�B��W6��Q�����h����l/��a�k� �X�u0�7�ؔ���X��cu{|tf��)+���� �,p_�|/e�x�����iܶ;�N��N��Hr88@�M�F��@��J)�4r�ǔ;����S���F&���; X��
���F���j@X?���}���Z���l)�>~���)����4�?�q
����1��lCQ����MM p��d�flh�14@��*fk��6&�y4����),[̭Q0d�[L�C��س�P ���ְ�)U���\w*�ݩ]]�r��;��w,�i��I�{�	#`�u�@��(
�b
 M�	�R)��	9ǻWÈ�W/� k
����Im��w��-�C�}�zx@U�y%}�Mu^p3����5��+�3����& ����"�G).�4�`�ިɲ��ʸڙ@#u-�a?��lu����s����NMnV�5i�}NL�Qں=���ٔ�~�mR�/Z�T�{u��v���R+��]���5�L����{��{��.����U��u�#�+U����
�����s]��r@5�Z�l�g��-#��°J�J�Gˢֈ�E.\-x%x}v��O���f���H$�n8�$I"̱Qˢ�{��4/2�}��C�F<2}̢@Y�zz��ݬ�	|ڋYU�e�IO�f���Q�X�R�>����[�I[O%��9��D�\�Q������;�]��΀4Y�O�KD$�K8�?i͐:���V�+�����$y�<�؟jj݊�y;X���,�}U��(`��Z�#�!6� �rl�F'�0�f�,C��a��:��*�I����:r^A;��
�A�>{}xB�쳇4��@'0{"�<5��rMSꑣ7փ�.5��"�;��1ty/��0A�E�P+��Noa1dw�q~D� ��c�=%����Y���[��@�$J�<kq�;~H�Z�R��h��~0�դc=`ܛN�ͼ2������y�\�y�T��J!���9��'.W�'�*�����Е'S����rP_�0Q�;L�[VT0���u�H�s8�c��H�(k�in��
�P��y�fX`0����NΚ/� C��L�$��e�p~���E[��X]Q�<�L냳E�M�Bf�ۨz�o�äEƞeQ%9��<�a��f9y�F�P��F�z��z��O�q\���־�%�;U�� �k��MeSv��//<5K�γ��I`2չ�G�	ҵ�h�b᧯��=G�\)ݧD:u�������O]�{���OP�!�Rșu���y�f�*���I���N���-ԅ���t͞�"����F1|	�=��?o";��Nh:�f�<ú|u�̼�$�Y���2=>x�a�'r���O�-	�<p��=9Ƹ:\�ihՓ�+v��Wg�N�h���

fvp��{��|�Ct���3��HIW���lu߷�Ӹ�+{�)И�N���!��0FH�
(V�ޔD%�����l�M����׍���
K��ȷ�d��-�a�c�/�e�Ms��܎�V��yۓ�2�kƬ�A:t�Zhq�L]Dnǋ�oX�GI��ӌOi�$�R~�P3��3�Fꎭ�g�?�~47�Q��R���`����Trf����
���ZKr����.����k��w׋c���S�YË��W�8=�!R�K4M����W�����q��vЪ�I\1����8�W2�ފ��렶ŠO=�r�르j0��{q!ev��BB��LФ�
I����
�V�@K3�'N��.W�e�8d?=��A�F�cGRR���b�D4H�5y/���!���H����ڀEG:|Lt:����`[{�V�χ��jW��b^��:��5 0\�&&BH���ro%��V1I�#v�����9��2��;�8�����kN5AI v��)��Y��/�3K: [���i&��HV`G�� o�w@�����G�&T�:f��|46�-cm���〔����6�2��/�\�Q8������?�i5l��i�`�v����ڣ��w. �>&�w
1�1��,���%ʪVj9��%�1�y���E|��X�J�3���1�ҩ�z<F���n�5H������XE�~̔RȪ"+�.,�Q-VsLS>��l_�����K���=b'n[��C�)YGoL1���������mnbo��J���?�Oz%��BJj`"6��Į8t����L�6��]
v�5�]�9���/�U�'J��P ��xEI���= ��( ��xXn32		Q"9�	�?/c36�Q0�,��Ϭ���3f�d����L���֑ܶ�юbs���Z�$�M�K�y]�d���}�R}���yb��yJ|cx��ha�i��q|�]�\�Ƕ�Ӧ�3�q��|�b�1S�v�3`���7�1DWg��X��S�������{����L�$I��;�4���X�(�Uo�L���Tƈ0!!C���u��,�l�����)�!�#+�k��j5/��m<�6�l�������.6J�#�K��C�P+�߀��]v��~@6ƬN༅ƶ"m��՚5�=,a��7�O�\k�<iس&�aP�O�Q�5jV�e����f��j�.)�0���SQaq���+�v��1��L\}c���j �_ϔ����ӻ\%��t���ڱ�*
�p����!�~ia�TY�1�(j�+�����G�d����߇L�3�J�Ohh��6-,2��ŀ~I���v�OO�{2js���]��6�'+8��J�L��Ӭ������h�_Ӗ����Zv��l�+�`1Lz~�g���:�%�1��)���V�t�������z}����I������4Q�����V�8ˁ���Ut�/e1��_߽A�����?����D���;�j�������r�"w�(�����p�,:Ъ� ��2��-�׃�׿?�ރ�s��-���c|oId�v����eN��Cp�w�QHʶ'P��@����L��xO:�M����@��ܣ	��[t���*�:���Z �`$�6 �US��S�G�[��jĊ�l���E��^��*����^%�q�"G")����Tk��r)AOg�;s�D�1p��Eذ�S��x5�"�s�;�v���}p;��+!vu�)K�����φ�^Y�ݲ���D;N��-�j�/���
'���]	���*��U-V���Z[rW�O�$H}�6n���c�
U!5(,4�#�'?7���+/�d���=J�~^�1�t�1�myNt� �&lRV �����	ah�g�ӕy�'�>4����GQ�9��s�no,b64?2{rXf�Al/���<E��[�F�<��q�m�S��+g��XCG�<E\�� ��c/�e��|�z��b�CalPv�`�@���\�vX8�{zBj����V"�������1*��11�7��ڜf�$Sr73�i�Pԯe������B3H�I�c*�� 9��^�ڡ��4(kuט�J[V�=��8a}yDӑ�gB������U7GX����.@����5gei��Ɛ�5L��&I��wU�S<I z�Cŋ){c��hl�fJI�U����B���Ɉ#^s��kh(iN�n�BeU%���)\n��l��Rb�%]��%��ݘ�R�B�˩������6����~�p#���Բ��L3J0�A�$�l9����"I�)�k�e<������7�-��q�LO�w�)�=�|0
2S�KtZ|zOQ�VZ���x�d�v�����E�y,�+�c�t�(�����>|s�`r!�Rz-�
��R�cO�D<(�]؜/1���L(I�I���4�x@l���t�l��������z�Kj��w�2�\)a�"��Gd�>
`>m�V�TŎ�A5#�V����ٵ����:�ި��1��}Ć�|�{�~|�`P���G���¨=�ߐ��B�l�ف��Q�q�
��|��&�|�a+�2�h;k�Uu�=��ߴˆ�$�{�*�8�	F������)�Z�+p�����2�#h��r�a����G�0jEe*���A����"�U��&�uۛ�����C�1�+I�7����&���彤�^Y'Qg�#|����hY�$��p|�p��i�ƌ3tܩ�G��P���-bv��U��~�T�w�s����NlE�I�J�3�o�O�O�A�}�fi�(����等	�E��Sbtd���:� �pu�Lـ:�¨I��4�F#Dx>���o��'�m��k��k �����?Ėfy|��L���ȉF���F�:����؟ѣ(��6I�Y��*Im���K�L�ŀP9��n����bV:z�(^����8O�ω˲�4k��)�J���9�C�S�F�Z���$�_��f�f�NG ���z�ٔ��X�z��}=.�e5Y߳����2nlS;���ޅX̦��;Fv���>6/��۟����8uYԈ�i���d�{2��h5
��(��9���Scؖ<��-A�r��fe5���<�b����cC(1����=/�q
�ܿ��̿���˝���i7��	�.���*��]��7^�α��߸5�7���A���#�]����X��V���UUךm\(X��\����� ���J���i=�/�^��ÃE���|����bD/n����׈����c��Y{�D���ɳ�W<��3�z��0��9oSN���©(^��v��&��dI���潛$A��v'�H����1��<cm��t�СW�~�P�&͏�\�[n�O,^�y,�O���84�K�]3��NҶ��z�րj��o"r�ӓq'��df�Q�N|��^��P�b��IR�!�$�XdWkiH�B�����f=V����Ky��$�S,��H]�^ԧ���=�r�3ZY��g�Ff���������y���
o����6�+X�UHY�2�v;P�a�c7e�Z��&��n��-��o=1�dd6p|$��4J+I	]}�B(� "�k/ݺ
�[��P0)��w�H����`�GD|ᛟw�h<�����߸�Ytp�h���T��N𛽢�㹉�$н���>��u��ğ���˜q�\�������(��*���1���E���xɁE�=�LmS�Gn��A�n�2��n�f��A;ꚩ���/����<�:v�X�7��V�>����ۑb������s���3�<첐T����Nښ�����s��0��$�A�Myv�y�ŻX P:kV�xfUJ��o�d�x���)%��� :�Ɇ�Q���s���$u�b�K}�>:ue���%O	���C�%3$�Kl�TL��֔A$\e�"+�oo�����8��l��� �A Q}6�L~Q�F���YV�����Jm.���gp�d��4:��04Eԝ���C�|�����C�|\�h���v�.�81��+�D*�%��o٪�և������ɁӼ�(h��z��Y�3�Zf�{,�F=%��@p�������3K�4�T����ߏ,�)_��m�X%��O�YBT@��
�ן?9�?mon���Pl�tx����;���{b�.��_�č
�@�έ�(Z'�F��V���n���DC[���-�2�D�x,��'Δ�j�Ss���� �L#�
H3\O�����@�ѳS�L+!�}��_�8��[�;ߙ��"�������R��k�Hf�l�\���d]خ_Tn��n�N.�X�7Yo|�X��y��4;�

����� ��KP0�HAF�-kcH����t��7�k�9@O��%.q��2:�0^�*����C��O�iL���FEA3rG(������s�Z��ry�(�2!�>�jښ�W
M��+��o�����Q�>��Ht���$�h�_�$h�U�F�`���
0�"y�4�����J���=�a !C��0 ԑ�,!ܴYn�uq�844C1r$j��U�bT��Ҩ���v��Fy��C��vK�������w�����2]j{@V\�$���f���O��][�aI���B��H����Ü�*�J&	YZa����E�Pl	���(M�,�� �����T��a�p)N�_:� d-������rB�ͱ-��	��\Dߣ"#�K�����\
�4j��y
u������,t��@���2_S�m���0�<#/!�����C��E˒:?q��K�1��� �q�t��O:�żߵ��8!�? ��h�n�ԗ$w/��\��<cGo3٢Q0����x��}5>PJ��1�mӂSA�ox��d�q���HK�Մ��9©���y� �A�w;"��j��L	Q8.֦��4�1�s�����������m�׷��wꮪG�f��g0��\�,�Z$��\�~���c�«'���eμ<��k/‐�EbC�Ʃ��W��o��0���g����ф��e�s����i�R��+7ûu1Լ���z6�V����$ZF��y����
 F��󯇊O�Bl@y4K��IF
��(i�.;�R����A�X�p���1���_Am�9zBG����w%�A���ǒJ��/�o*M���'XK���c�����	+��L�?h�[#Kr�Y�P�r^�w�ܰ�P�YG��Z>x�m�1�9��f�3���&�?��Cʑh��ϔ�+��:�	�L�$��bt�H�ܻ4Ol	D�R���4�U#H�!���&�����Z�3��j_�P�NFa�1�=�I�׶7L�9=��\fN��Ex�NO؋��ۓo�� g4���{�H5pg8٥���Gmѽ�1	[�,�\x#��.��C��u�6C��g����&C�<�K�bԙ�N�`��SP�:�����I�fb�:���S�)���q;tl�T�Y�S<|�dp����Q���@21���;��M>r�N$�ҌN��?�Fg�ux�c�N���bs���ɔ�6��3} x��!���̸[�+:m�C�2;J�$Q�����Ke��f�7ѓhs�&m���؉�o���/����|��2�oy3�E�
@,�І��0��
����k	E�r�3;h@�"�;v�������m���^(�����R�r�#�^�8�c��YZ��:O��H���������(��3f��+�L��0Pz3)�d\ad�~�
ŷH!)������b镳2˯ǩ�x�I����$mf���D�G|W��3�z�����h����փ� Ʌ^�m�� �{��-��wj�y^����`�k��e��=��P�ȨЖL��ymT�4z�'mR�����	���I��q��
��>_!�!ă�� 4�=�Hӂ�c��47`�D�O��gʄ��V�S'�����\�o�dϮ�2�Q~q�'q]�8��߳Me�ƇJ,������s濦�rhW����C��@u�H�$B��������
a��")4��W8�{�h��F�]�p�̍F��$���)x��\��Ƴ�t�nT|"-�;�Z����qޯ�d�S&�pe7dP�[�:3����8���J����;�U�ca��J����G����Kބz�|O�QQ�5�g�[��7lٚ�k�<]+'�=�+Vŉ�x]H)�T&�]�J�H\��Ĥ��%mD�ᨉB� D�r62ID#zt@?�6�U #��9��>I�vV8�P
�w�'��M��Z�ANܹ9Ri���:|#7���ZO1�K`�4�e%g	u�W�����`߻`+���������99M�ܣu��H��1��m�G8ܷ��^'�
���j0���.�|a�C���ݩ���q;���3>`R)���1H��f���+��K@�N=.���0������w��$�ѪOKyi�cb��K��}�K�~���;�������=옽�Ŷ`�S��
{�S�Fq�3{�i^�M��$�hf���X�S5S�f�/�^*X�ؑ���02���`��������6���\;kx��;H�DE�4y�gnҒ/s���k��=Q/ϫ�A��j^�;n%R�+M+x�z�u��j�hK��>�[$�8#-?"����mӅ(�3u��� .t'���U�8�+
�`դ8�!��������@a�ȟsb1�������(Av�'8�(���N��0������$�<h���Zqo���;Z�6����MˢI�2�(J,;<D��\�̝���it򖧞o��`-����aW�U�v�$R��gf ���:: $� �i����4}�UĜ�I�͎��L��(�4χ���Z���`5ܪ����U#�Ճ&J�W��z�I�,���l� ��I}�������	5za�3�o`j-z�S�q�J��w`)����c�w�g�Ԡ��m�:BH�h	щC|��.���Ly$R$pSѓ�}�A����0h�_��qy\�������y�UȘ1��o?� Y�n�LZ�%��w)��ȗx3$�z�t�!�>�F��Z�"��'9�~t�_Y)S�
�e`����kh��Q�-�@��;
T�S=g���L��ʴ�y��*�O�a&KV�%~#Ǝ�]k�m�~�u(��0w-s��V1��7�����9S����<��ʃ���������$�6��uO��	
aq��g�Hb�k�Tgc���w:�^���V� e\�kXs�̗W�x?7���h��Q�����+&o<���H@,>º1�ٞraG��g����@��{�0��^�+�d���xbs��^zL�I]�͍�|��I����C��ڑ����R�����Zz����>n�t�8�Ǫ�4�(��M�94�����9�;�'5ɩ%l͂/;���nA 2���uRհ}d�r���̣]��f��=_fm��s&���t�r��=Cl,��Șի?�Ƙz��J�q���!����7���D)�ǜ%՝��~I��B�7�s,��$H�'!��jB�j��d�`i��x���~
�[h�����۔eI�����Wq�)�q�瑕Jqsma~!k �)n1?4��ĩ�aO�������y���A��9Ͳ��(�|H��̡:�K��g��/����v��c�XR6��m�k���]��я��x��m��uL!xe��ߤI���F���s�(��k� w������1#�&�����S��ca��I��6U����(���Ȃ���%w9 3��2!ޔ�HY��P�Q^*Y.�?����3���VyH�_�Y��W����n}��$���=�X�:���G�m���q�z��18hٿ�e9	�@���]Ph���o��mw��%�*����pLo��1���g�E�ékS0��!��y���r�c���GA��9W|��,�d&���2)�Y��L�e�g����}�3��	?��U�F�<<+�j&�6���3zeZPX`��*Ԡ�:��"����e�[,�Ph����n�1��Zm�����������p�2@M�KX�CQ���0�cY��6 ������	lp���P�׳�����[l�lCJSAV���d܋�a�ި����,�U+e�Qj9��ĪO?��@�����("���B�ɰ8��?|xW���
�pa��G�1�c%�m_��̱�R�߼I� ��놳�lUb�ϟ#sʌ�`��j爠u�îP���rpl��܏��\�xR҂^����1�f��c�;�`鼑���B�ʒ �jʷ���9�kY���ƍʚB�����'I_��/ w�H�2>�V�L�o�k-Ql�-E�
P=�1MҎ3a'�'j�ۄ��|���"�������3uh�,��ا��[����-jj����z�:A�H��2��G<	tʪuǕq鳚&KS���q�9�K�\YÇ������6��1��!����Cv���%�5Ӆp�O�����R1;j���D�� �Ҙ�.�����=U��N%��H�ӻ����v�s��3�T��� �Gp�V��'A��tOS���8���٣qӫ݋��8�I�Lo׈a���"F]����M���D��f:�0�4u_�W��$X<��]s'���No/tA6K��؛���*�Wͮ�ƽ^r7��� ��?E��;8Ҩ����V�3\kyP7)�Ǳ�U��'JY��g�}���5R6�1���X��g�0,�S�Ec
���i`���D�\ǜ��\aT��VZ�;y���_O�)���0�&{�y}W�-�n>�����Xt�(�ەfd��I;���kݸ?�+vxGaM*9�];�ބD*�»ڈ�p��G����tQ?F��ܪ�P� �Q
��ݜgV��\ڝ�+PS�O��US���!��g8�LN?1�a��J���|��!����Q�ְ}�Ð?���y.��v@63��3k�-)ǅ�èc��5��z�QA����'��8�*�cBք��i6��ss�4�`��_?�8�yu./t�*Sߴ�&��q~h�(]���ht����U�q[b��s԰W��3�G�=W�l�䢈gɌT��b����d�P?\[��i�P�y�P����&�o�t��m	�e}'_;�0�r�.�B��2���F���(�����zj��{�:F�0݃ݠ��Y]�۵JS��\���׵4�>�x��MȖ-�g5"5�3y]ܧi "�.��|)z�g�!e2w =�P�<���؊c����Nj�W�UP.z�L
���oq]-"7չ� U>B;��y��}O��u!��r�K��՘����ɻ���f8��6���_/��T�n�<�k�ms!����+�,�a�7el���QI�������|�ŷhC�P���>�?Ү���|�q�X�ΝZAH"�՗H5p��-��dԌ�
�7�I8{.�-��y�G��vX�S�54#���4�?�J"��X(<X���D�;4V�	���k;�.��0*�n�EE�W
G�2D��t;ߒ������\�B�Ic�)�;��V���Uh<�f�[�1�J�M�7��St�����&�9ߚz�/N����_:k�U�{)��a�:�Q�k�����xW��� �_��1�l�#'���,��=b�;q�bn�6���0�ua��Ğ��nӄ��c�N������Dc� �7um�
u.���YL?_+�x4ܞɪ�P��,������Eе<�-�,H�[G�
b�Xl8�J6\d�N����=5���Aÿ������N"��K��8n��D~U��V60��Ve���HXļ�Ϝ��X���r�e�`a9�M2�,�a���ɍ�.���qc�+�p.�Tv:�	�~]D���7�~o��bX����CQ�v������Tt^ 1z�kY�pX!���G�m��!��Z�-M�c'���z����ʏd�&�//!!r)	���U���_��j�-<z�Y� >�`�����DT�	W�,��ݞª�A����g�Pl����k����"�_�W{�,@4���ʚ�ͥ�E�{MM%���Qs���,i���m��n����D�?�����y���3��4R��5NY/��@�SY�(�P�,��&(�UW; ��`�H��1_9P���I#$sE�kB��@��c��^;�)��{��/�U���^�I��t���Oh1D�'u�t�_����-��p�R~y���߼��0Kh/���TDz����a1in�ʇ����E�������*L+�7BH�W_��s�~h� ��l��b'�x���>T���N�a�	��`*�#����Ìd��*4�=��qvϥJ�4-���S����lH_�o����LQ�|İ_��
�ڠط(c}\��B8^��