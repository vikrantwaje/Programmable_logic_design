��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&o�5O ��2M9.��G|usk��5��-q/YC���=����['9���V�C��̶��:z�!-��}��{ʰ%-v��u�'G���nWD0.���i�	��Ӝ����X<����)�K�K��Dn�t�~�4��̜괅�#.��]d��� f(8	�Ј��Ve�.�sR�v���8��Rs ǋ���$)��{�:���N�r�:E��p^ÿn.Ģ9�5�ړ�~T�W��xd��#E$���i�?�� �ڠ�@��yP����#��C}�z<�L������`���Թ��S��L|i+�U�΢�Ȥ�Q���U��at�p�d������;��rX���u�������.<B�QL�Wt�e20:��vlh'��%����1ʽ�A��$Q�_폿`���t}UN�C�v
�����cb�\(+�^�5�>u�]3��Dp<�4l�L�u`��Ǌ��`JR�t��
�2{���&�x�3o��t�s�C��-��������GD�%�̞^t|��N0����S�K&�#��%���2P��G�ep�y1�ǹR������O����Gy0t1���1E���fc���Դ��b�\�S�Wr+���4�i~`?{�td~u����߄˻���V����=��c�
��v�j^l��֬v(a��K�W����o%yJ�8ks,�3�1R;���ʓ܁��7H�G0�������M�:U(D�]m��c�]5��F4<�\vf�s�X��`��:��L�ʻ�� ���j��cYQ���|L|('��:����MA�j�dLéc.�/�Hh���5���LHկ��>�֡��'�Ӛ���޲��]��,2oo9�ٲD]x�B�v�t^��t��¯2�$pBb�ŏ����W�Q?��P]�:�	 R-^S[��W1@��/�������(^@�m�c`~y[�����f{b*���ֺ�tI3w#��̑C�Գvo�Q�?�!l0K���N�^(C[��~��WFyD����Ze�ܟ~����4�!fh�)/WBp��)EQ?ޠ�P#��#�7>�5�Wy�~G���f���Ps�?�&�8AE�������m(*rIY�AN��26�>FjU1��`&��N`{�%L���&m���ep�,u���d?���ˣO��SV�]�(�Dž�^�2��eΗ�8�V�ӵ��$�m&!Hj�:�����������ji)#�7/��p����9��z@7�<��(.�q^N)��y�D��s��
2�4����.�3��f��]�b:�'��b�v�T�m����-�]��E�e2ʉ�Vw|��뇸��../�2>��t}��G �5���Jʿ>0�ܖ�R�kW��|2B�`���F��3��5@��e�ZGB�i�b2x���ѵ/x=����"		*�8�Q@=�jS'�.�<{�?�f�J�'Q�}'q��
�\�����B�8��~���>�cɤ3�&)b����3�2�Q��IH�b��O�.!�$�h�7��%9��,u8�Bv8�0�u�kZ����"A�5Ƙ&�%�>QDxdfcK�}ೀI���)��]*�H�pƳ��4d0|-�� Ⰷm��O�,���mR%`�{xg6C�*pg�H��Q3��-��7��M��O��h�Y�4;V�-�t�Y�3��]�Pxn���P�gbm�B��K�H�L���#������N�޵��WY��E%΅�9�F�,7�E�'z`DgIzҟ�-��Y|��=�٪��#���x\S#����L0��ďu����Y��b�0��)�z�Ce�Q���22��h����iu;�0��gc�@aF�r7�A%"�"%yrQ�q�VQ�-Y��jQ(�z��KW앧���5��>q�+'��D�*��_�$X�+�a��:.{`T�uJ��|$����`ؗՎ�5;�������XN�S�}#%e���u�[�������9ٍ�\��nȸ�"չ ����5�N����3������)��3�-��v��� ��� v�FU�_~�AЋnת3}��꽶�%�`�&mq����7�;��I��hyY�Ih:|�\�[L��>��~����+�-�o:�pP�KT��m����Q�,c�[�%5�]�<��ƭB�e�b�@ʍ�A�r��k�J�~���̗L=�����,���P�ͻ����6Ր��&�v�'Y��������N�d�'�8�u�Sx��d�2�J���=XA�d����8#�����J��Ú�j(>仜N���o��2��ΣHnj��n6=�j�o�wh��{�ا�U�$_CFV���$��yX<��KA{�#�A�]$���R��r[>���1� �p�p;��tfї���a�����g{���]�T8j!�`&Z�{����/	�3���7>���ģ��l�>&�"�L�!E�%R�]=bo;�W��Qۗ	���,��,��%��	��H�L9����rZ�Ű�f��H�y�C����F��kX��f�Ѣwx����+D1�w��O�y5��� J���� :��Kׄ�N����f0änHL������}�禶K(���#��H�BV�X�8K���3���1�d�%�8��7�D;��n������Tk���%]�2�h�ۯ��:ǥ�3'��4HE�l��=�,�G�F�����v����� ��ׂ�8
S�C-�O*���C�H��9}���7��SR�+�7I)�5kƢ�iT�����5�gd�[* :^�F�H!M�G=�Y�k�I��+�2�
��s�`>�R�7+b޴�S���C��zm�H�������у�uO�д\x��7�ŷ��{��}�T��Z&�� _�̪v��{ls������e�ǄKoc����,A2H�G��v_7A�:����n��l��Q������8����>����IZ�]��zz�]�'3麢�l�;�?�(ږ��^��K��QLP������~׼(&=q~�gPE1�_�Z.b%��s�Z���Y/��z�)N7�VZ�bO��W�x Ws�ԎD�6�zYK�5��]�N�q�?ZY����Nmd����
V�}�5����BZ�u��3�sn׈&���]ʲ�E|~�
���Ӱ�K���D�@���R��Hr���AL���/p:���3�g:�yy#4���&������xF
pA�9��.�[D�T�|�tb[ك���a�7h�+�gE���� �Z��qcU�� �9�Vg�~��O���˛z��[dq�W������{��ЫƩi���#��A�\�^j@_y����͛u�+�%ÅR�-����k�W�>�`6��S@s�n��s�g��sH)�)K#�2��A��8�5�%�S��p` ���w���:6��n���?i4�Pc��֢�A����[��6-1��^��F�'������>�B��YUO!�䘻{ᇧ�.��i(.���M��^�Je�be�,�&�����������mC	��my��mkU5+*�}�����d�M�6��4]�]B<�U����\�+�]/��4�0���IPN�x�c�^QH�>�k�N��He��x#fF��3�#�������/<e	t��J����4"��O�'�`��o~��нהH�F�@q���$G��fhNkۑ��y�}Z8lx	g�a ���bYAh��Ϗ�-FBG
���t*�H�s�;$�H��y�6L��H*ˊ�BH.O�sV��C8A0�ٲY̦��NH�|{�H�Z���Ns��0bLV��y��ʯq���a=��M�4�p���-�}�����'F�����KG8���[�q�9�8�g^x�HG 6�����Z �j�2I�N��ʞ1y���U~��:z�Hsfc�I��H�9�*�y�ω�i�(0|����g�m}z��^��.su��{��[�)��x���G.�5Q֦Z�7Opk�����f�`P 10��d�6?Y��Yt��vjY,�9~;�T�D��Vqs,�#�}/M��!��:�t� �&F�cى-M)NP��d�������4G[��PB<ys>/aE����˧*���]-IQep���P;�o���m�����-&ŦeT��G�J���m�l����
�ݾl�+��|����	��_ C���1+�}��͛��F��_ �/ z#<���s�@)��E L�T[O��5Q#K	~�H�lz.1�[=TۑJ>���S�8v<�'�&�Ӳ}� �	K�0�_1��GΠ�y�����Aǉ�_g��r�ѦρK=�um=1ޖ��w�hy�k-^0��}�6��	�~ �6��Du��t�Vs�"C�Ŀ�����8�;_T��@���};Q��*�����Fڥ�����E؃�1{*�B1/�6��R^Yg�qe�ݸ�K2�]!��-��R��a�!���V���P�F
Pg\=��V�X�/� �^8�A�l��;��;Š�ڢ@s��i�D�M�8��36�>�����x�΍�D���;�WÞ�N�k.�)<|z�g:q�{�2��̎���L|E���`�}۠~5��U6�q-��s�Ko���R�E?Q�C���G�d��N~2UOo~.�b6M����(��za�_#�#�;�k�s���m��Li�����<��'
���Sg.�e������e�Yc�c��ʄ]�ՐɽZvݖp<�����7|W.܍+�`�uA��ĩ(ܼ
�/de�A����;�w������7�;
��|{n�;����l�;*�BT���r�\l?AK�ĸ�a
��O ���#W,�m\{�&�+���b��;�-=u7�k�f%� :��0fB���Jn��s��K�N&��m_�!,Jr|���Xf��/.�e�z�7l�����J��l�g�(䱆qG�-��,��YgkI13Mb%1&�M@���w��F9v�6���br�O��JX���]#t;�}� �eS�Ec�KT-���5�d����"�#���`��K������R�x�ʻ5:�=H��E2"����_���8�oF�|:k3��" (�����%bK^^��y�iP�����<�|j�辀d��ZOƐ�ǭ]p[�rh{�{�<>@��¢[����I��u�Y���B�����%����J�w!�� K��%�����rD��X�-�%G7��'A��ӛ���M(�t�Z�H���������<)�I冩Z���0?�� �/Ň⦺�������;���;���;)u��s�[N/5#�z䈆-i�Ul���1����B'k{l~�,��I9��7�}|�����{�l���y�-�x o��ay`h5������\%��e"l�p���bC���n�#�t���L�d=�D!���Q~X��z�^$�i~j*� &,(���� �,t+��T5q.�u��������g�_ ��a~ZT����i|����mbD��z��f�d�H��j�<�S�PX��c}$�(� �l��<2��]��p��w;NŅ��<��k1��
3��,�?L��������}�U���3���ka5V�&�,�Գ��P����@P�ݗ��+�¢�i'$��]O+����!��vS��o'LӿM�6x�V�4c��Y�ߩ�Zt�o����(��mgl3�h�鸸��HW���s
�WS�EcE�U�.Q^�:�<L��P�|�r��P�4���3<i�d��⤯N�G 0��$e,*(ޢ|�����w�_�u���]Tl����P��H�]ٛpfR��g/l��
�_�����yx�Մ�C�S�>gL�y`�ֺ�3�nI,Ѥ�[��0��l`=D�K�FߠU�17�(�D1�)f7�e�yLL�ȿ&̎�Ax�i0�����-��:C8>�@/�9P�WWm�+�Qp�XA�I!7Be=>oJ�)��M��!/k�L���'��q��]��9�Ҧ>��Kr�m�/�hj��L��s��m��Yc�����
D���
 S�uUw#zy� ���!�\����3��k�Tv��wc��ՄfW� Pĵ>����Y��w��[��(U�> ����z�ߔ�jq������NFQפN�E6���R��R���V]�)��y�i���ɱ�����=�s{\�mE��keX�b�}���4лB+
`�2����;�CK��1��T��_����]2Q�� ��_l+��0�C�@�z�9@�t�G_ȥ;|"=V��q�)L ��,���!�SXMw"���� �%�th��l���
����m\a
��Se^��#Mi�Ĉ�8�ü���%\ۚ�Z='���!����Ov�US'U�l�a�x
%2ؾAhxP�잘1`�e�\�� ]rń ^Ip��T��PdBp� !���e�c^�2;thL���&gX&��>1����:��l �P��`��M��>YTOm'F����-��Z��&�k%�ݼ��9fP/�p�A|5/���nױ�~=v��k�;�#�oi�S1�]�\�`*�h�JxK��7m�|����4�uը}9&���U�	��@��ܛ�U��8�qY���v��vUpɛ�E^(Qʠ�u�y���s��R;㎽��/��)\�倩�<-PHj��&D@��_(@@�Ґ#�-�cN���� !�<��wi��mR��7��.�h����&��	zH��;���b���k,��?>�M�u��L�?V��`z� ���!�d#�"�i��[jT�*ګ��t�\svr%��m=����ƾ��F��o�)i42�yN�I�c
l�4�x>d����*$w�������R4?k	�۸X �,��Pt�3��3�`��������+��%�;DEf�7ض;# �q?�{8�'l���͜�~J�ER�K��%�6��Bh�-qn�M���0�")U4 �'�1�R'�7�(?���y]M@��,e�����HpJ��ٿ�2�\C�ICCO g��Dx�]�
�����j2����4��o�d�]�/�O�fnl�5p�9��#:�l��r�.R�[�E����3�k�ſr�?��
89ݔ�����{��"�;-y�˿o����Z��wI%cJ���c�Pww�7�5�l+`k��S�v�pLϕ�q�UǗ�2�ٸ�L	��e���Á���i���v�"Pr�\3wف��f�m��%�㮗ည�2Y�1�� �i~y0ؾ�ʅ�͖�Ft�JU�-�BrMht�����0��|)��>	��qT��E�b2��,���+��j $���{P���zvr{���6����R"�d�k�/���Z1#L��8��k���RߩV��(�BAr��T��N蝦����`ۮ�<�OHQ*c�7�fo�M򖫸�L���A��NUg`��!P�ce�9/,67�i�H�����JW��#zAj�NC�^W������5{د�8H]1��-�X}H��5�5�k����n�����V�6��i%f,Y��p�Ã4WY�=�=@�l����m�f��V�6�%��#o�m�����C����ʱ�g��-ȶ���^Ͻ��y�9CI��#V�@�������饈��\�n�:B�&	/�l��A���/�ݽ���7w��X��I�g&��� ����t����X�Qf�����)���H�6��yiOL4�,'?�.�o��hp�ÿ�֑�M��ȟ���1S�B$��}�ϙj�^&���C&"�iw�r"�ru���[qY��š&����9 ��V� �B�BB8YT�n�u�驪˽zO��矾s0��@X֐}�Z�bUuh�6F\Cg�$^r>]�4��?S�]�7��q?y�I�3q��&B���wY&e?0i�n~vUGxѐ���E�>3ֻ�$s�B �aI������E����
)CH���'!Ѥ3�mj�EYsD�9��"g�ۗ���*,�	�O5���p^v����G��Ru?�C���s'�SxO���/���Lmf	���p���y�m�G:Z�hT�W(g*���(P�xK}�V���A�G��*Ԝ]+�/q�rS�4/0�)�]��I�*J�7[B�m��_��þC��g�n#+`��}��M;��j3vGܟ�kP��rh:t���M<p�ζ��L-ٮ�Zԗ((LsG�!Nj���ۊ1nl}�T����8�ª�U�x�ξ��D��;�&V�-��2��a�U��!ւ]qc���_>|%��$ZΊ�VZ��5G�9oD���e��^\|g���s� ��k��Ҽ3�$�\\�{��L�ZZJ�0�"!�R'or�L����;#��b�������7q
�U^p��/s�AY��_4jGz3�RS�z��x��k+47ߡ�i��ˠs��$'��сB��F^+ �g0󴈱�8E�
 ��j��Be@� KÔƕo��)R�(��M�Z�j����IZ[fH��zaT%$Bg)Kt���\(́Q�ڸA�>�	@����4<R��ԅ.ֻ���HVGR�1FKX�?!��l��n�����Ƃ-�>���j;����3
�g������D�߱5rJN	D|��kP��tW�Y�m,K1�&L��xy�'��H4o�6���u��̻.-�������KDne!Z�[�{�AXG���~OCC#$0�SV�p�ː��7	&KwYY>0�����k��*��-�� ����FZ��jP9`ʮ���n: D@/���ٙ]��~U�����|���A�2�Ҝ�`�w�^���Ƥ�3��εImy�"�{�KO@���D���8�a���v����&�vQ���r�?І���&]>���r��\I����x�D���<���"������!2��o��o�Dۢ�#�kgJ���r괒Hy�!�&�=[�E�Z�DE6�A�(lZ8?�y�	p�o�H 0Zs@�+�Q��X���/h��R����V]q���TAUB�fԎ�R�6��I�FP��^H����|���:���	/9�PQ��~[�}��s�"��E@l.:�����)r%\@���Dl���'�hB'�!{��</A��^2���@eB�>&-����x?��bO7�Y�
�ƿ�þ�Y���ү��#:���Ą7r��P��v��N�kN$w�R��/���W���A�/���ĉ���Ҹ����O�İ�X�^��>�����6��>�^� B�ۤ��a�@�'�e� �&��.BaYp܍��&V=և3��Iu9�m���X�����+6��l�
dV��x1UϹ�[#U���`Pd��:��D���AT���@_�x$l����>� �M�$y�
��Qp�N��i�a���S-��o�����m� �R��Z�I\�6|(#��&٤D"Ȼ[�±f\�>}����y@�������ª�[P�΋�0TE�ӡEt���A!�h7���t�����j�|zS����~͂0=T R3���
�.�|Ư�_���ސ�3�P$a�1����ͿV�Tgt��3י��J�B��@�E3b�f���W44V/!��;�$�^ p1���W�W%Bا�:5hY�:D\�\���@^�Y��@�cL�`�8̗��r����� �6�L�N5�a�~`���M@qz���Os��38so�}��u��{~�=s�f�(��Vb	+M��������:��E��{w`3�T��h�ug����.������9���T�Ĭ��
#�]/���4!�$SQ�t�Fgg����L�����(�ʸ#x�t��\�v���D>�M.>���p����@��Z�G8[RX��O1�i�ք?�d�,a[?� KH�?]T7���������"�:��v�s���"�����j��:�j�i>����Z=��-�H�p�)(��RY�g����<S;��J9��ja�GP9K�<7L{��=����C���{���z�1���2w�X�$wY.]�̉T #�'`��H=�M�*F�ץ�S���_�s��wp(����vw��:e����������n�k*�!�rҺ�v�D�T0|+_�8���^�m�q?ـo���q[Q�4�שǗKRp�|�,�(h^(E��`qަ@�[5��S���Sd�1*��m�v��O*0#� J90�h] "K;�����D��B#C��
�i�����y�������Z#H��:���{KpvjH��˹|�}F� �J��������#�UM��졧�N;��!��~`r�W�.0���_�Q��w�r>�O�:�� ����x-IB�]>�&	ڔ%(A�Jȃ��1W$ט��33$�ح/X����.��+X)��{'�ߛ�5�+Le�|�v���ψ� ��1	�����?Va�2Ŏ�h��Vz·y}6a�d���9�YH�{O+ �8�5e�����;��ΞL�y�C
�NWpH'a��a8����B���fq;�=��N/T�,��%�5�/\_3#����f�y%�w��u���!���9��s/�t98s��c֝�/�+���g8>1�L|�A�D��!%dI����K��੒�PK�U���_>�MG��w��/���Kv8#�yzJ��C`Ry�lAK��#>����_�w��}c�p]��ʝ<�N8�0�^�$-�����Ly�%M�'�b�Cx�������b ���G3�K�G�s����p~���̩I$H
�m~��[GV/D�]O.�d�;
��R��N�~�%�����{E�S���*܀x#��H�n���c^��1<�
�o���R�+�:c@=�v��ۖ?'h'�
w��Q��+z�\�x�S<<rw�E@�0s+5�cd�sa�5�E[��mx3������`?�-���)_t�tpr3�E�Ggr�v ��g[U�x6Ʊ>�݃��Ы�*��ʁ�婕W�@�sؚ�����R�W��b�G���
DW�o��1�)ֽ�v�5�\>�x���?铅�V�-˲��\gf th�#��*~�j�%���H ��	��x�z���r����b_$�VW�W�/���g�i'V���h-��c�/�N�{_@گ�f&#�9)j]Kʛ��� CP&��v�{7����`��°�ۻt�T�8d�ZI��-�zJ��`��x�|����ʢ�h�|�<2�$�O�ơfY�R5u������*�xW7�ci}��{ȫ�9�܊���0Q]{�cE����<[�i��i����dm�W��@۫�\��KA��� �O����]t#2>����[W��������w�J���-/�kߘ}pH7� �(����3����{��Fc�q�68�e�8�A&��x\�V3��� 3W<�7�JD�"�"$�D�L*��3Y�B@�y�j��bXvS(Խ��4t	Pp���T0h��e����ޣTI��k$j��X�>~ �8�R륆Ǐ�]���y}���^k72�jTT8��w��C2�B����z����8)K$�v� �##��#vflGP����!����G,p����Mb���ϻVV�������t�g<:^u��t���Pt��1��|�Ҧ�����Y��s8�0Oc�w'A�V��O&^6b���.�Ԉ�LlM�Ws���<S��k&-3{;��=3�>�"h��(TCr���A��晹���4h"�>�n0���p�E�zP�r�һ�\�ٟi-d�i�2 ��ZF���������&��'�M
9s��㟒�.�-�p)t�&{�Ϣ����𓇑�Tɂ��s���곁���?ʨA�U�����PI����6p�֏�����A���HJ���wA�1��aт�L8�9��bx]~O���:a,��X�e����4	�3����{8k�������6�:�,�a�h��h���xi7��Ϝ~P��y�2��T�N��� �]#}���(܃��k(�B�1�mB���p,.�BTC'�_�{6k��vV��y��f�����)_:~�?��,;e~x�K�qX���MQ!Rp�(g�M}x�ϣxכݙ�V\=#��ň �-5� KV��c3O���VV0�:;"����J��v�ff����,��w�{�`Az���1�b��HF2�Z�*���jɵ���-Ոi�Y�_�K��Ai>ȁ�~����M�?�y�x����4��c.v��cQ��W�}��ld��ѳ���8Y���ߑ	:�S����d)��&�o̢ԣ0�=k���L�K�j�&vΩL���t����m3���Ts�����`6 F,_ە7�I�X��qƟ�ia_	�c�/�
���H� ���FBQ}(�0+eV�h�\��`p�����$%��$E2�[�f���g|\��;[r��H2�֔i��,Ɗ�-�1��f����m�"���9���>�����\$j	�	�2�� ��\�Yvm.��m��j
�W�����&����~��P��9L�h��L`��P1���C,} B=r^�t83B��gZ�>��h�:2,4�}s|��[�;������30\�6��CDcW�z�AfCCF+��9/U���F\����PC(��Ubh,���F��ț��FP(l��U-p*�|�z[/ �P������7E$|1�v��˿Eٕ&s�d�%'���+��y�����~�R�衐�̍����ID���� �@�!���wZU��
|�9���Y��V3�/�kD ���qk�m��Ů�1�	��NI쨳.�x�J� ts):!��@V�m+:�7�/$���n��zp�|)X��X���8F�����Y��*�0q���i�>�nt
e�}���<B�$�D4�\��<���~��<�jo��$gI�܄�J�f\�������TC�)�	z�R�^ޤU�ᑂ����Mz�.��ە�
�lo�v�~u�eb�_�GgE���g��(T���*�&Y�/
�v�B���㔲���1�r/J�&[�#�ToWu�.���Qa�i!���`H
�v���ZJ��	��^ċf�-�x�4hk@�!�*�p��o|_`M�$��T�io�T��Y�~a�RZh��_��]��7@z4�0��D��#�����+���-<�Y��
3��B.����(�&��e�_��	c�	T4}H'"6Y`P<��fH���)~SA{+r���VE�+�y�(�WDSJy߅�N�'��U�oG�:�x��'~��e��3�jz.M�5��'�u{ ��AۓRk�	GL�=*�W�� �S��)��?֖�l�2�+���ϭ>2jk`�
�	�Gh�B��`��v�+��R��CeO�nk �j||WLK���gs�48��_Q��>�t*�GL5���^��|Ʉq�}C���O���6g�j�@.��RTX�Ґ��^��4��u��3���0�g��*L�_ˉ����c�Ln��	��!wE�o[��z6�o::�&p��-��b��������U�%C��c���&�P�2s%.��
�{���cg4D}u'�dŝr#~ю��K.e eY����{��|����z��{�^O"\9%��w����vi{`�UWjgC�����pr�9�y��6ڷ�k*��0q%���*ʅ���x6Q[b�v�iDp8�8oc=���i{r��¤��*�.������禤Q"��Y�*yx�?4���< ���P�N���߽~J쐎|"4=�2���0/��r.��a�ꄁa�.�H�N�F����$���@�PԵ��{�E�?�Q�_H5��e���������I� 1��D�PS�\ll��e�G@��n�1?ёg��x�)������ו�ò9n�ΐ����Ăi�d̰�))CGa�[�)��4�5���.�`
��ǜK���x��KӟTC�l��P��E7�3��>��Џ��������B�'$о�i�}�
&-r��-ցra1�tw[�S�>8��r���0�y�}9k�h>(GJ�m  �S&<�$֮E�
��@f8\�Sq��.f�Ӑ)�*�'�&�!ND㙨���*<��]�?�9���PA��eU�*DBs^<���{ɤ����(ܵI%ʦzp=�g�חTb��߃�A�t���n��m���bzA�/FU����M5����1�]�����}+<X��>I�є�Q���=�Tk�����~�ѯp~!�g8�Qz�Qh����	�_x���+0q�u��4mf�,�6��H�j*	���«���V�4o��b{H�����K�s�Q���듚,���QWN@*M��-��:s�i��S^��@i��y�U���0�à��6��F�R"��u�=b�;H�U.�Q���m_ؚ�Z5#�>W��qw�|ɠ-x�7�_�shq���-�AS��㦻�ð܈p� ���@�f-d(���Oo��aZ���#����<��&�hw��� z�b�i�p�My.���_��Z-:{��R�1V���6I����fKio9�U2 �bf��S#Y�<Uv]q`G� eJ�*�;�'wԮ�Y��S�|�"d!ۨy�~+���ḽ ,��g���8�G������:��/��œ�Љ�+��QE����B �W֙Y�Y��`���TM�
|�mt���q�K�h������e��B}���~s�ø���^9���B(����6�|����6�t#ŧ,��OF�?��� �y�nX�6�!���М��w���+�D� ��J�ԼL~7��R��p�v��bA���*t^ަ\��o�a�Ǿ��6Ao�����nO�Z��#?I�5�0��}!3�|b\6#�F���~��B\@�{B�$vAmֽ�0ܬ%�E4L�&=��g,�	ѿG�8��P-t������n*JV.A�9Y�h2�5���#'�����| ����,d��v(��.����h�%��G�G������Oخ	�l�J=�u�\ǮlE�J�>�wg���#�uC��Z�C��me����+/q��_Q��&��g�-}��֑�4a��{7�Q%=dk����O�Ms��ӝ���^SZd�6�
5��H�31\�O�v�����Ϯb��dDY;�L�� %��Jq�k@���IW`{Ӥ�^D����<�۶����j��9�A<�ì��B�׹׈KGOCc-�X�� |�r1��,q�����P��E�e����~����G���#��@Ǳы��w� 6�1>����^�W�hؒ�T�w0���S-VZ'���dS��(&��j-��)$�گ֣&n=䈦W�	������6�B���5 ;�
��+�湗=dMLļ��}��1�+z�`89���-�*O˦�2#�X=W��GIs.�ԗ*��'�|���r"�4�P1�V^����Dܒ(�I�T��a�I��:����]��ݙ��s��x���U��ԁ��'XdAt.�^�X K��C���0��Ri�Xl06K������v�r*�#O��^��3�C�W��N�I������ѯ���Fah�����Ǽ� +�7D��87訢[Q�0C���!�&7��$�n������a6<e7�n�@�<����W��wŲ*Q%��裩�Q�����G%�$+��Yz'9"�ę?���͘-����+\4ֲ'�"�K�&$b�3ˤ��W��m0���:r��mnǰ�(M�f��Ϭ��J�l�c��&�x`�
�|jm�]�jOc.��d�3�l���h�:u짷��