��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?C���zb��+Y�GXP&fO�8a۞�sI�k#�٬߲ "sA������w9'�(��q��4;�8�K��G�	���s��j�/+.A)���o��BJ���t����D%$�$6^C��G�fO�.\���md�vVF3�~��e��\�k G���iϐ΁�O�W�ȝ�v��a-BCO
\w#�0���SQ�Ƈ&���)��KRؘ[g�����>��>'��\���\.&�����H[Z��&��3qʭ,�]��l��nB�D���ֿ�=e*)�p��'\�J"��\GR�(��}��W{4�[�홋S�9�4�7�l����;���L9��Ul���Bً�L�[��-]�Kq�n�:h��^]�_N�9��犢�b��������Gп�$m��8N�jӻ=���X�(�ˬ7>�Q#��rX�hj�+S�6� ��!8��I]u8���F�It���M`s�(q�D ����Kԝ�T@��e�)M��LPޗ�U�qR��sL��^�����������J���6�$u5��-?��0vJГ�e�
��c0-�h�����A��{�Z�/x�-�VF;6�m�X:��z#~�&#�h\O3�@�6���BԵ@%���N�d�V�2
�l�5����M0�Z�#��K��ɟ�l$$Sޓ��y0*�n�Aܹ�%��b���=����!l�\6��I/���<sm�L��q�w�]M��a���(���6e�{��
u�96U�����	%�Ñ��E�nX(]�}�_�*�(eԎl�/KB��,�=0�Q�EB^I�4ZXy2��j5��=qmCBE��YA{e�ՠS��>��x�X���sI��Vcc$�H}5��г�KD-�t�{g/:�Ry{��Y�N�tWD֊D�pTC��<zU�M]�7S�*~����w�1dE��/���&�a�C��+�3�M�O���D�I7�w�a�gBG��?L��˴ҳ�"��K���+�:f�x�,����4r����יh��0� ��S���y�H3��k� ��-G!�/]���1�G�8�x��$E�_3|�-�s_ע�������_���l��G��̜18M��eᖸ?c�����?1���<���� ��Xϛo����=�ڙ�ujD�ܔ�����uAG��g#�ܲ8p�{��!��VG�\Ĉ�p�PI�W�g՚Lp�>����$Ɉ�"f�L����K�@ۿ��֘�����Q�d��@	;����۝��i��
z1ل}���&��?z��,,U2a�X��5M��9K���B�,;D�'	#��go0����8q�*U߽��Z*�{	�3�Y�T���8�ո�)#�L��.�X�*>ާ��u-_ܴ7Y��j��3�(���ŕ)�l��Z�<*D�'ϘS�f��o��x����6�B��.���	��CS����V�a*i�c|��P�@R4���R� �����J5�����uf�D�Zp�v}	b;n��)P~�W��ǛZ^��һ���=��0�W�d3���V����#�'VfE�S�d��VX�'�,!�I.��2���y�P�d���z|����/��n'��C]��K�]�N��W{���;�<����hoQ݃�X��f�:X�OK����;ȝ]�V#�*�A�1���8��7;�+�����n��YƂ�3)�/��eE�:S�O�P����Ћ�`W��?�v�gY��m����� �lr��CdR��ǲ�����i C��q{z��8��¾5����SW}��)[���b\��"'�ݕ�Q�s�K�z�9#�b���a��US$C���1��(�.�Yy��I!�jiE�;�*����}	��%,����N��g�u�4�L������:5�<�^��%���c9a~7:���yg]����<!?<��^/@���/g�+���VA'�'�����|ƒ��sq?����V�j�ݕ����]�k�"M��(�x�]��1����6�O�	Ք^F�,L*�sO�Li2�1���\'�J�D�����g�����u�g}^آ��
���t2p���)�kwi�!Pę����xeh����?��j�Bh�h�G}P_�6t��/�nK�a�)�機�����#U 
��P�N��0a�eł|_~�>�?Q��)�u_'Q�\4BB'�	�4B��uQ�Ͱ��TY��i��1��,H~e�a;���?����� �]����\�$� �q<L���!a�c�Հt��K^��L�z���������Ƨ��$/T��d���k3�NL	g�i�W��vgy�Z��l�Ӵ���}�V*I�}��[.k�xqKv7R��[G<U���,[���"�����2���o{B1�oh��N��x�r���f����`d�12�#�ǐ+S��D�����/|�A��~��֒��:A,��@��vv��n�j��7�`���"�%cU�dɧ
�;���/�i�)��b}8�3�z��Gػ��<B��XPqH$���1��U@o���ɤ��6*��p,c�6��b�7m��0��H�:���S��^��C�ډƨ��k���خ�ÓE��&�b�ӧ�旯
vVD���n/��j��ո�dsaIj	�y�f��Kξ�Q�Q�[[�V�@�^b�JK��$�y&-�M���3Mie�%����{2y��3�_=�������r��O^�n9G}�˾r��-�	;� ޷�+U-�ygs�T�i�z"w��.���8��޼�2�� *��0x���W��^Uh� �t�\�iv'�¥�L�;R(	�'���=�E8=��Nx��%R�ns�h ��!�!�0G���ܦo�g7A��u�T�(��vM���<�x�gl2r/�zv�	�|�hu�y�g�/� 5�Wo[@p�oӆ��oU��Y�o'U�up���u�=���Fu��H5cC��c��Z��cn��!��nj�v���N�-��6�fxg�&�QUAu@Q?�L���{�Ld$3���3iT��Ӿ��E�����\��%�{ȿDuX>�h��Z����,gB��H�<�;���L���;@�]�¿wO���)�4)aն�m�L�4��g�M�i9O�o���X���_?*l�ܐ6%����ϞcʦL�$!(aE���W2'���h8~��N�Ks|ؠ}g��v����u\׆B�9$͵�`NBx3x,|�襤�!ע�u@V�w�h3�c%�uC��q�uꌚa�'�|"(�!��Խ�L�=:Z��L�[���:uӀfq8?���T��)�g_LF׺�	#���r�㵄�u�[����X6F���*֙Z��<�Ak�\��i�����aUr`��P�H�&��*\z���<��J�8(��zۏ�-+[�k[j�!�"��g�;:�qu�+0�����Zǻ=t०�F�C�m�%蜿��Ȗ,6ޥ�G���<lU��g01�����2�ϔm5��$��V��K��#�L�؋��hb����-�d���
H�C��H�(�V�vN�\ִ�CQ��\��br2!a�IY*�+�N�\�F{�U$t�c���Yǽ��ro8�f? �b��� #�u��	��q�"�3��O>L1�Iܴ�qi��)�.� ��"��"ʽᶒ
�y��4 ���c�軧�yu�x�f¶O��',{%�v�[_SW�C�q�-y�6i�VP���.[Y�� �(����$~`�N�	�7]HI_&��e��ⷱ�)5�xf '�p"�mdrj��ϕ��(�I��/��+�D	�RTct{�,�\�F_��
���(��fQF!�æ�sy��]�ft͒�FV !��Y���yѕ�!p�q-!SRi�lk2�Y�vS��Uf�Re��w/]y�2��S�T�y�?ViҾOt��}�ä(6�M�)��(#l��;�����9��0�2� �9ә�W0wirby �MR02��~��+�������n��^<$o��"��D+�'���j?%v3@�wH�����f�1qh(��l�*�W�5��/Mt�-|�_t�ES��͒#����Ka��D�L�kwq��Wl�m�wʻ@�`�7!8+@kH��1B���ww�lںAn�P�쳮b$޵���rH�V	���HFx��-��$%\�(ҿ�j5X���t�B�؄=8�r�=��Y��bI���k�e(�����qϻ�JtCr:rL��n*�b�}Skw�o$բ+���ô�O�[�%́�Qu��P(	�{8)e�=��u�����j�3L���+�y"�5-_��HT�EoaQp�[�a�������g5+�\�Lڣ$��yP����(�i��ʯ�'QY���7�hl����=Ut@ȷy���:�����b�/L&��X&��Bj(�3�^�_�@���؋����5hQ�o�/*u��Zf�x��TW,aץ3���|�N�5Ԉ���E�����4�6�w�!�*���H�Ѳ������	�]�]c�3T�FJ�q�l�3`=� ����� 
B�0�4�{��k\7^��O3�/"�o���Ėè�0
T+�������T�ߺ�l��u/e���b���>�ψv��ٿAs��$u×�	'�`���q��&j�]h�5�Ә���ޠ�a��	�	-��N�+vʅ����p)�f�'�
�VE.�\���p���a�E
7�닶7�X�'tp��p��y�x��[�}<��4�������������C݇�o<���:)R��h��ua�Gpt���J�ԮX�WP嵤ۤ�J�n��i�upa��ϐ��X�z�s$�`��姠^�������%g3�P�]q���6�8&���Zy=�J�z�%R+"9�.瓤�xٟ�`�7���*DQ��6�Lɱ�F������D6s��~��H�$Xm����W��ke/��t�)4��8B��$1��]����Y��>���ba*�+��I1@�P42����8(���d<7�ͽT9��مd�>Z�^�$>��Pg��w
܆��տ�.>��o�]���S^>'H��{
�������Ưq%tM��5���r&���1�r�N�4��.	L9R6�"s���#ze�I�á�S����gD��w�U�:D��1nhxR�&��ˣ��hs�e�-^��鋟�-^U�66��z_[�L	r�i�nˆ�nvvH�b��x#'4��VS�Iׇ��r��-�D+���;��5���W$.HƵ�^�Ì�yDs;N��B�Me�s8�������o��o���f���.��E��f(ѮҖ�8�0�����j���"��UBI�o���/{�G^�YJ�֡�;n������7^ɻKu�t5t5\8�D���߇E,�2���y�iԨ��q�4M沧
����gĴ5$N��n:�Ы��}4���I�A��;��;k�v��V�Y��^(`�o=I^�S)ڤ��`RY��s�u;��ǚL��~�r�U�G�xSIF*0֧����Ъ��3t��oKG9rae���c�5�j@M�np4�"��Qכu�ܨN*3�LU���Q�-ī�·a�T��g��p
�#������#�ߡE*Ej�n�4Eg�Z������ ��bT�w\�6D[nmԕ_y�bV�s�k��`e�#A�����}�cq��F,'ad�N�5�v�m&H�-�����?
�3x�w~Dو������'�}��\�m��}yL�C:�����S��f���Ӱ=�4L��0v���HrL��x�����1�T̓qD��cf쪖ׯ�Ğ4�E�2�|���$�:���Y.�r�iz�`����g����ڎ�[FhJ4~Z#����9^C�z]�P��! O�W�6��t94���H�?nڽ�Xx���#7X9�`�o�h�k�#���`NU���v
�V���ז��,�|;�$h�(�`Y�6
3��-�4g�	��{U�$oO�;�c�F6�����M�5���6wb~��Ϡ�1M�Z�f�0>.H����3��g	�߉i�I`Y>Y��=Q��9�o�I������7��)q�4��"�W�<H��u|��T�}�ͿڸP��_F&�v���P�����p���.Y�Q��:~zZ&6���t������[���F���eK�V�7J�]��T��m��Xc��i�C�]�߲7aK��p�nX�T��+�%&�&������t۟���LĆ82\�a��*4�8�i�����:jK���,=�����
������6��&3X���r��>�\�h��d����[Tn-?�G��/����s��l�T�������sã�\#��#���gq:�ԩ�X�{4���Fz�°M������GMuLg�\�l"����pS�u����u���z�������*�K����8-_C�L��t��)� �V���ҝJ�'�Kj��� � ��A���"�5�L�c�c:Bn�Z�T��5�ʭ�w��x�)��Ɉ��?ِ�h�b��\Y���d͍B����D��)����-�G��O��3����'��
�JSM����$�?�rC�����xK���8��ó���s���w�c�p�*)�#�%TD�_Y��UV�������O(��1 �+�I=�M`+#>D���p�s��h-�6=E�n��r��mGr+W��- T��*�N�)����T����t����^�t�HYD��QFRX��ڏ	���s�g7��EG	�D]�KW1^��}��L��w��*zO2���mC-g�坟��U%�ZB,jߘ�A׊s&� &�5R��~�z��)K]B�f���9��H��g:�[;������b��3{6�E��(-�(ig��^jKС(��;G*�i�wV�{qФN|�$��a�t��<�oG���2�(�R��Y���Ռ苪̐�k��B[�����o�AK<6ʻ�����J�X�b��l`� ;��3��g���ɢ Q�%1�}�h��ɣ5��ܗ��Gt�#s"d0��mtQ�r���^�a��s�9
ZM�
mR�n���N�#�ύ�;��R 4 q�Gn":��#�I$μ-cyll�A�y1�>8�t��7,��\��mq�z���բ���Ǿm�u��z	�N��$(��w;�n������5t�u+)��#t6ʞ=ڑ}Q��c��\Y�����\SV̿w-����62�����_�e��Q}i7���~~4a��C�J/�^@��D��F}q�~ͨ�
��"�.G���}�Q�<�Uc�/�͗�=��S/�\^�P�A�ͥ�|����lΐY/���)8r�.L�KOq_��^C������I�|E�Z�N�Wco���$���	������g�v&g�p�8�Q3$�I�C�-v���u�Ad���8��u�E��
1�Gx�C���@ �AgZ������E��:�zJVϼ�<���H�>�r�u��K3us'������C�R��'�z�iāy1�J���n�޼����Z"�*�k#0�.D�����n�`� `^�8<��Lq�SC��`G.�"��fHe%{z|3���wS��TB:%pW#��]5B�+8 -��K��T�mA��HI�ղ �HB3�����B�M�'�i#[�3������?r7�*�Ӭ(�g'r��R@:)�D�2l�" ��Zs6�_t d�������dD?Xy=�$;n�S����L�z:$���3��',����A6��O�.@,�+����5�P�!_��4���%����_I/i�Y�a���]_�j("5uW�M'���>Km{��TB��y���<e�eH-g=�^nd(s�����Z��M��b�2b�����a�����g��7�\ b=�2�dM�&)["��'E�b�FT�=I�P�rd���J[x�QZ@sQ�g��H�� ��.b aѲ�$PjI��<�CŐ����Yp�!(�߷�n����D�M�A
״�-"�J!��B��Sswi!<	�W#I"�F������.�!�+�J�Bia�mY�����P�v���[�w'I�jI5�?��	�Ԁf��{�z�ӂ��bK\��V*���/R�K'�,��V� �`k)��f��=v�2��9��9�����%G<�~)������h��<BD裢���@�pG�m������^��!\O�.Z)���m�����|�r�4Ԍ��t�K9���a���%���Z���+=c��!sL{�3�z��x��Y��܎����}�����=�k`L4=�Xki�������$h�BV�,o��%Sb5^����f笒4*<��.��ֹ��
vM�G���V��a��"Vo�d��Hn:I8�}r�K�ڞD�L!v.Eb�V�������d���0�(�{�!߂�� �3w�bF|���Ë�c_z�[h�yI�8	u���V����Y�N����<�����;���ZI<c>�C�I]�K_�T=�2(E+5�¸#�-�l*ݥkA/��G�#~D���r��$���D&���O�o��6��[�����ݢ�+��l��0��1 ެbd�Q��2�2��H�ށ*2�/E�ư۠����6�qLȥ�Xz{�P۷�E@lu6�ƫ����2�\�J�O���A'���Hc�"�$���Î�1\��߂�����	�$��>}��<��'ޭН=a�V/3�N��f�A�E�_ڈ�ɳ9���& v��h��-�؞�"�B�eD�9�I�5���\Z��)D���ڌ���1�_�HK�����B%�>�N�h�7‏�,��^�1H�)�9�|^��_����.ʊ\r|�����W":p�#��R<�i����d��@�~"���:�, �B�M�[j>5��"���!g��8��h��\�/��*e=��0Z�w�1۱��������xI���
`C�{�G���Or��9R^��~(_]����n��r�a�M�h޳հ��,�&�A�+bL.΀o¡W�$ �P�"g�@��;F�y�аV|�p>?�q�)�����9a�VJ`��i>jn�	�fo�)�1�'���C!M���e�?��Q4$��H<y���֑I���v��Z�38��W(G�}�T6��&,�Mp+�6�9�lk����u���"����$L���3�Hr����v�M�1��%�3��W�.0�fa� ��Iɾ�4�)��s%)�(X�7�C]?]�c��`��1�(-&�z��)�ǲ�4�Z��D�JK�WeC-���m���vLb���=��ە�RP��z������L��K��O��bJV���|��.[��9��֔���Ȃߐ��[ ��g%>��og8�� d�x���eP���uo�{�u7�^�|H�[~�F:W0T�㙣��m��E�yJu6��WM����ի�ۼ&�r
���#�s����$Au��g���2�J�Ox=��˂� =���:�L�G���=+��o�G�C��=y܊�f��W/��5����xg���"!7h\B����V��_�	��j-��k��$��X�M~�b�2�%Zpp��t҂K �6�c�xVa�w�d��U֟�D�3�^���ˆPvw*�'Fl��yBF)�,(�V+���m��0�.e�L�J@��!)\� I1ԛ���.k8����T����Yщ{Y�4g�tQ��c��	�鯏��8{��oј43�lff"��v��KI����0�%9�����Mx!0�V뇈�R��7:��}��X���\tn�3i�YKF��/���ճ�}�im��"��Ö�vE��ԕ��ͪ���E�l���4�XWU���/3.B��Cr�a�m�a�'�Wi��� ��j��
��l�0����8���W��9�n���ʉ�v:�\�u�n\��,�P�� ;�4G̥cMi��O뺣cXR���!T�g�m�4z��z�^=�o�2l�$a�/��n�6�l7l��ĉ�l���+�R�w�3r͢.2���!�L�֬�Ro�T�/�X��	'��@��GWL�4�##�2�p���rh�U�H�������(�S��E�TUt�$�J�Κ�`1�/������/I�Y&�i͞�iGmյ}gĸO��L)����G7�U=!z�g>! ����<3d��g�+��^��\~%Chu�t���/C�� ^�٫�Y }�����߻U%$-�'�_��&�0U��9�+'GBmE�x�H�H��	��M�U3�&n�8��u����8���BNs��s-g�}ѣ�$І��8��	'��/	�\
0�$Q?��:�9�ũ����n�o~����٥��U��$�<P�h9������)ｨ��m
|�5w���y�����I��[���~�,����ڰ ��m��Hn�68&����`k��e� {�s�ߝ%���bI�H���I�Q�ܸ��%�%�WA��sX�1�¨g'�Rh>��%�.��}��Ԝvk���S:Ҩ��r�odt�M*$�1;�w+6w׈x��e�nشV*�R�e(&��P0%�h���M��Q��.%>JDK~��ǋ7�ܺ�h����M�W�e�*��|���L��p������Llg�G�{��<���N��of�kP�wv*�N7�e@'�L�j �D���ď���)��L/6|�ܛ)�~>J�@�`~������ˁ��Z��8��%R_iF����	?,�o��W{����<�z�ߵ	���X!bb�q-LTJjka]��ݚ��9��O���㝀}7Ic�y�Ag&�r�`���EP������Q�ӱ'���*�럐'3����-�u���GS˚�~BT���ѻ��ʴ�^]���/�����!.�*�kZ_�&16n�VA�`��h0U���Π{����|�o
���8z���S�:���ѷmϖ�b1���-IS=v�"��?���g�����0���jrjO����7�	�>!�����}���;���d�_��nc[�:gE>(��
�oK�T��
��S�:���e�VT�!�k�S[�3�l|�zq.z��F��0:��ߖ����H�
��#��4ih.�fK�g|��j����Ì|!Z~���;#*X��]F�������l���q}(2��#�����i�ɤf�����?k��Y��ch��)τ��ʓ}`�4�$ԅ-�!C)�\vu����Z��P0�`.��8n�D!�w^F+����2c?�d��ܗ�*TJ���O���1R\�8	=�-�8{�2-\���
�4�� ��E����A�b�$ޯ����LX��	ha�n�
���.�XS�bi?����h5����S2&"�b=����.�z@����%�Z��Z#��/fJ �b�޵�hч܎D.�-'r���/��}0Nz��K�S�zގC���ϡ�Ui�F�	�锼��^�l�m^qo��d��"�4������s��![FE񠴚f���,U���T�+m��u�;�E��Ì��?+&�2��aO=�U)��ZH�����n@��v� �iw�p���#�
�R�q��6&n��jtH�P%��S��4x�Q�2ͽ�c�^GRF���de43ib�(�\��\�Ɂ��+�i���7a�p�穯�ET��w1] ���/�`���"q��:qm��?�(4�  �z�MSt�aE4�|آ7�NL��X'4�&p��VL+q4��Lp�K�Z�I=���ױ������`G�;��_�N��"X��}]�2w��eɍ�4���ӗE�<B��3������������<C��O	H�p�:��\���V�װ��@k���Q�2^�)l��i��HoǷf 0+\^�\�Qo�<ԣtz���T�~Ӵ,Kt_`�@"Ԫ�����!hpwB����@u��(��X�@�75�e��yq^�ܧ0).�p�{QN�o��<��qb��M��?��%�6�u��y`����L�t<�6��\�4�y��!�GY���#Yz(_#X\%Q�Ҟ^]��9 �L!��Ό�6+1�Z��t(���@p��P��u�Z�
1d����:)/(�5�hGJ�a ��r�&ܶ���XVr�*�D�1�9�s�g������WǶ�HJ}��b-6Ю�iNO����Д�\^����ZD���5G⼺��i��[Fz�t΁���*3@i������I�Iw�����H��	qY�%�D+喝x���j'�*����q��J�%lN�k���|��
{�9b��!������x�Q�U���� 臑v:1|B���I��b�"��	K�NZۄ �Bf/9���H9Sf��6�)�+�DT����S}��[,�F��/�S���+�h(�����!z=��b�� �8eل{�#3zd��#8��r�W>1��l����A����� $��c8���yu�!�&�����n��Jg;���6R�{aj�?m�n�M{R,�6u����t<��W��s�3���q/�_�� �j��#x�xǛw�5ʍ�:��j�;�ECV��)5��Z�3;yj���#�]��OL�]�a	~�n��Vp��++a�k�>D=&��T����m�� β����̉#�����SN�<ɋ��["]1_q��ic�YL�.����6���n��Q�%ͨY7 N��ǁ�_:�
�mc�[/���n�K���K��h/k�Y%��l�����ww-z1�fn]�1�O��9���V�h����ڞ+�gff8r��
�z?�_X�e��u2:(��?��z�H���zP���h�V�Q�A�[Af]d�8�;���_iSU|c"^⩮/��y�*�V00�`�K��})!'3)��'�&ȧ�HӾ:uS\0��Ԃ���o�Qh�DAI֡��,�:�n�!'�i�/~�3I,�B[
|6`�50�����d��Or/��	������73�%��+sN�9I�;i�����4����E-hQ�����j�ǧ0�H	��-��><�/�����,h�U5�`���A8�dy;<���L~3o����]1�&��
���w �FM�܏o髀�k0hWP	�fw����Sw���� �x�8��d��fy�Ry���p�O����2pU��t3�kY����Fd)i��{��a�Y7|�Z����͛*~�S�S�!��@���i����tQ`z�a�H��*M Q�;����d��)�x:�maK�ғ��aZ����#Y6J|4��؎�.P/
���5\�{� ���'�x�~�$��y��om���sJ�q�.M6�W���]�l�S����Z ��tuL�K=y�9���h�O���jH����Ȝ�j���ɺ�Q�c
�����9[�X7�3�Z�h/k�V ^���ʡ5��`������,v�Ka�b��e�/�H;;�\����EKn�cN�9����f�刧�ˋ'����ꁢ�E%I^���1�.Q�5�֞]X�}%�.�@[Y���5�A	�u)�u?�FpU�I�ڗ1�<$��K�)73% w��Mm��vW���2kKO�����߂�J��B�>c�p��3RT�{��'����P��Y:hp�Z b:��CǇn���z�F /v+���E�j�c�����5��Ng���,p�xo��QH��y���/���*	��%�xpel�4!�B4a���8����M�^ù�� c�6����)O�ּ�'H�����+I|��~�c9�@pBY#�=�`KU#=���Z�Wf `��ŭ�^N��aVq�ֺ>�T���>��~���SĊ��i_��!�o��f&��Э/)����<&.pC���ެa��W&�1R�����0�i�wr[=�(��z��lzs/�n�7	N�.��<Z��p������Z��?�WN�#c�)�?��B8���rmi���H.����e�Mv>��-��!C"��R����W�4�c��Sr7�o�?̞05�S5MF�x����)(�7�DQsM�T��hJ@�v
V�j�a��|_T��:=a���	�D��X�0�`�P�+ o�#�P�Qw�����訌��RI��m��ù~�n��'��{ΜA^e~���bf�k�d�U`D�O\L�e���(��m]r<�SW���C��AE2-�� 7Y�ϩ%%��Y�X��s�X8��o�7e�7v$续=H�|���_e��F4�2s�C��[ �Ų3v ���on&�Z�l��ܐ��4H�����tv��Z���e���D�N"�l�G�5��->Μ��{��m�	=�S��5�*tq��̳�c3@ �X��G��
�A��:ܠyb�8�Y�� ��KeYR���А���tȀS���V����!p~8 ��y\�e��4Ŧ�]�w-�zh
�d��f!gN���S���2|V��7�󤤀sǦ@ �LŠKQy֙��|(/������G*&����K����8<O))1- �BE�>8�/5]p��G.c�DP���!X�4 ݧ/&�i�3^��/hȦ�B�x[lB���2z3�9��<
�%�i���X'�b�HZ��g�Ə��S���B�vѬ*Z�[�ֲ�U/�c��>thނ���ai�N��4�J�۹�A�[��^N�� )�I���ycB���O�=���=��1E��	ۮ���cX0B�I?�wݱ{~')�l�,&�e�$ޡ��+��h7�����F�b!��p?��H��CQ^�{+-�����Q��4�u�p�Wnu~gs^\WQ��l��:d�b�B�a ��bm�/br�$,-�6�F��&��,�� T\��ҭ��Gl	;aq�fb���Y"G��K�I/�4X-<Ց5�V.��}���*Oo�sO�l�Kb�2���Y�N�-�hH���e�S��|~?��:����i�k��՚��LX�2*�Y_��/����������V���-�l��M}>����s��!��>�.ƨb��Uc�<�/M����e��\�e�%v��ʅ��� V
�Sr��/^X�,6JNA��o��SJ/; �T��Y�_�p#ެ�D�p>�.�il��j!㉗�$��"��  *�pi�-�~	c;�z���U����	��d�E�#4�VK�)�H��`��J@�Y"�I���F��3mQ٣Z���m���`lx���;�R����9Lg�h	?�P�]�2��cM<ȣ���g"ز�����X�?��ʀ3xXM����
�pU�`�83��Hu>MEI0�\&�v��g+�m.i:�b��+�d'��;�kA�y-���>�̥Ϫ��(b���`c�IK0���GCq_��H�\Hb�MO��g�o%�/�^�pF�1`1��}�����CSϾ�L��(3���-9��k�����,������V�N����xY��:v�^�W��NAf�1�m0&*?�3�վ��?b�#��hԤ��p\�&>~c|�U'�Kc�V�>�&r<}��ӧ<'�&a�o��9)��@?�"�}T��,���8���m�SSS����4�@`�H�0�r	��k�JR�rdYo�mR�����8AU��;�_ O��2�b���t�$R~H$��.�3�?LQ>���mD�M���79(]n[�X�%/��JQ��� �Y�?���Ļ-q�S�Aܚ��w֨�|	�M��s����k.a�]������$�g*���=������TW�tKw&q�.��,ြd޺ �N3��̙�5d1B+6T�ܖ�6���=)� �E��ߞ����l!��門;]�t�=�>j��|��Ώ�C�,ǃ|��}93��KH��������"���w�9�ֶr>��N�/-��<��t��&G]�F�#�,^�XU1U�(�>]���[�:��k�>�vW7�����p��h���3�7�5�f�ݺo(�SiA�_H,�@�&Y���ܧL�%oK��� ��.�z�+ -�gO*JoN�b�Nvg���6�/�J��#e;E)��@jz+���>�nv�>D`�G`�eJ��ҏ��$�򝈃���Sr\H�~�����w6����Uq59���������}�Rq��j��
ف�����I�P^��61�Ŵ9�;��𤾣j�}��x�s��I̒�p������������]�u{,L��/�0�E�^��MUk9z3D�X@:F�0��6_�J0� ��rya�����on����%́��玈Z��r���W�Q��Qa�R� �V�h V/��HD���[�[HQ��qg	�2彤�a��Lg��RE��x盎!����xeJZ|�������s�`6�L��U#�CL\LU鿌m]f'�̳�������닧<&��X����	>6��sQ��E�����6��Q[kʀ�"����s��ۗ��R��
�`�Zb ��#UY�]��IQ�N���Ľ=�(�g�G��Ā�I"@�J%�SBm�Jx��!��kY,��Lg�x�<�7Ub��	��c�i)��U�x�j�c��0�k���Qp[_܍�p)��|�~�AAu�Xܜ��a�ܟv�N!�����H��³MZ�ӌ�]��Gʉ�#����K"ۢ֒�[_Ϝ{Q*'�7k#� \L뒊<�׃�Cƛ$�����Xs��z��Rz'y6����x�%� �s�ӤK����U̥�hH� \��Z�G>��ۀO`�S�Ԝ�\s�h����ס^zJ�٬D�ee.��:Fj�ǝ�$�h��)�A�?9�X���r1��CFYד>5'U����@�sǾ��=p��z��X�OՍȋj)[^$88nE�ܜ랗���<���<����<��*�کjKHZR�`��F!����[�[-�ڄ7�(�D�O���n�}�?y��x%�( v�PNi-$�f�Hm� �Ų�mb�kiݶ���]k��P-o�ޞ��A��.�Ч�-��P.�!�c܅�&��qy׀r���[��%^ #؂n+����#���q����j{�L�_�ʉtk����Mm@����RCL���� &j$�P�נ���e]9����[�R��\��.��	����8���?e��8 � ��-�u�:�uL�*N͵ 7-�f�O��z�N`��3@`䭘Z�Mrx� ~��R}�W�4�dV�")��{�t:�9{i~��MC=����M×�=���}x@��3NХ��1O��ݱ�\Ca���a���|lWᆮX����gx
�C�A��ip٬�?�:�Ne{�� N�2q(������U�".jV�=50�)���a!��Y�A� �:3)�ٌp ��Ѽ����:נ�����.�Z���˲!1pu���7I��H�~�.�ۋ�оg�Vz�����o���,7v�y,�{�B�����?�H��_�<�UҺ_'��%2�I��ޙ�# ۱��}�l4��r����+5I7�7{�S�XW���H�?���+{��g	7�ԭL�:�|3�"\wp`���Վ�A)!-,�����H��N�X�,cw^[�]�f\� �f.#�G���^�/�\��BB�`�1�YӰ�Q�`K��od�8� �sl����Lƛ?��W�=ɼ,�Bt\�;�Ԛ��?��)�ch��)3A���5%�� �`p�	�9�N�����Q����k	�*�v'i��; ��>ǹG᠟��ٍ��f��#w3,(��ӵ�
'd���mMݣ�R�V�P�EZH������%�~�Œ�^L����R�q�:�*�7	+BR�`�h�"������]\O4Uϻ�Q����E�/>8Bb�X1�Q@~���β(F�˄�Z��nI�=��FΫ�B{�2�D�E�$�����л<Q�n�ZLsKdW�E5rFrH���u'��w>9��5�c��ɬ
��N�(�/��dVf|���MF�%�̖"��F���q@� N��?M���	� �hq��B�N؄�+-"L��c&����3�f��L㹅�hª��ٚ��x�4�5�Pg7�z��ŸF������6��я��V�,Z[T@�v@�w�t���G^~
�V$�~>o�k;��jܦ�z���HԌ3�MT��O}����i������9=]h�S�:	�@v���3<6ˌf�>GB,����h����-�Y�&���jh�=������j��~
�D���s�{!~"����
���L6>�z����tA>�xYH��]/��0\ʾ���gR��'������c�M�5&}!�V������}��̊�!�u�Z6�A�T�@��3����L��O���>CO�k�663�5�d�������9��yƾc�d8h��٥���H7*�Rf��&��4"v�`h�bk�'���b�������6D��ż(dY���wp�b �1�]�𤋮+nR�!��Bv"3��|�M��5|	P:R0�}}(0�`����]ǰ7��~x:�N���r�X��
:+U�>>e�Tv��N�U�8��H��7�u����T�uܽ��U*�|I�r�l��/��Bj�W�ϫ���Xnt��#�Xa���^��/�zX;-���9�r��+u�[ǻ�U�-\Y���g�ɬ�5S����¼��kO?q�h��M!�Y[v������L[���yǣ���,Ԇ�lc�
�RD��ȃ.Ż��ɔi���;C�	�����&eyl�9��xQ�l!�8
Yz����d��rx�H�]%E��d�b�iPL�<��)n�.A���=m�q��r���GƎg̩�)?G�$�	�s�9�ɟ48����+<=±[��r<�D��;"��ǂ+,���U|=�'��w�w�d���l��)8E2Z��`�;�Np<w��(�S�
�5$��su$�uY�!�%а��x��\�9�,��m_sM.㍈B�!�L-�_eCr73҅R��P%҄�mx Y�vj�򂹼����ty�A�kE�B?�� (�3`�y����"��T�T�a����ˏ���~��������Z�ĕy#��E�q���d�u�Yw�x�eD�7�+���i-�|7ɘ�fZ���m2iL��f��х�%�al�g`"�]�k��P��A!.l�O�_Ͳ��]7��5膚}w,	E���w�*���P��]n��� l��@,T�����:�R��:�X�:�
�$Ku����P4@a&O��8�=1�ףs�.�BX�de`�f�l�H��5��-v�����Rz�O߫_�Y�^Eؿ(�Z��0�1�H�}��Y����.q�m��u|J����|�����<wA���%�tS�+X����pxd�Q��k}U�E)R��_E^5L����7�\_��Ugѥ��*��΂NG7�AK2�D���⇨n6��lY6�C��X)m�zIx3��l:���9��,U��cd�@��|ɺ�7)���� lV����@�e��3i_1 O��´��K˂1ouh+�@�5�q�/qq�����I��Eތ-H��,�}��T��pg�����}k>�p����@<m���C�����������Q������W_,h2᦬�����F�����b7�8�Jj
#�oj�� |�ZU��);�k��I&�u1�h�'=����;Mh��c-%�2�)ђThfvl��v��a��~1ss�웋�������H���a#cΑZ�vƕ]Ÿ>��
�][���ݸ���S����$� 'G���ɠ��Ҥ����+�Ӏ�/��%�K1��}���,2� ��n@�
8"��0���J��%���9�I��>��߬��sr���A��moۘj&I �B�1��ѕw:E�h.<n/Mr�)^��#Zt;@�Hz5����t�SI~	ܵ�I�`�?p����*�A�I_ P�xF���� �Li�8I�}Q�x6����F0��'F��Y֛�B�7�����+*�?��>�T��/u�g����a%�MX��ۄ��I�� �#-�ـ(�o�>�Y�iC] kbB?�HT=��ٽ��� i�=�4��ͣ�F��zj�=�>�r�.��GD�z������X�Xe�e�N��$8�f�����u۝�@���8tM�/Zt��OЮ��Ĉ�6RR��c��K	a�i-A$c_TO=Э�U�J�e���%p��{���٫��D~2��}ńaݭ�n;	Eo������?��:�L9�"S����"�}�2��"3�"�{���L�)$P�[S�kx���E��]���"w��Tő��Q��=��׏�ِ���	�$t�Kݒ ��	���l��M޳�-ό���	}Ky����2hr�g�[�{OZ;n�:,�y�>���s�j%��B;���y�e���U�z�-�_sD�L�A|Z� zf�HĨ����N��_S-�;T������aԢ;�ss�wư�j��G�8N	���[fJa��ҥ�>����$N\�'��e4�:H�_�,�U�������=|��L�8��pC�-����B�&Ӆc\�����"Kdj�iC��V���X���6 �P�� � 5��®� -;Օ��v�Ϙ3���'ˣ ��-�)(=`3�Vd 0a�įI7FѤ�p�;Ԏ\APa�wĞDE�3�ѷBI*|��EY>W������ �Y�Æ�h�=��>�䫮<�G.$�=�*!�� &���Tȸ���(&ZcFҰ��$�")C�"7X�ٜ���+	ǰY,��������v'�2F:=I-�؂ GXD�����V9/��s�77��r�:�V��I��*-�4$
��tiWב� BR;*�c�mX2�<�Ȁ�K���5��0tXS� ��v��X��x3些UxuS҆<�ߋoF�u�:.B�?AO�⇘�q����+g�ɩ���ȴ�K�T$�>zd#��EÒ�SC�'����س	g�?���.�#ʙd�����T͇���6|�w	v~=�	��|��%�#B�-6C�E�q��rҠ����zY&K���A�RjS����TE�H��,O�jņ#���!�w۔/����f،��;����?�y$�N�5��P"T**�a�޷�-N�R��Ř4pG�dF���'DDA�*�k���0i���ȝ�)/wN���'�%�%q�ٚq�]�odu�,�G|��T�X8�e�Dz�V��4�cl.X�k��:�C��)JF�y�4v&ly �VΤk��q#�|�2��兙e2k +]�R�<���$V�.�,]�
g�I���v�Au�Ę6$0� ��d�=�kJ/I�G?��n9���G*F�\k�����,�j�"�������c��}FǢ�H[w��~�*�+1�+~�ӊYsO�VՉp�pF�Β"�������������y��${)�����ͯ��<j^\�tI=��4o3A�re�5;�î�-��n[+�,�P�\c.AX/؉�����=@7_-|F��(��rjڑ�����ݬ��~�hL��;�5�0�u)��FE�:_����?��Ň��P5w�U����ܦ ͓�=$(09�7 R�¿�~��\&�RS쇔x�z6^�k�&6M�`g�e���33�p#q�a�'`O&�s�GC���MH�c"n{6ؠ���n���l��T��>m{Zgw���y=�tG`n!xwH����<�М͕Bl�w/{x� �=������d����˘�ʨ"r���R��%�����������7�M��g����-���r��]�����.��ȮI�f��O�/��I��apt���^cZ�l�$��7��v2�;2A���#:e\v�Xg]��K��Fc_����BmUQn�!���N�7�X�["x�B��stnG�m=g%<}�*c[?��O�V_�$[�̱�C%@�����M����^�7P��J����\��4�g<�dα V��-&��Z��lM�^�C�!�f�B�*ɼ�.&d�,I�lqޢyY���1ȏK��w�N��4k�W�S2x-�o�	��mZ�H���*�6N[N>�3���ue��m�7%�g�嚤�H�3��캈&�! ����W���p�4�r��]�j�B�S�yN	���E����z�,q~M;WJ"�rc��y�yZ���X25��(�q��h�b��a��z,�c[��K�k�-3�2l�����ug�ĭ�|-�U�A�ɐ��U+��S�|U�y]���^�&���Uو�+M�v����y&%KW�r�>���<���H��A��x_m���7�v�$*�S��}L?�ஜ��iq�TeGW�;0����R�o�ٵ�-�f9M�Nc�-{0|�×�>��1�ϼ�;�.�>Ӛ��ǹ9n$�B��-*��),T/z~�&�)��	����O�E�8�����_^8�3�3�0H.�C���u��£6�=��/?gY_�����4|���/�ڳ�����+���7�	3q�2&G�*���eJ��H��-�K�iKhY�{Xbʊ������8�TW�#Y^�����R�@�=G7S��	~8L�h�P��⺳;K`5�c�T�3M���
�[�6@) ^t3׍ŧ��t�+��r�4��f%��ʱҏ~r��Y0�/9�LJ*^mZ���__�۳>�̽;����aC_w<ʡ-����:t�G��g�������cO��sBls��A��C��-W$�����@K׭���m3�g�A�-DhX�<z����n�V��6(���	1�DT *"dg2q��%K��D'L4�l��5_~�K�� �p����b���\h��B��J�����t|�������d�Dl�ת'��j��ò��w'ذ�~PLQ�?�a�����!K�2>���������J1ؕ��|��ӭΎ� 
ƃ^PHU�]��a��#�1&Tqo�XN�\��/����:Ԑf��v�<׮>��bAM�K�M���:�|#>d�f��;��+ϣ0�r�G���rSIC<����F��5jI�}�eC��j+�(���cE�Q��.����Tu#�(\�nu=v�-�Σ��Y�ND/R�G�?9�����d��@�	���.��p�v�UC82)']�3"�N3��� �4����!���T�ұc��1#�v�H@��9f�jU[,�d��x�7/���m��vԈ�)=#��J0��:I���&#6ܫ��n!�Y@0Zbz��o��+�`Kt#i�י:yWaΤ�(؊�M��!��C��S��`$tfF&%(�ķ�<�衏J��/��5�9$��0y6�Z`�Ry�9��2�)W�`<�;TZ�[nO�<f�խ$�_z#��bQ�D��CtN������KT�>=�<�_Y�
��m6R
��ߝL��ƬL�Ν�E����hb�e�5n#���%#%���=��R*�y(�����d&o&Gn�
5��!���$_M�
(O�B���m��JB�~(y�*��ʅ��kliۘٱ8G��VV]RI�*�v2���^�C�L"�?��:�M7�V�w�闟��
V�(F5X*_��/R�$�Ŧ�0�؄�9�f�o��˟�D�������G+7�s� ���m�ՙZ\�a����l��5 iw�F��7"�X����~QO�/d��uu���L6�f��%��亷�㾔+]����^�=2.XN8��?RK
�?H3<�Da���|Q����͞�\��""�C��C�C���O��s-ͧ���Cm��XdM5��� ��>֥�j���8�I�[���a��ؔ½�^�B>3����*L�vT��+���l��v3[�����.�p#�"�psxq��ɔ�o�ß��a��'Y��p9�)\�p�f*�V���. ��A����s
�~���Ү��Ҝ�d�����(����z�Y��Χ�i�H�ցU	��;�}$$�)����1n8��ʗ`�N���F`Ϯ1{�&�{���f����Y���_��]�G���/��*�����y�~���;Ǿ�\k��qLn��qYI��P$R��܃��L5Y�)_g�0M�F�E�:��B���_w3����)$��e��q����k:���{�y�]�&ߨ@��Rx���.��*\�|��h3^��'�1���,HoNXۀTp�z9=�,�;�IW�\' '����5��4���6����4�w�^Mˉ�@��qzV벞��I֢����Fԫ�zt���e��n��a������!ꠔ$���h>���1�-M��rV���������eܻ�U��_şU���3�,9vWւ2�2�:��S����m1��>�Is��n��U?�3��VrޭfE��-��,��%�m�E&2��~��ͅ��
�M���|��OXl�*U#�ȷ1��� ܚx܂���@��){�khS���Y�b/-=	TN*5�t�@�lRi@t�(���*�-%��m��̆v�qc���u�Aa�x�h�"��
S�F��V9������yr���3��kʗ�z)�NI��o ��t�=&��ȼ�:�`�0��g~���]�4�)�Wn��"�n�Y�f'��X�s�X<w�s�oٱ�}o�t������� N=�i���6��TXf���$���	����������%�>NP��J#�ـ�;���~������R~TQ�u%O������cJ��(�B���`���Ѣv����X�'�̂�fO��괭�s)���q�[v\v�m�����#=�<u�9m�A	��|`~�bC��M���<æ�b��Y�]nc���1�]�T�6��͖s�3u�g� J<�;���IAӬ�r��R�+�U��~�m���8��E�=��f8��'#-5:NI+�^p�_w@���D�Fpޘ$\���t�xN��L�<p�5�V��xF����w��X`R{J�8�#l�|cG���N,
S�M;�IO��Z����ݠ-��ƥ�y*��eu��IT-���E4��E$ʙ�ASNE ߉��C*>O�u�4���i�X7}y]�_����K��OQ��}$�D�?P'U�V��tC�Ɏ�N�8M?PH@�\c��ǿ�MGd[�6&�˝�CA�ZU7O���h0_�%����t�S6ɣ�mߑr�`/�:��:� ��P��^�rc iPoe���PQ��씆K���!�K�3��'�A�0�q�ϕ�-��s���"�8���*���VX�@�?=�Ϝ��w^���H����:ci�K���]~ְ��/rILv��U��烏��_(3+�����＜��\�4:y���ǟ�(�|7�<"�@�2eEj`@=��7������G�6�
�s@cw��D���'.Y�#2ւ_�VF�)π1P�,(��XK�c����(1�V��2���I��y{�1j
CM�vNʇl��R��P�3gP;V����l9��!_j�����h�p���P���$�jg��RH20�-��ROӊ�~7�~�8���3��NjX�u���xAY�Mz�#:�v_�~)8&�r����������j}�(�������t��8���L=�o�I޻�'�-Ԉ����Jn��d���G�����X�z�H�)��MXR�0��nN�4�êq��.͂� �$$|�~������,����e6�-�z
��a�]Z�_~Z6w6����ymL�.޼�.!/3�J��a�B�Z���kw�����Z�e�����Y���Sf�3-7�ZK��I�W���}�X���,�'{�Զ+�Q�Hɨ.pC
�p�����&���@�6��W��!�kĦ�����5�>cN�Q�P1R�&�x"�co��!��7�*��$LH=�!|���o�;�E�ĝ�*�{��\'���J9�"؍����Gk�.��V�;Ro(/���^3>Q
��V3�S��z%髇BZ��{��N��oI�����o��v���Z���?��卾���X�7L��5���>��P�Ir����3�n��v���&t�A0�����ܦ���@Q?V^b��t*o }��0ƠΣr_quE�cP_�n�����ӊVAq5���:�LW:�:�p��p�:v!r��3�[�� 4~Q���ʹAUIqŧ[٨�H.���ֳD���.�^��{��m�w5�W烌/�R�_9a�'��'RT������G�Bڔ��8�ͯSF�EIs	if�*e��2b�0�a������w�a7}'��3�'9�s W��@"����}�
�L��<g�9Ӡ�ZWw�9��'m.��'�AVj��a�	�%XIj�n���:�6��tvhq��
�Ԋ)����q�X]'�=s��g�������5���<�ۗ�9���I�"����������r$�#w�b�qjV��E1��ݢ�Ԏ5q'�w�d�\Q���9�"R����v�_�0�f�	�3䉬�\a��b�� �H��@gEi;>�N���_S�5�z�����C�7�דqR)�v��z�pf���<^�-��R'W�)��w�h8uzg�a���\q��t�� �S�Ʃ?��"��U�MWfuΙ`%a5E���B�YY�H�6Y溣ŉ�#x�=J�����^u�3�r��k�o�ma�HL��8+�|K3^�2r� ���*%���a����s�����> ��D�Ggu�����1�:���ȶ�cܐ̡��yF��o�*8N����[��g5lU#M��R��AAdHT�b�W>���S��ܿ�6R����1���� �]����ԃ��`��W�����;Z�ڱ[h�mF�(
���Y���\S9kIL��?:c�&�iE�v�����]�>�&���k�(ۓ�'���ԡ G�ױ?�h�vךL4YgĬ�����s�G�Z3�q"ۻsҎUCbkb����;-���T�9�Ǯ��F5'������9�w�(�p4�#H��;��D���!�'u�3(�Z.���D�]���2�g�DA��=J�m�,�*�_�ϸ����!��_�Mqx��)����!��C�#??bp��ӭ����k�A�� �8��|z�iȹ[�7/�m�~�U�P��hK؅F��X8Ә93�TJ�(��:Z�h��gC���/e�?@�
�Hܕ�`م�o��B��&8�8�k��$��F=K�P=�:P�pv��Ҝ� :9.��C��]�QoY��C��� �ql���[�{���Uu)�5~4 �2z����z�.��uε�AN:�IRω&�,�X5�!��k��nR)A���HxjTJŘO�fS]D�¤�a�lG] =��G!*��KX�eLj�E�E�ʆ�a�df���y��	ne�Pw���T��M����/+5�O)Jp��{hg�����F�fz�?��<��Fʧc$7L���:w>�7�]�u,|� �
=��9�1r<�A<�u�X���䴿�N��S)jzƓ�Q��o�G����q��ͷ���'�� /B��OiX1�*@�c�oҠ�۹ܼD;��C�P˫��"g���}�-W*�H�d����t�IVxN��EC��J�����\�Ӣx0v5��1��[^���-������ݴs�84g}��L��)L������exOc��t�U�����j���D��uZ��:���i�!�be�CFs�-���d�OW�$��lK�+�|" ���#��s�	�+L�)�Q�j0���n����e�`b���č��Sx�J=��H蹎�d�z,�N�`��x]�䦡]�I�Э�|b���}���+�[�oq)U�g���.s&׼cs͛�3j��</�f�K��i5�F.�P(^���������uO#Z��ڿ���>u>oN��8%���>����%�ź����
�X0�j������f�
*qC���i>��K �S����k�8����p�n��`"f�GΠ��'GJ����0���%����Q� ��ٺ&��#�<.)�Ŵ��rQ2�q̷�� 
�O���D'!�����!	0sË��� ?��d֚>���_|X�_9��l��{���!O �ⶢ>��ҷ9<no�V��P�ؓ��̽��l"lX0227!6J��Dݮ�^��z3�p57g�v�Q�{0XGjÉ%�y4�iX��ρ������7��s@�WSg�*�y���%��W���7��tqF��5?��e� � ԫ։������.��;�k���!8׬	�d��=Ӯ�L��D���z粭F���G�Wx[O�`�T�Ȋ|&��`#=�n�z̊��8yi[�Ӕ[��C���٫�ޒ�-@:�����t�h`�I1�-<��4_oc�����&T�R�i�yקG)����0�$ㄪ�5B�c�_O����x�SId� ��ĵG�Xg�x�P��fp"��{��'�@˪<@P X~��ņ��W�<e�� ��f��xQy�D��3Z����)�w��Ha*N�{�/5Ȯ>p~{��Z\�ؠTW�A̩��E)�;A�g�Q6�:r��7:s�=�c,<�4��ˑ�:��&XGk�݉�O��*+\-;�t�f�N�G�̕��q�[|2ѵ�g)p��+T/%7��c����KsP)0���
�hm�/3`_e)�����]U۾�-����ߠ?�jq׾Ҹ�bF�ޘ/��&ќ��'߼� ��|j���ۑ���}ܒ��[����Ix4n�$w�����Ѯ��9c��]í0W�4=C�p��0�����2b_�TO粼'([�@�(+k�hY�KdA�U��W���~�;���3歺ݒ�R��84@�L`���m��*��!��8�/��'�Z̢���MCkZQIA�M8ֲxA��Çc"9:�k`X��b9E���ȍ��g���|0.԰g��Q�'I�d�,���n+��/j��1B�J�f5M�����L,�+i+}f'�qe�Z��
k�`z�';r��Ak������K����l��I��yM��r�3������2啳J���EWX����O=�|I��GMc�L9���V3J�\:�2�΃i�P�/*��I3�����w�dQ�c�7Km �'��n�O���Q��i^ć����yEp�����@m�m����t�Ԑ��i~1r2��!�\f n\�I�s��ç�W�&D��u	F����aƟ^��#��,V��VTk@	}���A+z�~o��5�Ŝ�p���j���`i���Z0�v4ZYC��R��Y��T����"V 4��雍�3��n�C��
FA2�G}4?}�����we�rS|�֑�D]�t��
{��²�|I�G��XFw��<%��l���剺����C�'}�1G)�a/_�f�R���~=�Ti�ͩ���U����u�Q�,d*�5`�/���d�:�$8���5\���I<@[���{���9��(}��S`����l ��I�Yk'`o���#�<�J��y:.��w��L���3��L*`���ǐ���:��23��2Y`��֟8�vsu��Z�4����V��M�����Fk�N=,�ܐ>_3��wv�s�u�ּ��4o�.��(lJu�X�����394�Ɂ�6ƷTX��d: �Z�o&N͟Q�S�{�3���0 6/c^���1���6F%  ���/Ʒ$�|{
�k���W���&�$��ƙ�٣����࡫�m6�a~)�d�E �+�P��#��(�Ѿ�n�n�޺���+(���k�N��J4L�Si�&G(����1�X�q��!�al*��588ȓFQ`������H]FE�\��O U���(�������MR�F��'DO.��e2�B�p]-�"	�V��L\�+���6t%K�dT_�|Iʖ$���ٔ�e�j����w�.p
��{���j��:`����2)6�7ׂ��:k�����)��؎zh>AT��a~� �
��uԆӯȋ�B�aw-;���o�>�w����R�#�˙����H���/���R26#��)\��:oյ�T#��L\ۍ�w�KQ��&���Cu2�e-��9�>�x*�B��$�ƅ2ǜӲR������&��D;N�D���y�E"j �b�=���$�\E��[E.Q?��%�ޛΊ�s;GO�n��*��AZtY\�Tm�lL�'8�^6%��?�v��/+b��v,i��y���a�������'n4����/�ݍS�G�@�{�
Qt��w�Wx���������,���A���n�J)�_��]V?c�X�!c��mp�'��ڂ���j!
��Ce霩��W*�:lӞVB�N�nMnjF�sɞ��&Ѽ����Ճ^�v\����.�g5j"|	���jS�
\�� ��	T��$8����.��8�m��Mub�-�PhYSG����b��S�x2P�
B�C6�����9��dga�Z�D)���4*.��!�V߃9����wZ��cפ�H��HFŎ$Q�?�'{�����E@ޡ� ������3���l�|�����7�	[�2.��Zr�t1;k��p��Qu�ye�F��gJX���㑯��bB }A��ǂ�`O���!���O���}V� ��qz�I�����[��~q=��ގ.��&��J�@/���xlDB����0g|W$6��K)�R����d�A䓀.�E�$vM#EjH���3K�ꙣ�jX-`,�v��f&5�^�|����&��?��a���nY���OH�K�i2I���}�߆�JNyR|�f���d���F�}���6�4r�g/�����#��W\����nJ@|f������񂟛S8��~�$t(4�@��uԀ{��?C����� ��n-�4������X7���_!�����۵��=IJLZ�X��\P���3�u�(�Z�eMٷ8杜��
�*G�׮�U4t��f�֩Յ-OT�J��Im愓.�����"b:���c�04�ќO��l��X�'�3\���<�</w�@��dϖ��N�u�V�����+�l-�x�*��yY�`U2b͘W*\gӽ��&���ʟ����7�y��������d�x��_��/�M����{dOGK�|�"&��W�j$6#:c����:�+�l7WO��N�h�4r/��Yye��I�<�$�!��HKx��F�9��6q*_<�#1�"fi(���`��C�+ЫՎ��SX�Z����um}�KQP�O�w��5�s�@�J���'(�QB��0Đ����l"Q�HG�bD�M���*��װ�S��}A���b�e���-�#,­��X����6�v��ė��IinͽE�Ώ��|����;��7��b�1�v���ŏ�� ��(V|�W *�nA��K%���%�B�9�DdTx>-���� �B,L�)���wi�˳�������:���c:F��+@hs�d�x�84MS�6����K�
2����!��r;b4���ع��Q��?\H%����)S֪2tu��Mm%m](��Bܜ�-�hj�5	;�._}%+�z;�"�{ ͑l���ǐb�ʜ�mެ��G��.Q����(6ؠ�a_��aW�GfE�ny�0� �&2�Pד�C����y�q}s,Q��T^Ǆe|$�P9��U$��b�[w��9�莥
�R�"��q��>���`�{���k��w���l[2�k.�����-}n§ύ�˘�<��;v���yH<��F	qvs-r9j�����t�y�(�(įn)hѼ�s��w���2u�2�4����64�-^y2�gMiG���v4N"��S���83X�,��^������CaI�=>;�E*ҳ<v�����ta���+�R�Ih��D��h��?���3��E��N9���j+�������1
ۥ?Ms�@9�r��y��ݝ�b�� �}1d|
�!>���]>A1n�4�>�X~�>�E�@��_���I'+����zg�$��=��ѫ�:�n."_r�W�e��'c2����?�o��yU��2WP�8z�ȳ��� \Hd��"����xso��Ep��[^�&��)M5��u-���%9�J��t �����?½5eYmYD���d�Z��t����s!?f�S����c����6#k-=Ⱦ�] ~����7+� ϩ��� ,&N W�Z4+y�žoH�πL�ms��쯈�tI���� $Y*֑O�W���`�PCD'�$R� .��R%��P�`�Q�%Q�#�s&���CF˨�;��N&��e�����>�&F���U愲\����e��$���9:϶>%�C��۬�ψ�%�Ò�A3O�0]��;W��/z	z[l`�B��
wm��i�\�j��ί�j�h��c��%��B���%of���xsq�IQB�,I���z�W�Np�H������Ҕ�d�d	�c�#ͺ.�g�q��$q���>f�/�P#SĴ�������\�*?��Z&Rd����
������i!�\�H)���x������l�R��E�޿uW��o�V8���	T���,2�[[K�'���%�[�9^�[1���w{���M+/Bؓ�b�`���fh��Ӆp|��F��&��3!������,d�'�\�4YX�<�<�B�+>#m�Y<����J!H *į���9{�̴ڻ��̝� �!(�9G�.�Я��g���:߻4�t�'{(��p��X��{L�&s��7��=�=@���j*�`Bzx�(T4��qSex)�zӑ檎�T[�7�A��-e�f ���5�Z�([$��D�P�b�y���Z,@��TT��1v#�j���	���/��������&�م�Bפz����@���������4�F#�0Kb�z��߰�?r�T8�����p�˖dO�Y�&��G 4?�ŵb�7������$�P��m�fД�#Þ42V$�ԝC�A�
|�<1��z���տa��t��Y����`���`�f����z�61���3�VNL@X>�nYm�RgV�O���I=�Zngʚ�[���|9���N��_gM�/�	�k�(�}�+Gbɮ����Sr6d�W��J�y��M�B�Y>!���[m�b�ؓǀ2p�(qF�oD�yz����������6�S��PK��æ�B�U���U�����0�/��C�
�5����ݾ�$g�&E7L.Z�M�E�:N�K��vG�{տqe1t2�s����\8
+�:�A#8�B�{1��獡�@b~p�&#2�bu�����a�δ^�q+
Rk� ,Bʋ@�Ǳ��v�WG�NsYA_����y��M_�⚨q#�6`aĞ��xc.�R��N�90.p��S;e�EJ�:����MK�T����X>��f�1�L��(?ɍLUR%W3�x���n�j�n{V���U����ʁ��KAr�|;�~������@d�9�Q����d��3��3�T0��� UgĴ��y1��d�G������2JU�@�i��a9#��vAB�M�+Y9?�8-�|�l�܊F�5�mo�; t�q���`���40�@=l���4�F6'�є�7���v�\ӹ[�������d 'N�������1����r��#9fZA�f�R|w�JF�wUy�#
�B��7B�ߵ�D���b
�R��93;��
N��8�7+��c�I��b j$�P��v��D������h���1�e.ʾqh��	�CQתB�q�O�D���C�l�W�h)��߇]_,xN+*�T��?!0�>qQE�W���L�iǯ73��5��Q���<���A1���������~he����r��C+�D����Ŵ&gKB�gy.�U���d����.�h�#�����ƴQ{h�+씂�c����ف����M`������ zT���;=��J���Ͼ�맑�f��*�����6^��O�>����-E%��]:����tȊly�&d���[���������My�!�OB�X�$�!z��I�c�Hz�~�D���U�~��v���҄���d:in5��}�7���]���`o|�#�2	�K�Q���&�Sbr��7�{�L�a���3@2�Me���l�m	�o>k)��{<�/�q�O�̽�?�c�(�ykCt;�&o�`��+;�������k�Q�%��,�CJƇ<��{!BX�(ɕ����B�М�T�S�n����X�� �-��i�Bz���I_�(
)W����T)>�1�ڞ���ؙV��OI8�`��s�'T��*}ag���c�+h��<����W1�.�!c$J�[��A�������`�0TO��L����g�f0�i���� {�$-W.���h?�t��!>=c����Q��<�����D*�a�n��&_%3��=�9��`�0�������&��"ҭ����u���Z���^���aC����	9ҡr�j�f̳xU�i_�zPU#z�����x��D�m
"̕.d,����4F?�UN�����!�oI��A�v�%E�O4�����W]����>\�o�G(�r�G���
x��ρq
%���NP`\�����>y�2�i��������bs1�B f��(�LW��B�>$��u�9���薇0O�� �X�0{`]�(������o�v���Ɗ��L,Y���#6�llj��g5IH�&.l��88e�k�L���*������O�b)sd��tpLD�{1�GRD"��.Ї�3W��'N^3t#s!�}3�أOH~9�������P��d�����9Y<�U��{Lf�@=g�����Ol6v���՝Жv��qB��w��a�*W��j�Y�֟B���Y3�z,xКm�lu)s����[E�@F�)q~j�L�Ɲ�2��߿��T�q/����Np�G�ԫ}�8@z�G:��f�2���H���c ,���؍ᥝ����)�{P�������U����/u�4�=~��@IgK}>���p�+�[����e���4$�W^���`���<ۼޮm9+��c�-��0о4Pg�`�8�L�	�8��<g���[!��L0�Eu���fW�����|�(�����T�ΰ��J"#�O6_c���I�3�"��WՂ=8�<��/�u���}�wRzz;�hM=(/.&h� 2V��~��m�ڗW^�n�!U�)���1^���#0?dEM���^�.�`�&�:�*	�����f)����.g�7ǈG?�<3��ç�n=���W�{-��x�
���/���dI[�H0V��A�O��e/�����|�b/ȍ+�~;��⦧���{�N,u��%���z�E���AHz b�^���o,�Ώ����Ѻ��H��/6��J�J�X7ȅ)߮Eb餖���o}wܕ�'��"�
\ﶰ:�?!y��<w�~UA^�d�+��j��谁�R3;h��TT~�siE���#X|f����u&{stk1"ĽXc���"�Zq�7��׶BTI!���\������pf�ʄ���V�i2d0���Ko	Ц�._�E )��%��7����ޮ�����C���BYSSuX����!V�vV܊2F�ik%m�3UIF
]�9��(�s��� `�rQ*����u��G��ϫ��
�{�(����(��D{-�N�"����e��5�l��g�ހ�XU��'�/�v�����[�)
z�63*�J�+���#s�"��n�NËϭs�|^g=X��tj#��g~R�^��t�i�V�/�
�.f���]|Lˈ�PZ����
"�d2:�$�*�a�K=�Дũu����� ���:�-�-�+��o��a���L>����-� ��R�7����c��f��22�+��v��?�%"�ώ���QN?R�_r��v�q���Y	�M �Οע��HQ|�7� m{U�ׇ�����<�O�,Z.��e�tb�^��˪3��1i���	bY\ރ���D� �G�W�#�l��)Ɯ��sj�A#��PV�0�Bw��z~��zT���)�CyJF�ǏP&���H^zIw�����2�����*Zc}kL�ݱ�J7��ZU��<���a ��� �YAY�F:�x�2���)E3N�,��椉�����7ӣ�a{aCQbH��&��P��w�����E�z�F�Ϣ�q�K6M�%{��wnu Lt?�2��#!���?�~ZHA1�u�r�!�Rr~�Wq��������+nY8���v���I�Z���D���}]Q�%V�����؛�-��b��D�0x=z<ѡ� �f@{Ԥ�A���Ti���s�k��Ĉ��n�^֯��	�>\:�_tk꿏+B˺��31^�{�_�`L򙡫�edD�V�wѮ�fNlĳ똮3 o���`���,�md93�QY��(׈�,S8��A��1�-����pa� �a�[��/�C���<��B�B5S}��fQ�����ëf^
,�bF���� ���3�wF�4J��Ճ8�2�|�������a��!�
zĲL���ǯ`�����HCm����ۘX�h�K��4%�<σ�8�E_/�b(�ɺ/\c�a�E�B�����
�`89�鼘�.�0t���i�i���h�G4�,hR�-��c�����x������)"R��[�*��/���fB�nP#ʢ/����^X�6��s
��@�!r=�q�Ӿ���Y����~l:�g�s>�R�C���-�	�+X2�����̂,(��8vVSI��r=����L��ڱ����?�)�]u�9 � -�>8jr��P�V򬽮�l��/duV	�pʛ��:��IIBY������E��P`�*����vw�L�ȵ���H�_���� a��l
O���yx��9&3�z�-N�r�WRu,����*���A�Aѐ��8#���a�����"�DH�<���#]���V,�H$7M,�x��Z3��|L�	�.�������B�7����G�����X��zSu��ܬ[�Y	X/� �S�����v�r�+�P�'��k�c!r^0#�!���Q�
ũ���	�t�Y��=��Ѓ�SxQ.IX�A ������~�9�N��z�_�*��I�m��F���e���x%�߷��?i�i�m���.o3α��~�f�����l�!pt���B�ge�'&��u([�E�x�}0AOo_f����u�GQ�qf����T��d�^1!�
![��~
���<G�W��Y��Y[�.���tǹ倡���2 P�������!F�����{R:Q��)f�P)4Q=}�jr�����'�T2ׁ�~���<L��ʖ�8�=���'�k8��:g! �*o/[b�CX&�I�)*�Q�<u��<R�;?&f�d���Z����1���q3��z��;����=6�b^h�J��p�|��!�������K5���Q�wˡ�6A�����ֳ��� Q��K�,������(r�u>9M��ɝ�ɀ�[�ݽ䞐��=�YjƧ�L�J��uv6�Xo]7
dqD�IkQ*��}�͹P-�wU��8*�S\�3��V�k�C�'Hз��]�� �v-��/Ȉ~%�e�
w������3Ѯ�R;��HUF���h��QӮ�Z�+�[e�ӈhDJ�x��Ho}� �����SQ�&t��WBK�f��n,�;�=��*|4�PO�U�%|k��6p�k>�e����5�i�9�;^2�<n4G�����c�h��G������8������3"��lFБ�<�O 1_�DU��Z�G� �*p�6���_��ޜ�0Υ9��Ԣ����w�����B9) e(��T����?��T��V��g����8��K��˴QY���kHo�}C0QUJ�r\���($��NK��A����w�ye�!N�y�K����іi�E��&^��[`��Q]c�o���W�UՕ��=��K�BR�����L�f�y�_���8fY]x{���l`��j��?	6�u��*���>�gtH[+�Ǥ�A�O�T��	ו^��`CY� 
���2І4���g�x76Lt�����àN��mr��-��[�)�:2�����c�R�ܝ��W�Fo�*v~Y-%�N��t>���g�U��˹Z{s2�O�\�G�5,��<���"tr�YFP��U��w�!�-'�X6�&�S*��Y_=�m"����w��A_�ew������C���F�Q�y��Ƭ�*0䧅ł�����Q�`���*��?='x9��r�jhj�{J0ݗ�/�m�^H&ݚ�)R��=�@u�q�2�ۺ��.O��g��F�H>���e.	�\ L_~ٱ ]����J�&)w���	���l������
��,w�*~p{Im]��U���!*�B� D��W�Z�i�`+=����[�m�!e�CUa��	c᥉�<teK�\�Qwa ��R��.ƌ�G}����t�usn�@Ew��z@5.�|sc4$=�5ϙ�ge��>�|������8�*%�K1��]d1�qs�xQ
��ʐ�E�+��1����{	�Wq]kӮ2o����蠍
M���m�tl}C�h}��^߻�h�Ͻ	�J��~Æ���E��W�;It��\���)j�_������v��zqwso�p�OH+�?TyaOp��6���(��&�	S*r��d������Y��iYҵ�	��e�P6�i��h��sؠ�����w�H]�w7J��E��D��F<�ʼ�~ދ��U'��uA�T�;V,֔H�p���NS�<Bo�p��z��?!2z���Y��xV6!xw�l]�C��n�!��7I���a����+�2 Um̓��ޠ8'[.��1���$�̵�p^2�*�Qi��%kz�%8dE��(�3<��U�a��S�"��#�.�#�5���(3���}����TG '�q��4�#{Y���)_�����<���$�y����rOݡ�Q����q0�v b�����&DȾ���_i�9�ä����x�1^к:�6hEN���Sz Αٮ��e6pҪ�e��[)��B<��h��@#L��*tr��,�/�_&+��0Ba���?��6�iU�������&���IZ��*��a:�H� �W������S�ߴ���o(ʫ�lyGP�߼~#�r���(�R�|���k�z`�6��������ϖ�)�g�t��8c}�1�u�5"M��	��o�	)��P�����U���WOXk',8w����!�14j�P�p7�3o�M�t�B��:��}.A��h�4E��V"�MVI�-1��a�AlBл�G�vt�H�u�B��?�,�ӓ��i�X���8�`V�^�#%F�I�Ms��\����Z.vj�ZsV%����� �C��~��(�4��>d��Û�޸l�f�N]�{���d"iQ;��m���,<NdD�EP�s�Z�?Q�#}���<T�sLԩ�QRg��`��G�ޠnM�ͽI�����&��;����3l����Va)�;�9K��tl�.L�U��ؕJv���Ve�b��k�64�@������f�fRd(e�YD~�=�"h�n�(�ӝmYr��9�u�9��ǧ�0�U��4Ȩu��@����q��s�� �^o���%�l!�W�n]�8��]>�*��\G'$��Lk]��Js�t_V�͌����\H��fr���.�ߟ��N�7d����:x<y�Z�2�G���8�����)=}jݙT/0Hg� ^8Rf�kʈV�I?a�0	|���r�g�����^W����o��'�y�����Џ1������qri��f`g@�J���էEF���<�H%t��M��5���
�TH$��?�/��"��2�� ���J�`'}�r�ʡ��oQ����Khrq;�j"��	b���[�o�:h��Y�n&$"����p�K�]��K�����a����/�N�w-g0kN�����L\�d�
��T� �?\�b�������?���P[>�oWT����΢̋ψ���3ox�E�/����^����|�����O�-j�Zb�uB2+�G��ۜE=T�2}�짴W��q+�+�-��5��?i�D@��R���M�7��:-� F-/��rC�H)�4U����J<ޜ��7't�jښȏ�\�ŋ��{E�����>C�2o}k��$o")�
W�����۲��C;� T�r�zJ�˒�(H��
��:�שj�V��+GK��+�&��[Q��N�@�N��Z����s�Lrl��>G�!�E�$����������,�Ӑ�������o1���̰C|��u�,X���jE�l��q{1���e$2B��
���s��� ix�bhƸ��d������h������aǐ���!�F/ɮ)�/Y�N�G��@������L�yY�Eֈ}"��� i�U�Y�T�H�z�˂�	\��P�O��]
�8���%����;��u�k1�m��"╞�d^}�k�[�%�.�Qo����}G���i5n|1(W���`b�l0��S���BM����ME"׈��B�\ј1.�r̛�Շ�Ig������_E�FĀ!cO��WW�|����j�n���R�d��:��Kn	�r���b["���v3%��~�� ��|��w�?=�b��=�����<��}��1z���){���V����F���u��ro\�C�<�e-,��
���u��zt��?�R\�/O*�{�:�E{��:zն\=�7�`�V<0T&DM��,)��!*�����N�$#?V�W&;S���0�m�Q����WX~����j#�N�I�cq�',�kK��Ŋ�����E����NF}�ͭ��M*���O@����|���)�w�@��J�	�J�C�aG��"�WB�r��J���Q�Xɚ�N;?��1��
7�v.ȸ8�v�|�w2 ?Z*TnL�f#�~�׻��N�˸���O��E�3ZΏs���(w�zA	��>�S�UhI��w�L��Ag�W�]1k$�и;v'MD�
Ղ�;�a6���t �p�w�!��_Xk���M�@"�ER\z�p<����9��Y��=Z��;�H_��2Z���dA� �S�E�A',���2Z�ʗx�	���%g�2I��B���]pN6U����U8<��Qv����/~b[ �q����;/$>j�	�
���PY�z�"Q�,���\M?ȗ^�-���hКM�3���L1�Ҋn�N�D�_�s�t�6܋v����U��&������mlFT*�T��2�1Z�V���y�\b�)(�e_���1�\V��u��*�(����Qa�q�`�	�����?ܖy|�Kr+n"$���5��;E���B�B#�Xu!���1����:%�`�a|P�/�ͨ��2��k���u��5��z�-k���@���O�S����Z��e�Y�Y���J�d���f1/ɀ������i�Ϛ5��4�t-��V�lMܪ��]���e����g��Ie�=ScWK��(-�����"6v�Fx�.O�s�<����Q�������Ӎn~F�d�U��Zu���!��s�l�
�R�2��kȢ�B�5�% �ؙ��4'3�f�E1���Jp�
���L8Z0q7��J�U�o7cc�������������uތ`f�#D6'w��+��w0"Y⫟h��k/�hP��S[M��섢��(��9,�:���o �v��1^�.l��7Ma�c�'5<���W�U���W�qx:���$��)�,����Б�{��	K��Y,&����$�3��׽3��8�'�P�\�`��U>��G |�Su��lqB�9�xs֢���m��d�<<pd���8$9�Ե��i,D����;���)��}'�;�5�Z�y.;��qD�nGx� d;֦P�j���)��J�2^��% �PBP1�s-0a߳��hp[3��7�c%�BN|�댜�.A����`�� ��(��y�̼����ͫ�^LJی�0�Y����3\��$�Oo�	��P��u3������%O���n�i��PTJ=���|��{7rӇ��C/��p���c�M�|+
\q=eR�� �0�����jdV[�m�bPn$(�1`��$=OH�'o��j �/���b�R��6�HRn�k�K �����>�7^p^��}L��ͭo�P���#��G��.ڰ�X��'Y��2�v�m�P�g�fg����<"���̧Ϫah8���=�٬9�dCcm=���3�o"{��?��>�nB��2�����}E�l��q"�>���T�����1��x�+�&ȂՂ������$l�%R�k�4�+��yC���H.��څ;�ֵ�7��~����Ö�(|�ט��M��l���h�H��~%/��Vf�����֪+�e�P��ʗʎ�
�G�J���s�Aq�Z�`�T."��eӘ眹$��q���fI��i����C2�]��ӫ��Ex�^3*)~h!�ڬ�f� ��})H�&���V@�V��$��������w̪4�N1L�0Č��*��1���^=:f��H�'��v��"�x�1\.�٧���b�X_��~g6�P�ws���Bs�	���\?�q�?c	"�y����wW��!��x��)G��
���^w��e���/u^�S6 =���:����^���S���%�0�~�R� "���hPM��T�E�; �����&/�b���&U�1	�J@�J��̧ru�$�C�����V�<r��_�r1��-��(m�R�@�KK3Ӗ�K���j�\���N�KH`�K�_��6j��1��K�9Ο�ԀF ���y�u!����P���<�K�*#/X��hY66�N����n?�|�7�gL�s6Ĩ�1�H�����=�n��}��#3�Z�w�˒�r�ۘ�#�y�Ok򵍛_�l�Q4�������)ޣ�ҩ���cS#ؖB��y~^�f����8��е_�Dr���2��eė-���P$	�K���0�7]�sB�E=ջ�~AO��,�P(�����b��Z׏�)��d���Q+�Ll���g��5�uwR��8�c5b@�J?����d�>�0?��ߝ{��?$�H��5SZG��m�	E�����/�#&ou���~*��]�7Xq��卣'��A��gm�������� @�o�w�n���2�@-��5�R��§�6�
�3&��c�STҋ����V�H��Y0�X��t�G~�@78Bf��E=���+���H8dt�%Z�2F�ƞlU g���i����zW����Pƚk��fG�G��~�
�ZM6*�����\,7�܇J�H�������ǚ,��|�5y��pu2X�ȫ�cJ�g������x�g���ߋ�;	5V+�=��A�#
����(1�B�����jU=��	ݑ���
����$�滝h��xAA�:.Fx���k$�-W���_@r�5�k�$�ƭJ��F:C	hnkPkM�GM��Ԑ��% &7Vm5��P����|�-�pY$eU����~\�V�r֮Ua�}-�P�Y���F�Q���9�0)5���8����F���Y7*�q�o�<=C6Ӟxh�Rd]xhf\"*Ey��O�m�ׯ���H,�_t��[�Ю��.���|5EqD�9�]�p��5H ��+룔�b�=T�Id�Rh�S�0�wTcg�c��+�kfʈѲ�.�+��"�+��1��m�$q-�/�K�9�S����>�=ܼ屮h55o����Ǌ��;�޾����)��a��2�� �g/�!��o@�n��v�=��dKp��r�,�j��(���V(�k ���ѐ-	*�Sl���K�Q�2�T�&Q9��C�-F��Yt,>&�(!���&���{��M
����G�=C���^�5�+�3�{-���9���^C�w�g!u�Ux�t#��|�Ċ�7m�4L+�XB�� M;L��GU30���~(�^4��n]&�/&�{d@�,��Ԝ��DGf����g����tc��j�$�,��Iᘺ֒	�'����,��h�2�z�z���U���V��SWW�ԓ����ȩ��b��j.�^�A{$#+��`9@[o��X�:M�y�F������f�c����C��G���������ؼz�}�w[i:�����c�� ��0)'ǳF�V�Vſ�-��$�n�,�J��ۦ�ЇA9c ��1^�1+��o�f�&ҷg����6@N�'��'DH�2	�� I���x��,�^(��,&-�W�?R����U������M�pWV �AzS��o�-�ބ%��h���baC:[Qo©�{e�qk�f2M��� y��; ��M�!���Z�6����a� 9��.3յ?�x���9W����	a��a'X�8a~::�����:'0��s-�b����k�U��q'���<��N�\|�^C?i�l�11L��nE?Mc�S�o�)Qc�1_�D�l���(V̏��.�.ظ�5�@u@��#%����>*՝�a��� m��O�7JKS��Yf!ylh;lhc<��ӂ�.can�:�ӽR���8���-��
��1[K*!W����{�Zv�,=H���Q$Bu)����zΡ��3q7�\j}=��e�X0,P��<!�O�� ��`�"%���?�O������,#�rZV���
M���U��:�p<�N)ZQ��
̕/�>����37Չ3�#���z�o;���~a��-l��C��y���>S��؈�؅�V���/��#1�5q�Ao��nr�9y8��|�������1�y�l�$�Z�_���8:�'��"Qx��V�G�S�܍&�>b~TF�%/<%�-99�U��D5v�Bq .-�����G���o��͘�B6�/�.�q�.�J�n�kTEY��x�m��u���%+��,b�a���{,��I�6o۸S5a�T�)��1����kֈ
!�IƋ�H�RBX&���� cOMc��g���&CJWd�[�2ɏ��#20U�_��c�E���i!�`XR�4Δ�M�ڧ`x��g����M�Π2��*��m5V�m\��"
��d{$��38"̈́y3�e2��riǹ�����^Դ(���zɄ�����vP�*n'�R������2�Y��|�2D�,&ܞ�Va��\6A�5^�aXX�r>5�&	&�P��iK��V��.�����PA1v�.21��m���Z��;�~2�@e�v`�x�Z!�b��b"��},Ǧ�M �c�{[#I1�g�t�5���eiu�sW�S֔?���(�[�5�!㴙��M2�8tӱ5�)���3!}W�V��SӦ��/��6�|����O�hZ~��L�"5�E�9�Et�1u��L��m=�� �}y�lBm�  d�5K���({d�&0ϡ�h'=��=<X˱*�fd�?�����v�Ѽw��"ơ��TM�|N��ߵ�c9/�p;c�i��Ŗ�]�^=U�9�I��Ш��Ǚ�����-�v1���+��B{'@(E*�;��<�o� x���T��dg`e�;�#ql��d-�]����A��u�^0z�F1�v�v��bM���E�ʏ�r:�.�o�}�?��s0��U�f
<B-�#ch�?$�K�D�{�]��=�m+/�H:�]�v�{"���*S���=���2��N�SW8v� 28T
?m<�\��w�~����-��n�`�oh�,X�_D���@hDw1M~w@��6>l5񒁦(�o�]W���Lޥ&4�� Oȥ]L�r\~��p��Ϩ���~;�W��֘M�-4�"&�@E���qB��m�ٟק�y��c�!�ޏD��A�!�M!�a�br�"�9�"u��{��Q�]8-�1����'��5 �|�]��(��Q�~2Qf�K��"�UX�$�r)��5\A���s�s����������r6�N���p��m�ڀh��xi����J�l�2U(�c�*�e�L����������T�9�ѵCO�x���)m�ݱ��頝 �\�R�������-:�[ M���O	h��M���O�F���&���4��5�ֳ�e�b����c�ev���]����f�o�qq�(b�_q>�����UJ�B>���G��ܚ����Ɉ�q�h��](�fkC4Gmj#�������L�vo`1���p�N�1��{9�@>����Cq�c���)�>Z���vͮ��nm�3J$,97�/6�鉟c�+'�De�"#�D��5��k/��y�T�r8�0
�>��`YS� �V�殈�s�Il/��޸]u�oxIʲ��WWd��)�J~}�?�'��-���YG<�մz�I0x�q���L"���Q�A�)��-�
>��Gu�T�ۈ'�n�TJ�}���W0|[��fXL-XL�lΙ�����v������>�����F@�:�e8��3����M�-8��� ��Z`��4�1��v>�)]��6��T6�%bc��'�S�Ұ�V����!XKv�{��w�3���t��7l6��v��t>B(���F���V{_�I���j�+t����y���^�W ߿�vg�ލ� ��Kj�[)����+V�>6�mm-�%f�qXX�OE��Q]�dY�OOK_���4�V;�{Y߀<����~��n6_��Ie{���e��P���n�����ƒ�������YX�	Aq����;�z��!l�D�}r�s|*��������Y}hc<l2DI-��(�3~~c�!�t<-���IȒ�j��Ƌ�]>��E(q�
�q`DR�C5����ǒ7bV���[V)�Qo;Ό�ְ9͗3&z��2�=� �
�E�ϝ��ԑgF~���X*)����9&� U�U ��c�A��>�3�?�u����Z�놝�H3�,��A>�.�A��$�uy�.x�ăK2L;�h��P~��.$���_0�ʔ�c�3���X�@�S^!�"k� �����Av~U���h�lB[����j�P(�lB���H�tM�c��\�౟V2n� \G���[H�ϴ7(h�ٲ�6[�Kw�9)�냉z�a�eF8��NbR����l07
�p ��i54�5i[-��+�v%^x�^�t��SPƑy4h�S)�G�7�8Jrۃ�]"RE #Ct�#���Sk1>X?�-٤��s���E�A5�����	���ɡRw�KgXM������F��a
���W���V\���]�������91<��>��*�а��F�p>�0Fl�	ݭ��-t[���!�ֲ��6_7s�%/(@���#���K��D+���x4�d9;Q\�ٯ\����Z��@:�{ln�&�	�x�p����Bz?Z�r�ZK+̙�^�pz�@�bQ�������e����YZ��.⟎��C��E6�pU�RAK�~UD�RPh���q�m��d�Sqf Gf� ��=��+��|�^��}Z��F*�jAQ
$����&�_��:"İn��Xj�eF��P�\��zA�Ċ�I��|�(��5�fx�%�DC�z+�jы�O��p3_ yya�8��JUC�0�ʩ���>a��݈!>ʨ6ѐ-�D>Qy����˝�*�N�X,��H~~���K)�z�X�7��j����(�p�V��d�;��aY���!�^���>g�i��b�w�ѿ��9|��i���Sxv�s�����m��{�s�&�e	��y�(%39�5-�e�v�(ō����l+Օ�u���MV�X2�~�L�~���K;E@!�yj��{-\�� �w�d���7��P&>�1Yo�A�!=127��)�i�]���<�{	�Y�.	9�ڈ���d0��׼��&���H�����.=�R���A�7�����w�:�LW��Eo0��o� ް�@j�
.��8���C��5:�$��圏��no�q�בf��>����� ����7_�'"�ƷzP�j��&�{f�0���"�j.*�q`�͍��e&�ťjlKa�q��W��I��M�n^��;f�o��ª�c�6V0�,�\0��_���� ّ��@�_�%�My$��&�/~�NQ����ۃ���_j�8?.;a�\���S'
|��1����b/���[x$���l�4���asW��Q���cE&G��Gq���t�����+h��&��;_�/�x_(�]��'j�>��d��|�d�k0k�~�m&���D>x�q��W�-�7ҫa�e&�P�ǛIa?��^l��fp[�Y4�rńT���U����(J7�k�fc��:k��@�!���V�z:)�QY)���c?����&2��<�����G�2t���:�p���
	*�@I�B�	�=��DF��v�~C��Wg$�o���|Q}`�LSw()�3��~�0`�4g�*xGHq��xEG����e,�ƀ`�耮�������=�����Wn�FC�2�6���3����C�+��Z���	�{�]�w�[������ԩ谦�=�8�dN��}\�5�N*[�	SL|xQ�^�v�^ތ���iM�6L�{/�3#Z��"@n����a�'�imť�%%��w��k�g���>�X�̓��Uɶ�U��.%vO��BS�X��.�l��\!������3
�t�o(Յ�A�>/%1�AGP/���{�J�t�m ��S�#��k�Ϯ!�o��=�#1�|�is(`���q��j�3`�
Dyǌ�����Q
;�bG]�����=�@�c��+� |�fl�=�����A�����9Õ���gT؋la��9�xv-�7U
r}���O�?Hǫ�zXXo�y,d����uJ&�`��(U�N���xL9(
h��4vW��x
=I��Q�Ί���5����fd��֕�r�y�?�$�������B������|��	ܲ�<h�5�%��12K��0o��	e?�d��
���4��'�J@]�����,l��ԍ��f;�0������n�8�t�F���.(�E֤1de�[Gc�%�޺���xR�W���WStC�����_ү�2���,F�Ӑp.��!�bl�Pۨ����܊U5ӏ���[��G�K��9��U;�8�N��b؟_31�.ѦF��l�0�� �]��O'
��nIqp�G���(���.X
(=�$f���/x��8��I�!�B^�%)T�,j�Po�t�-�cv�����D�8����e���"Jp�l�Ik�2�	9G�k�n��v!L̓>�Z/��CW{���Z�!;!V �J����c owhU����`V��mz�CΏɀ�ܱ܄q>�+n���aڶ#����݄�*L��i��J!�ڗ{9%�عN�Ki���<����b�*G�[��lC�V�g�0(Eu�>z'h���D9����1*���oEm�/k2��Qon��ʸ��(��J�c)��ױs��`�w��g��<�q6N8ʣz�����W[�E��0=Gt_
�5���)�E���,-P��>�/ssɶ'�va�v�qd�Z���e��Z,(��X�7҄�R�5������W?����� �a]Nx���Q��!h^�Y1lHJ8vZ���]����ku�@�//>rzaB��]��6��}w�e�C��\*?� �/�W� ���F1as�G�ԲL��Q�ds��i`{��c� s�%��Y�L
?�2Ф�>{��XF"�� ��<M�j>϶��i�U�v�!��%,���~�Kx�� kEpG��9�̌_[�	�J�x�8��̻��w�Q�{�M|��@ͺ%9��8� �D������n�v��t"�E���]�ڄ��˖'%4���}�D�?x噵�B�ؒ��R�^��Z5!�e�"�A��?�������S	�#�=o"�����s�(E�?s���D�6Hp�Q������# ���1S&��M�i�c̈́�3�Wep����XP��d�H,줘b_���̡�H�3���X��d�KW53��#u2�PS�<ݫ���}0���'_[	���@�����Lq>t$���2ѭ�.����`+)R^��&P�A3��{���U��D�,�k�8�D�p���yT(�=���i��G]����.���WJ]}���LU�r*-h�Ir�7$S���I��m��C#��
���sB�"���[ r�"쨗NpF[q��������EL*W_(N֜��7[���OGM�ċ�_68S�J�/�l_��E�f�:�8q��	#o��[o.�ul`�.@��Z%.�"�Y�~B�������P4�:F�s��n#��ݍI�"�z�5q���	Y��Y �P��)�e����@U��6�1�otm��F��뿹���ѹ�j�'�URN�N�� rrX�ɉĜ�����